magic
tech gf180mcuD
magscale 1 10
timestamp 1699642504
<< metal1 >>
rect 1344 38442 40656 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 40656 38442
rect 1344 38356 40656 38390
rect 25566 38274 25618 38286
rect 25566 38210 25618 38222
rect 18834 38110 18846 38162
rect 18898 38110 18910 38162
rect 22194 38110 22206 38162
rect 22258 38110 22270 38162
rect 18050 37998 18062 38050
rect 18114 37998 18126 38050
rect 23986 37998 23998 38050
rect 24050 37998 24062 38050
rect 24546 37998 24558 38050
rect 24610 37998 24622 38050
rect 1344 37658 40656 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 40656 37658
rect 1344 37572 40656 37606
rect 21422 37490 21474 37502
rect 21422 37426 21474 37438
rect 26238 37490 26290 37502
rect 26238 37426 26290 37438
rect 20402 37214 20414 37266
rect 20466 37214 20478 37266
rect 25330 37214 25342 37266
rect 25394 37214 25406 37266
rect 1344 36874 40656 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 40656 36874
rect 1344 36788 40656 36822
rect 24782 36706 24834 36718
rect 24782 36642 24834 36654
rect 23762 36430 23774 36482
rect 23826 36430 23838 36482
rect 1344 36090 40656 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 40656 36090
rect 1344 36004 40656 36038
rect 1344 35306 40656 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 40656 35306
rect 1344 35220 40656 35254
rect 1344 34522 40656 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 40656 34522
rect 1344 34436 40656 34470
rect 1344 33738 40656 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 40656 33738
rect 1344 33652 40656 33686
rect 1344 32954 40656 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 40656 32954
rect 1344 32868 40656 32902
rect 1344 32170 40656 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 40656 32170
rect 1344 32084 40656 32118
rect 1344 31386 40656 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 40656 31386
rect 1344 31300 40656 31334
rect 1344 30602 40656 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 40656 30602
rect 1344 30516 40656 30550
rect 1344 29818 40656 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 40656 29818
rect 1344 29732 40656 29766
rect 1344 29034 40656 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 40656 29034
rect 1344 28948 40656 28982
rect 23426 28590 23438 28642
rect 23490 28590 23502 28642
rect 23650 28478 23662 28530
rect 23714 28478 23726 28530
rect 1344 28250 40656 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 40656 28250
rect 1344 28164 40656 28198
rect 17378 27806 17390 27858
rect 17442 27806 17454 27858
rect 21298 27806 21310 27858
rect 21362 27806 21374 27858
rect 20862 27746 20914 27758
rect 24110 27746 24162 27758
rect 18162 27694 18174 27746
rect 18226 27694 18238 27746
rect 20290 27694 20302 27746
rect 20354 27694 20366 27746
rect 21970 27694 21982 27746
rect 22034 27694 22046 27746
rect 20862 27682 20914 27694
rect 24110 27682 24162 27694
rect 25454 27746 25506 27758
rect 25454 27682 25506 27694
rect 1344 27466 40656 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 40656 27466
rect 1344 27380 40656 27414
rect 20078 27298 20130 27310
rect 20078 27234 20130 27246
rect 21646 27298 21698 27310
rect 21646 27234 21698 27246
rect 40014 27186 40066 27198
rect 18834 27134 18846 27186
rect 18898 27134 18910 27186
rect 40014 27122 40066 27134
rect 19742 27074 19794 27086
rect 16034 27022 16046 27074
rect 16098 27022 16110 27074
rect 23426 27022 23438 27074
rect 23490 27022 23502 27074
rect 37874 27022 37886 27074
rect 37938 27022 37950 27074
rect 19742 27010 19794 27022
rect 19406 26962 19458 26974
rect 16706 26910 16718 26962
rect 16770 26910 16782 26962
rect 19406 26898 19458 26910
rect 19518 26962 19570 26974
rect 19518 26898 19570 26910
rect 20078 26962 20130 26974
rect 20078 26898 20130 26910
rect 20190 26962 20242 26974
rect 20190 26898 20242 26910
rect 21758 26962 21810 26974
rect 21758 26898 21810 26910
rect 22318 26962 22370 26974
rect 22318 26898 22370 26910
rect 22542 26962 22594 26974
rect 22542 26898 22594 26910
rect 22654 26962 22706 26974
rect 23650 26910 23662 26962
rect 23714 26910 23726 26962
rect 22654 26898 22706 26910
rect 21646 26850 21698 26862
rect 21646 26786 21698 26798
rect 1344 26682 40656 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 40656 26682
rect 1344 26596 40656 26630
rect 18622 26514 18674 26526
rect 18622 26450 18674 26462
rect 17502 26402 17554 26414
rect 17502 26338 17554 26350
rect 18398 26402 18450 26414
rect 18398 26338 18450 26350
rect 18734 26402 18786 26414
rect 18734 26338 18786 26350
rect 17390 26290 17442 26302
rect 4274 26238 4286 26290
rect 4338 26238 4350 26290
rect 15698 26238 15710 26290
rect 15762 26238 15774 26290
rect 20402 26238 20414 26290
rect 20466 26238 20478 26290
rect 25554 26238 25566 26290
rect 25618 26238 25630 26290
rect 37650 26238 37662 26290
rect 37714 26238 37726 26290
rect 17390 26226 17442 26238
rect 16158 26178 16210 26190
rect 12786 26126 12798 26178
rect 12850 26126 12862 26178
rect 14914 26126 14926 26178
rect 14978 26126 14990 26178
rect 16158 26114 16210 26126
rect 19182 26178 19234 26190
rect 19182 26114 19234 26126
rect 20078 26178 20130 26190
rect 28926 26178 28978 26190
rect 21186 26126 21198 26178
rect 21250 26126 21262 26178
rect 23314 26126 23326 26178
rect 23378 26126 23390 26178
rect 26338 26126 26350 26178
rect 26402 26126 26414 26178
rect 28466 26126 28478 26178
rect 28530 26126 28542 26178
rect 20078 26114 20130 26126
rect 28926 26114 28978 26126
rect 29486 26178 29538 26190
rect 29486 26114 29538 26126
rect 29934 26178 29986 26190
rect 39890 26126 39902 26178
rect 39954 26126 39966 26178
rect 29934 26114 29986 26126
rect 1934 26066 1986 26078
rect 1934 26002 1986 26014
rect 17502 26066 17554 26078
rect 17502 26002 17554 26014
rect 29038 26066 29090 26078
rect 29250 26014 29262 26066
rect 29314 26063 29326 26066
rect 30034 26063 30046 26066
rect 29314 26017 30046 26063
rect 29314 26014 29326 26017
rect 30034 26014 30046 26017
rect 30098 26014 30110 26066
rect 29038 26002 29090 26014
rect 1344 25898 40656 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 40656 25898
rect 1344 25812 40656 25846
rect 28254 25730 28306 25742
rect 28254 25666 28306 25678
rect 40014 25618 40066 25630
rect 2034 25566 2046 25618
rect 2098 25566 2110 25618
rect 27794 25566 27806 25618
rect 27858 25566 27870 25618
rect 29922 25566 29934 25618
rect 29986 25566 29998 25618
rect 32050 25566 32062 25618
rect 32114 25566 32126 25618
rect 40014 25554 40066 25566
rect 15038 25506 15090 25518
rect 4274 25454 4286 25506
rect 4338 25454 4350 25506
rect 15038 25442 15090 25454
rect 15262 25506 15314 25518
rect 15262 25442 15314 25454
rect 15710 25506 15762 25518
rect 15710 25442 15762 25454
rect 16046 25506 16098 25518
rect 16046 25442 16098 25454
rect 21422 25506 21474 25518
rect 21422 25442 21474 25454
rect 21646 25506 21698 25518
rect 21646 25442 21698 25454
rect 21982 25506 22034 25518
rect 21982 25442 22034 25454
rect 22206 25506 22258 25518
rect 22206 25442 22258 25454
rect 23102 25506 23154 25518
rect 24994 25454 25006 25506
rect 25058 25454 25070 25506
rect 25666 25454 25678 25506
rect 25730 25454 25742 25506
rect 29138 25454 29150 25506
rect 29202 25454 29214 25506
rect 37650 25454 37662 25506
rect 37714 25454 37726 25506
rect 23102 25442 23154 25454
rect 14254 25394 14306 25406
rect 14254 25330 14306 25342
rect 15486 25394 15538 25406
rect 15486 25330 15538 25342
rect 15934 25394 15986 25406
rect 15934 25330 15986 25342
rect 23326 25394 23378 25406
rect 23326 25330 23378 25342
rect 23438 25394 23490 25406
rect 23438 25330 23490 25342
rect 28142 25394 28194 25406
rect 28142 25330 28194 25342
rect 28254 25394 28306 25406
rect 28254 25330 28306 25342
rect 14366 25282 14418 25294
rect 14366 25218 14418 25230
rect 14590 25282 14642 25294
rect 14590 25218 14642 25230
rect 15262 25282 15314 25294
rect 15262 25218 15314 25230
rect 20750 25282 20802 25294
rect 20750 25218 20802 25230
rect 21310 25282 21362 25294
rect 22878 25282 22930 25294
rect 22530 25230 22542 25282
rect 22594 25230 22606 25282
rect 21310 25218 21362 25230
rect 22878 25218 22930 25230
rect 1344 25114 40656 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 40656 25114
rect 1344 25028 40656 25062
rect 21422 24946 21474 24958
rect 26686 24946 26738 24958
rect 22866 24894 22878 24946
rect 22930 24894 22942 24946
rect 21422 24882 21474 24894
rect 26686 24882 26738 24894
rect 27470 24946 27522 24958
rect 27470 24882 27522 24894
rect 28366 24946 28418 24958
rect 28366 24882 28418 24894
rect 29038 24946 29090 24958
rect 29038 24882 29090 24894
rect 29150 24946 29202 24958
rect 29150 24882 29202 24894
rect 14926 24834 14978 24846
rect 25454 24834 25506 24846
rect 13682 24782 13694 24834
rect 13746 24782 13758 24834
rect 18834 24782 18846 24834
rect 18898 24782 18910 24834
rect 14926 24770 14978 24782
rect 25454 24770 25506 24782
rect 27582 24834 27634 24846
rect 27582 24770 27634 24782
rect 14814 24722 14866 24734
rect 14354 24670 14366 24722
rect 14418 24670 14430 24722
rect 14814 24658 14866 24670
rect 15038 24722 15090 24734
rect 15038 24658 15090 24670
rect 15262 24722 15314 24734
rect 22542 24722 22594 24734
rect 26462 24722 26514 24734
rect 27694 24722 27746 24734
rect 18050 24670 18062 24722
rect 18114 24670 18126 24722
rect 25666 24670 25678 24722
rect 25730 24670 25742 24722
rect 25890 24670 25902 24722
rect 25954 24670 25966 24722
rect 26226 24670 26238 24722
rect 26290 24670 26302 24722
rect 26898 24670 26910 24722
rect 26962 24670 26974 24722
rect 27234 24670 27246 24722
rect 27298 24670 27310 24722
rect 15262 24658 15314 24670
rect 22542 24658 22594 24670
rect 26462 24658 26514 24670
rect 27694 24658 27746 24670
rect 27806 24722 27858 24734
rect 28926 24722 28978 24734
rect 28690 24670 28702 24722
rect 28754 24670 28766 24722
rect 27806 24658 27858 24670
rect 28926 24658 28978 24670
rect 29262 24722 29314 24734
rect 29262 24658 29314 24670
rect 25790 24610 25842 24622
rect 11554 24558 11566 24610
rect 11618 24558 11630 24610
rect 20962 24558 20974 24610
rect 21026 24558 21038 24610
rect 26786 24558 26798 24610
rect 26850 24558 26862 24610
rect 25790 24546 25842 24558
rect 1344 24330 40656 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 40656 24330
rect 1344 24244 40656 24278
rect 19630 24162 19682 24174
rect 19630 24098 19682 24110
rect 1934 24050 1986 24062
rect 26462 24050 26514 24062
rect 9986 23998 9998 24050
rect 10050 23998 10062 24050
rect 12114 23998 12126 24050
rect 12178 23998 12190 24050
rect 13570 23998 13582 24050
rect 13634 23998 13646 24050
rect 1934 23986 1986 23998
rect 26462 23986 26514 23998
rect 14702 23938 14754 23950
rect 4274 23886 4286 23938
rect 4338 23886 4350 23938
rect 12898 23886 12910 23938
rect 12962 23886 12974 23938
rect 14702 23874 14754 23886
rect 26574 23938 26626 23950
rect 26574 23874 26626 23886
rect 26798 23938 26850 23950
rect 26798 23874 26850 23886
rect 28142 23938 28194 23950
rect 28142 23874 28194 23886
rect 13806 23826 13858 23838
rect 13806 23762 13858 23774
rect 19630 23826 19682 23838
rect 19630 23762 19682 23774
rect 19742 23826 19794 23838
rect 19742 23762 19794 23774
rect 26350 23826 26402 23838
rect 28466 23774 28478 23826
rect 28530 23774 28542 23826
rect 26350 23762 26402 23774
rect 13582 23714 13634 23726
rect 13582 23650 13634 23662
rect 1344 23546 40656 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 40656 23546
rect 1344 23460 40656 23494
rect 14366 23378 14418 23390
rect 14366 23314 14418 23326
rect 15598 23378 15650 23390
rect 15598 23314 15650 23326
rect 16718 23378 16770 23390
rect 16718 23314 16770 23326
rect 20750 23378 20802 23390
rect 20750 23314 20802 23326
rect 14030 23266 14082 23278
rect 14030 23202 14082 23214
rect 15934 23266 15986 23278
rect 15934 23202 15986 23214
rect 16494 23266 16546 23278
rect 21198 23266 21250 23278
rect 20402 23214 20414 23266
rect 20466 23214 20478 23266
rect 16494 23202 16546 23214
rect 21198 23202 21250 23214
rect 21982 23266 22034 23278
rect 21982 23202 22034 23214
rect 23102 23266 23154 23278
rect 26450 23214 26462 23266
rect 26514 23214 26526 23266
rect 23102 23202 23154 23214
rect 14254 23154 14306 23166
rect 14254 23090 14306 23102
rect 14478 23154 14530 23166
rect 15486 23154 15538 23166
rect 14690 23102 14702 23154
rect 14754 23102 14766 23154
rect 14478 23090 14530 23102
rect 15486 23090 15538 23102
rect 15710 23154 15762 23166
rect 15710 23090 15762 23102
rect 16382 23154 16434 23166
rect 16382 23090 16434 23102
rect 22990 23154 23042 23166
rect 22990 23090 23042 23102
rect 23326 23154 23378 23166
rect 23326 23090 23378 23102
rect 26126 23154 26178 23166
rect 26126 23090 26178 23102
rect 13134 23042 13186 23054
rect 22082 22990 22094 23042
rect 22146 22990 22158 23042
rect 13134 22978 13186 22990
rect 21310 22930 21362 22942
rect 21310 22866 21362 22878
rect 21758 22930 21810 22942
rect 21758 22866 21810 22878
rect 1344 22762 40656 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 40656 22762
rect 1344 22676 40656 22710
rect 19294 22594 19346 22606
rect 19294 22530 19346 22542
rect 26014 22482 26066 22494
rect 40014 22482 40066 22494
rect 16146 22430 16158 22482
rect 16210 22430 16222 22482
rect 23426 22430 23438 22482
rect 23490 22430 23502 22482
rect 25554 22430 25566 22482
rect 25618 22430 25630 22482
rect 32050 22430 32062 22482
rect 32114 22430 32126 22482
rect 26014 22418 26066 22430
rect 40014 22418 40066 22430
rect 14590 22370 14642 22382
rect 14590 22306 14642 22318
rect 14926 22370 14978 22382
rect 14926 22306 14978 22318
rect 15150 22370 15202 22382
rect 15150 22306 15202 22318
rect 19406 22370 19458 22382
rect 28254 22370 28306 22382
rect 20626 22318 20638 22370
rect 20690 22318 20702 22370
rect 21746 22318 21758 22370
rect 21810 22318 21822 22370
rect 22754 22318 22766 22370
rect 22818 22318 22830 22370
rect 19406 22306 19458 22318
rect 28254 22306 28306 22318
rect 28702 22370 28754 22382
rect 29138 22318 29150 22370
rect 29202 22318 29214 22370
rect 37650 22318 37662 22370
rect 37714 22318 37726 22370
rect 28702 22306 28754 22318
rect 15486 22258 15538 22270
rect 15486 22194 15538 22206
rect 15822 22258 15874 22270
rect 15822 22194 15874 22206
rect 16494 22258 16546 22270
rect 16494 22194 16546 22206
rect 16942 22258 16994 22270
rect 28142 22258 28194 22270
rect 17378 22206 17390 22258
rect 17442 22206 17454 22258
rect 29922 22206 29934 22258
rect 29986 22206 29998 22258
rect 16942 22194 16994 22206
rect 28142 22194 28194 22206
rect 14814 22146 14866 22158
rect 14814 22082 14866 22094
rect 16270 22146 16322 22158
rect 16270 22082 16322 22094
rect 16830 22146 16882 22158
rect 16830 22082 16882 22094
rect 17726 22146 17778 22158
rect 17726 22082 17778 22094
rect 19294 22146 19346 22158
rect 28030 22146 28082 22158
rect 20402 22094 20414 22146
rect 20466 22094 20478 22146
rect 21970 22094 21982 22146
rect 22034 22094 22046 22146
rect 19294 22082 19346 22094
rect 28030 22082 28082 22094
rect 1344 21978 40656 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 40656 21978
rect 1344 21892 40656 21926
rect 23102 21810 23154 21822
rect 15810 21758 15822 21810
rect 15874 21758 15886 21810
rect 23102 21746 23154 21758
rect 25566 21810 25618 21822
rect 25566 21746 25618 21758
rect 26238 21810 26290 21822
rect 26238 21746 26290 21758
rect 29710 21810 29762 21822
rect 29710 21746 29762 21758
rect 29934 21810 29986 21822
rect 29934 21746 29986 21758
rect 26126 21698 26178 21710
rect 13234 21646 13246 21698
rect 13298 21646 13310 21698
rect 24210 21646 24222 21698
rect 24274 21646 24286 21698
rect 26126 21634 26178 21646
rect 26350 21698 26402 21710
rect 26350 21634 26402 21646
rect 27134 21698 27186 21710
rect 27134 21634 27186 21646
rect 15150 21586 15202 21598
rect 22878 21586 22930 21598
rect 13906 21534 13918 21586
rect 13970 21534 13982 21586
rect 15586 21534 15598 21586
rect 15650 21534 15662 21586
rect 22642 21534 22654 21586
rect 22706 21534 22718 21586
rect 15150 21522 15202 21534
rect 22878 21522 22930 21534
rect 23326 21586 23378 21598
rect 23326 21522 23378 21534
rect 23550 21586 23602 21598
rect 23550 21522 23602 21534
rect 23886 21586 23938 21598
rect 23886 21522 23938 21534
rect 25454 21586 25506 21598
rect 25454 21522 25506 21534
rect 26910 21586 26962 21598
rect 26910 21522 26962 21534
rect 27582 21586 27634 21598
rect 27582 21522 27634 21534
rect 30046 21586 30098 21598
rect 37650 21534 37662 21586
rect 37714 21534 37726 21586
rect 30046 21522 30098 21534
rect 27022 21474 27074 21486
rect 11106 21422 11118 21474
rect 11170 21422 11182 21474
rect 17602 21422 17614 21474
rect 17666 21422 17678 21474
rect 27022 21410 27074 21422
rect 28814 21474 28866 21486
rect 28814 21410 28866 21422
rect 40014 21474 40066 21486
rect 40014 21410 40066 21422
rect 14254 21362 14306 21374
rect 14254 21298 14306 21310
rect 14702 21362 14754 21374
rect 14702 21298 14754 21310
rect 14926 21362 14978 21374
rect 14926 21298 14978 21310
rect 25566 21362 25618 21374
rect 25566 21298 25618 21310
rect 1344 21194 40656 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 40656 21194
rect 1344 21108 40656 21142
rect 17950 21026 18002 21038
rect 16258 20974 16270 21026
rect 16322 20974 16334 21026
rect 17950 20962 18002 20974
rect 18622 21026 18674 21038
rect 18622 20962 18674 20974
rect 40014 20914 40066 20926
rect 18274 20862 18286 20914
rect 18338 20862 18350 20914
rect 20290 20862 20302 20914
rect 20354 20862 20366 20914
rect 22418 20862 22430 20914
rect 22482 20862 22494 20914
rect 40014 20850 40066 20862
rect 16606 20802 16658 20814
rect 15698 20750 15710 20802
rect 15762 20750 15774 20802
rect 16606 20738 16658 20750
rect 16830 20802 16882 20814
rect 18958 20802 19010 20814
rect 17602 20750 17614 20802
rect 17666 20750 17678 20802
rect 16830 20738 16882 20750
rect 18958 20738 19010 20750
rect 19406 20802 19458 20814
rect 21982 20802 22034 20814
rect 20066 20750 20078 20802
rect 20130 20750 20142 20802
rect 20402 20750 20414 20802
rect 20466 20750 20478 20802
rect 19406 20738 19458 20750
rect 21982 20738 22034 20750
rect 22094 20802 22146 20814
rect 22094 20738 22146 20750
rect 22318 20802 22370 20814
rect 29038 20802 29090 20814
rect 22530 20750 22542 20802
rect 22594 20750 22606 20802
rect 23314 20750 23326 20802
rect 23378 20750 23390 20802
rect 22318 20738 22370 20750
rect 29038 20738 29090 20750
rect 29374 20802 29426 20814
rect 37650 20750 37662 20802
rect 37714 20750 37726 20802
rect 29374 20738 29426 20750
rect 17166 20690 17218 20702
rect 17166 20626 17218 20638
rect 18174 20690 18226 20702
rect 18174 20626 18226 20638
rect 19182 20690 19234 20702
rect 19182 20626 19234 20638
rect 21310 20690 21362 20702
rect 21310 20626 21362 20638
rect 21646 20690 21698 20702
rect 21646 20626 21698 20638
rect 22878 20690 22930 20702
rect 25442 20638 25454 20690
rect 25506 20638 25518 20690
rect 22878 20626 22930 20638
rect 14254 20578 14306 20590
rect 14254 20514 14306 20526
rect 15934 20578 15986 20590
rect 15934 20514 15986 20526
rect 17054 20578 17106 20590
rect 17054 20514 17106 20526
rect 17390 20578 17442 20590
rect 17390 20514 17442 20526
rect 21422 20578 21474 20590
rect 21422 20514 21474 20526
rect 22990 20578 23042 20590
rect 22990 20514 23042 20526
rect 29262 20578 29314 20590
rect 29262 20514 29314 20526
rect 1344 20410 40656 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 40656 20410
rect 1344 20324 40656 20358
rect 16494 20242 16546 20254
rect 16494 20178 16546 20190
rect 18062 20242 18114 20254
rect 25342 20242 25394 20254
rect 18386 20190 18398 20242
rect 18450 20190 18462 20242
rect 18062 20178 18114 20190
rect 25342 20178 25394 20190
rect 25566 20242 25618 20254
rect 25566 20178 25618 20190
rect 25790 20242 25842 20254
rect 25790 20178 25842 20190
rect 25902 20242 25954 20254
rect 25902 20178 25954 20190
rect 13694 20130 13746 20142
rect 13694 20066 13746 20078
rect 16718 20130 16770 20142
rect 16718 20066 16770 20078
rect 17726 20130 17778 20142
rect 17726 20066 17778 20078
rect 18734 20130 18786 20142
rect 18734 20066 18786 20078
rect 18958 20130 19010 20142
rect 30046 20130 30098 20142
rect 23314 20078 23326 20130
rect 23378 20078 23390 20130
rect 27570 20078 27582 20130
rect 27634 20078 27646 20130
rect 18958 20066 19010 20078
rect 30046 20066 30098 20078
rect 30158 20130 30210 20142
rect 30158 20066 30210 20078
rect 13470 20018 13522 20030
rect 4274 19966 4286 20018
rect 4338 19966 4350 20018
rect 13470 19954 13522 19966
rect 13806 20018 13858 20030
rect 13806 19954 13858 19966
rect 17390 20018 17442 20030
rect 17390 19954 17442 19966
rect 18846 20018 18898 20030
rect 25230 20018 25282 20030
rect 19730 19966 19742 20018
rect 19794 19966 19806 20018
rect 18846 19954 18898 19966
rect 25230 19954 25282 19966
rect 26014 20018 26066 20030
rect 26338 19966 26350 20018
rect 26402 19966 26414 20018
rect 26898 19966 26910 20018
rect 26962 19966 26974 20018
rect 37650 19966 37662 20018
rect 37714 19966 37726 20018
rect 26014 19954 26066 19966
rect 13134 19906 13186 19918
rect 13134 19842 13186 19854
rect 16606 19906 16658 19918
rect 30718 19906 30770 19918
rect 29698 19854 29710 19906
rect 29762 19854 29774 19906
rect 16606 19842 16658 19854
rect 30718 19842 30770 19854
rect 1934 19794 1986 19806
rect 1934 19730 1986 19742
rect 30158 19794 30210 19806
rect 30158 19730 30210 19742
rect 40014 19794 40066 19806
rect 40014 19730 40066 19742
rect 1344 19626 40656 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 40656 19626
rect 1344 19540 40656 19574
rect 15262 19458 15314 19470
rect 15262 19394 15314 19406
rect 17614 19458 17666 19470
rect 17614 19394 17666 19406
rect 23438 19458 23490 19470
rect 23438 19394 23490 19406
rect 23774 19458 23826 19470
rect 23774 19394 23826 19406
rect 16046 19346 16098 19358
rect 9986 19294 9998 19346
rect 10050 19294 10062 19346
rect 16046 19282 16098 19294
rect 17726 19346 17778 19358
rect 32050 19294 32062 19346
rect 32114 19294 32126 19346
rect 17726 19282 17778 19294
rect 13470 19234 13522 19246
rect 12898 19182 12910 19234
rect 12962 19182 12974 19234
rect 13470 19170 13522 19182
rect 13806 19234 13858 19246
rect 13806 19170 13858 19182
rect 14030 19234 14082 19246
rect 14030 19170 14082 19182
rect 15374 19234 15426 19246
rect 15374 19170 15426 19182
rect 16270 19234 16322 19246
rect 16270 19170 16322 19182
rect 20302 19234 20354 19246
rect 20302 19170 20354 19182
rect 20526 19234 20578 19246
rect 20526 19170 20578 19182
rect 20862 19234 20914 19246
rect 20862 19170 20914 19182
rect 21198 19234 21250 19246
rect 24110 19234 24162 19246
rect 21522 19182 21534 19234
rect 21586 19182 21598 19234
rect 22418 19182 22430 19234
rect 22482 19182 22494 19234
rect 22866 19182 22878 19234
rect 22930 19182 22942 19234
rect 21198 19170 21250 19182
rect 24110 19170 24162 19182
rect 25678 19234 25730 19246
rect 25678 19170 25730 19182
rect 28702 19234 28754 19246
rect 29250 19182 29262 19234
rect 29314 19182 29326 19234
rect 28702 19170 28754 19182
rect 13582 19122 13634 19134
rect 12114 19070 12126 19122
rect 12178 19070 12190 19122
rect 13582 19058 13634 19070
rect 18286 19122 18338 19134
rect 18286 19058 18338 19070
rect 18958 19122 19010 19134
rect 18958 19058 19010 19070
rect 19070 19122 19122 19134
rect 19070 19058 19122 19070
rect 19966 19122 20018 19134
rect 19966 19058 20018 19070
rect 20078 19122 20130 19134
rect 20078 19058 20130 19070
rect 20638 19122 20690 19134
rect 20638 19058 20690 19070
rect 21758 19122 21810 19134
rect 21758 19058 21810 19070
rect 22318 19122 22370 19134
rect 22318 19058 22370 19070
rect 23662 19122 23714 19134
rect 23662 19058 23714 19070
rect 24446 19122 24498 19134
rect 24446 19058 24498 19070
rect 28142 19122 28194 19134
rect 29922 19070 29934 19122
rect 29986 19070 29998 19122
rect 28142 19058 28194 19070
rect 15262 19010 15314 19022
rect 16942 19010 16994 19022
rect 17950 19010 18002 19022
rect 16594 18958 16606 19010
rect 16658 18958 16670 19010
rect 17266 18958 17278 19010
rect 17330 18958 17342 19010
rect 15262 18946 15314 18958
rect 16942 18946 16994 18958
rect 17950 18946 18002 18958
rect 18174 19010 18226 19022
rect 18174 18946 18226 18958
rect 19294 19010 19346 19022
rect 19294 18946 19346 18958
rect 19742 19010 19794 19022
rect 19742 18946 19794 18958
rect 21870 19010 21922 19022
rect 21870 18946 21922 18958
rect 24782 19010 24834 19022
rect 25342 19010 25394 19022
rect 25106 18958 25118 19010
rect 25170 18958 25182 19010
rect 24782 18946 24834 18958
rect 25342 18946 25394 18958
rect 25566 19010 25618 19022
rect 25566 18946 25618 18958
rect 28030 19010 28082 19022
rect 28030 18946 28082 18958
rect 28254 19010 28306 19022
rect 28254 18946 28306 18958
rect 1344 18842 40656 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 40656 18842
rect 1344 18756 40656 18790
rect 16830 18674 16882 18686
rect 16830 18610 16882 18622
rect 22766 18674 22818 18686
rect 22766 18610 22818 18622
rect 24222 18674 24274 18686
rect 24222 18610 24274 18622
rect 28814 18674 28866 18686
rect 28814 18610 28866 18622
rect 13358 18562 13410 18574
rect 13358 18498 13410 18510
rect 13470 18562 13522 18574
rect 22990 18562 23042 18574
rect 18610 18510 18622 18562
rect 18674 18510 18686 18562
rect 21746 18510 21758 18562
rect 21810 18510 21822 18562
rect 13470 18498 13522 18510
rect 22990 18498 23042 18510
rect 23886 18562 23938 18574
rect 23886 18498 23938 18510
rect 23998 18562 24050 18574
rect 23998 18498 24050 18510
rect 26238 18562 26290 18574
rect 26238 18498 26290 18510
rect 27358 18562 27410 18574
rect 27358 18498 27410 18510
rect 27470 18562 27522 18574
rect 27470 18498 27522 18510
rect 13694 18450 13746 18462
rect 4274 18398 4286 18450
rect 4338 18398 4350 18450
rect 13694 18386 13746 18398
rect 13806 18450 13858 18462
rect 17726 18450 17778 18462
rect 14130 18398 14142 18450
rect 14194 18398 14206 18450
rect 16594 18398 16606 18450
rect 16658 18398 16670 18450
rect 13806 18386 13858 18398
rect 17726 18386 17778 18398
rect 17950 18450 18002 18462
rect 22542 18450 22594 18462
rect 18386 18398 18398 18450
rect 18450 18398 18462 18450
rect 21522 18398 21534 18450
rect 21586 18398 21598 18450
rect 17950 18386 18002 18398
rect 22542 18386 22594 18398
rect 23214 18450 23266 18462
rect 23214 18386 23266 18398
rect 25790 18450 25842 18462
rect 25790 18386 25842 18398
rect 26014 18450 26066 18462
rect 26014 18386 26066 18398
rect 26462 18450 26514 18462
rect 26462 18386 26514 18398
rect 27694 18450 27746 18462
rect 27694 18386 27746 18398
rect 14590 18338 14642 18350
rect 14590 18274 14642 18286
rect 15038 18338 15090 18350
rect 25454 18338 25506 18350
rect 21970 18286 21982 18338
rect 22034 18286 22046 18338
rect 15038 18274 15090 18286
rect 25454 18274 25506 18286
rect 1934 18226 1986 18238
rect 1934 18162 1986 18174
rect 14478 18226 14530 18238
rect 22654 18226 22706 18238
rect 17378 18174 17390 18226
rect 17442 18174 17454 18226
rect 14478 18162 14530 18174
rect 22654 18162 22706 18174
rect 1344 18058 40656 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 40656 18058
rect 1344 17972 40656 18006
rect 22430 17890 22482 17902
rect 15138 17838 15150 17890
rect 15202 17838 15214 17890
rect 22430 17826 22482 17838
rect 22206 17778 22258 17790
rect 9986 17726 9998 17778
rect 10050 17726 10062 17778
rect 12114 17726 12126 17778
rect 12178 17726 12190 17778
rect 22206 17714 22258 17726
rect 23662 17778 23714 17790
rect 40014 17778 40066 17790
rect 27234 17726 27246 17778
rect 27298 17726 27310 17778
rect 23662 17714 23714 17726
rect 40014 17714 40066 17726
rect 15486 17666 15538 17678
rect 12898 17614 12910 17666
rect 12962 17614 12974 17666
rect 15486 17602 15538 17614
rect 15710 17666 15762 17678
rect 15710 17602 15762 17614
rect 16382 17666 16434 17678
rect 23550 17666 23602 17678
rect 26126 17666 26178 17678
rect 17602 17614 17614 17666
rect 17666 17614 17678 17666
rect 21410 17614 21422 17666
rect 21474 17614 21486 17666
rect 23986 17614 23998 17666
rect 24050 17614 24062 17666
rect 24322 17614 24334 17666
rect 24386 17614 24398 17666
rect 16382 17602 16434 17614
rect 23550 17602 23602 17614
rect 26126 17602 26178 17614
rect 26462 17666 26514 17678
rect 26462 17602 26514 17614
rect 27582 17666 27634 17678
rect 28354 17614 28366 17666
rect 28418 17614 28430 17666
rect 37650 17614 37662 17666
rect 37714 17614 37726 17666
rect 27582 17602 27634 17614
rect 26798 17554 26850 17566
rect 27918 17554 27970 17566
rect 21634 17502 21646 17554
rect 21698 17502 21710 17554
rect 26898 17502 26910 17554
rect 26962 17502 26974 17554
rect 26798 17490 26850 17502
rect 27918 17490 27970 17502
rect 13582 17442 13634 17454
rect 13582 17378 13634 17390
rect 16046 17442 16098 17454
rect 23774 17442 23826 17454
rect 17826 17390 17838 17442
rect 17890 17390 17902 17442
rect 22754 17390 22766 17442
rect 22818 17390 22830 17442
rect 16046 17378 16098 17390
rect 23774 17378 23826 17390
rect 24894 17442 24946 17454
rect 26686 17442 26738 17454
rect 25218 17390 25230 17442
rect 25282 17390 25294 17442
rect 25778 17390 25790 17442
rect 25842 17390 25854 17442
rect 24894 17378 24946 17390
rect 26686 17378 26738 17390
rect 27694 17442 27746 17454
rect 27694 17378 27746 17390
rect 27806 17442 27858 17454
rect 27806 17378 27858 17390
rect 1344 17274 40656 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 40656 17274
rect 1344 17188 40656 17222
rect 26686 17106 26738 17118
rect 21746 17054 21758 17106
rect 21810 17054 21822 17106
rect 26686 17042 26738 17054
rect 14466 16942 14478 16994
rect 14530 16942 14542 16994
rect 27794 16942 27806 16994
rect 27858 16942 27870 16994
rect 17502 16882 17554 16894
rect 21422 16882 21474 16894
rect 13794 16830 13806 16882
rect 13858 16830 13870 16882
rect 17826 16830 17838 16882
rect 17890 16830 17902 16882
rect 27010 16830 27022 16882
rect 27074 16830 27086 16882
rect 37650 16830 37662 16882
rect 37714 16830 37726 16882
rect 17502 16818 17554 16830
rect 21422 16818 21474 16830
rect 18062 16770 18114 16782
rect 40014 16770 40066 16782
rect 16594 16718 16606 16770
rect 16658 16718 16670 16770
rect 29922 16718 29934 16770
rect 29986 16718 29998 16770
rect 18062 16706 18114 16718
rect 40014 16706 40066 16718
rect 18174 16658 18226 16670
rect 18174 16594 18226 16606
rect 1344 16490 40656 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 40656 16490
rect 1344 16404 40656 16438
rect 21310 16322 21362 16334
rect 20402 16270 20414 16322
rect 20466 16270 20478 16322
rect 21310 16258 21362 16270
rect 21646 16322 21698 16334
rect 21646 16258 21698 16270
rect 28142 16210 28194 16222
rect 27234 16158 27246 16210
rect 27298 16158 27310 16210
rect 28142 16146 28194 16158
rect 18286 16098 18338 16110
rect 18286 16034 18338 16046
rect 18958 16098 19010 16110
rect 18958 16034 19010 16046
rect 19854 16098 19906 16110
rect 22766 16098 22818 16110
rect 20066 16046 20078 16098
rect 20130 16046 20142 16098
rect 20626 16046 20638 16098
rect 20690 16046 20702 16098
rect 21298 16046 21310 16098
rect 21362 16046 21374 16098
rect 19854 16034 19906 16046
rect 22766 16034 22818 16046
rect 26910 16098 26962 16110
rect 27682 16046 27694 16098
rect 27746 16046 27758 16098
rect 26910 16034 26962 16046
rect 18510 15986 18562 15998
rect 18510 15922 18562 15934
rect 27246 15986 27298 15998
rect 27246 15922 27298 15934
rect 18622 15874 18674 15886
rect 18622 15810 18674 15822
rect 19966 15874 20018 15886
rect 19966 15810 20018 15822
rect 22430 15874 22482 15886
rect 22430 15810 22482 15822
rect 27134 15874 27186 15886
rect 27134 15810 27186 15822
rect 1344 15706 40656 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 40656 15706
rect 1344 15620 40656 15654
rect 27022 15538 27074 15550
rect 27022 15474 27074 15486
rect 26238 15426 26290 15438
rect 19058 15374 19070 15426
rect 19122 15374 19134 15426
rect 22306 15374 22318 15426
rect 22370 15374 22382 15426
rect 28690 15374 28702 15426
rect 28754 15374 28766 15426
rect 26238 15362 26290 15374
rect 25342 15314 25394 15326
rect 18386 15262 18398 15314
rect 18450 15262 18462 15314
rect 21634 15262 21646 15314
rect 21698 15262 21710 15314
rect 25342 15250 25394 15262
rect 26350 15314 26402 15326
rect 26350 15250 26402 15262
rect 26686 15314 26738 15326
rect 26686 15250 26738 15262
rect 26910 15314 26962 15326
rect 26910 15250 26962 15262
rect 27246 15314 27298 15326
rect 28018 15262 28030 15314
rect 28082 15262 28094 15314
rect 27246 15250 27298 15262
rect 21186 15150 21198 15202
rect 21250 15150 21262 15202
rect 24434 15150 24446 15202
rect 24498 15150 24510 15202
rect 30818 15150 30830 15202
rect 30882 15150 30894 15202
rect 1344 14922 40656 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 40656 14922
rect 1344 14836 40656 14870
rect 20862 14642 20914 14654
rect 18162 14590 18174 14642
rect 18226 14590 18238 14642
rect 20290 14590 20302 14642
rect 20354 14590 20366 14642
rect 20862 14578 20914 14590
rect 21422 14642 21474 14654
rect 29262 14642 29314 14654
rect 26450 14590 26462 14642
rect 26514 14590 26526 14642
rect 28578 14590 28590 14642
rect 28642 14590 28654 14642
rect 21422 14578 21474 14590
rect 29262 14578 29314 14590
rect 40014 14642 40066 14654
rect 40014 14578 40066 14590
rect 23886 14530 23938 14542
rect 17490 14478 17502 14530
rect 17554 14478 17566 14530
rect 23886 14466 23938 14478
rect 24222 14530 24274 14542
rect 24222 14466 24274 14478
rect 24558 14530 24610 14542
rect 24558 14466 24610 14478
rect 25006 14530 25058 14542
rect 25006 14466 25058 14478
rect 25342 14530 25394 14542
rect 25666 14478 25678 14530
rect 25730 14478 25742 14530
rect 37650 14478 37662 14530
rect 37714 14478 37726 14530
rect 25342 14466 25394 14478
rect 24222 14306 24274 14318
rect 24222 14242 24274 14254
rect 25230 14306 25282 14318
rect 25230 14242 25282 14254
rect 1344 14138 40656 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 40656 14138
rect 1344 14052 40656 14086
rect 26462 13970 26514 13982
rect 26462 13906 26514 13918
rect 27246 13970 27298 13982
rect 27246 13906 27298 13918
rect 27470 13970 27522 13982
rect 27470 13906 27522 13918
rect 27582 13858 27634 13870
rect 26114 13806 26126 13858
rect 26178 13806 26190 13858
rect 26786 13806 26798 13858
rect 26850 13806 26862 13858
rect 27582 13794 27634 13806
rect 25790 13746 25842 13758
rect 25790 13682 25842 13694
rect 1344 13354 40656 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 40656 13354
rect 1344 13268 40656 13302
rect 26462 13074 26514 13086
rect 23762 13022 23774 13074
rect 23826 13022 23838 13074
rect 25890 13022 25902 13074
rect 25954 13022 25966 13074
rect 26462 13010 26514 13022
rect 22978 12910 22990 12962
rect 23042 12910 23054 12962
rect 1344 12570 40656 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 40656 12570
rect 1344 12484 40656 12518
rect 1344 11786 40656 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 40656 11786
rect 1344 11700 40656 11734
rect 1344 11002 40656 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 40656 11002
rect 1344 10916 40656 10950
rect 1344 10218 40656 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 40656 10218
rect 1344 10132 40656 10166
rect 1344 9434 40656 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 40656 9434
rect 1344 9348 40656 9382
rect 1344 8650 40656 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 40656 8650
rect 1344 8564 40656 8598
rect 1344 7866 40656 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 40656 7866
rect 1344 7780 40656 7814
rect 1344 7082 40656 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 40656 7082
rect 1344 6996 40656 7030
rect 1344 6298 40656 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 40656 6298
rect 1344 6212 40656 6246
rect 1344 5514 40656 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 40656 5514
rect 1344 5428 40656 5462
rect 1344 4730 40656 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 40656 4730
rect 1344 4644 40656 4678
rect 25778 4286 25790 4338
rect 25842 4286 25854 4338
rect 28690 4286 28702 4338
rect 28754 4286 28766 4338
rect 26798 4114 26850 4126
rect 26798 4050 26850 4062
rect 29710 4114 29762 4126
rect 29710 4050 29762 4062
rect 1344 3946 40656 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 40656 3946
rect 1344 3860 40656 3894
rect 22430 3666 22482 3678
rect 22430 3602 22482 3614
rect 25566 3666 25618 3678
rect 25566 3602 25618 3614
rect 29374 3666 29426 3678
rect 29374 3602 29426 3614
rect 21410 3502 21422 3554
rect 21474 3502 21486 3554
rect 24546 3502 24558 3554
rect 24610 3502 24622 3554
rect 28578 3502 28590 3554
rect 28642 3502 28654 3554
rect 1344 3162 40656 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 40656 3162
rect 1344 3076 40656 3110
<< via1 >>
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 25566 38222 25618 38274
rect 18846 38110 18898 38162
rect 22206 38110 22258 38162
rect 18062 37998 18114 38050
rect 23998 37998 24050 38050
rect 24558 37998 24610 38050
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 21422 37438 21474 37490
rect 26238 37438 26290 37490
rect 20414 37214 20466 37266
rect 25342 37214 25394 37266
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 24782 36654 24834 36706
rect 23774 36430 23826 36482
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 23438 28590 23490 28642
rect 23662 28478 23714 28530
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 17390 27806 17442 27858
rect 21310 27806 21362 27858
rect 18174 27694 18226 27746
rect 20302 27694 20354 27746
rect 20862 27694 20914 27746
rect 21982 27694 22034 27746
rect 24110 27694 24162 27746
rect 25454 27694 25506 27746
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 20078 27246 20130 27298
rect 21646 27246 21698 27298
rect 18846 27134 18898 27186
rect 40014 27134 40066 27186
rect 16046 27022 16098 27074
rect 19742 27022 19794 27074
rect 23438 27022 23490 27074
rect 37886 27022 37938 27074
rect 16718 26910 16770 26962
rect 19406 26910 19458 26962
rect 19518 26910 19570 26962
rect 20078 26910 20130 26962
rect 20190 26910 20242 26962
rect 21758 26910 21810 26962
rect 22318 26910 22370 26962
rect 22542 26910 22594 26962
rect 22654 26910 22706 26962
rect 23662 26910 23714 26962
rect 21646 26798 21698 26850
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 18622 26462 18674 26514
rect 17502 26350 17554 26402
rect 18398 26350 18450 26402
rect 18734 26350 18786 26402
rect 4286 26238 4338 26290
rect 15710 26238 15762 26290
rect 17390 26238 17442 26290
rect 20414 26238 20466 26290
rect 25566 26238 25618 26290
rect 37662 26238 37714 26290
rect 12798 26126 12850 26178
rect 14926 26126 14978 26178
rect 16158 26126 16210 26178
rect 19182 26126 19234 26178
rect 20078 26126 20130 26178
rect 21198 26126 21250 26178
rect 23326 26126 23378 26178
rect 26350 26126 26402 26178
rect 28478 26126 28530 26178
rect 28926 26126 28978 26178
rect 29486 26126 29538 26178
rect 29934 26126 29986 26178
rect 39902 26126 39954 26178
rect 1934 26014 1986 26066
rect 17502 26014 17554 26066
rect 29038 26014 29090 26066
rect 29262 26014 29314 26066
rect 30046 26014 30098 26066
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 28254 25678 28306 25730
rect 2046 25566 2098 25618
rect 27806 25566 27858 25618
rect 29934 25566 29986 25618
rect 32062 25566 32114 25618
rect 40014 25566 40066 25618
rect 4286 25454 4338 25506
rect 15038 25454 15090 25506
rect 15262 25454 15314 25506
rect 15710 25454 15762 25506
rect 16046 25454 16098 25506
rect 21422 25454 21474 25506
rect 21646 25454 21698 25506
rect 21982 25454 22034 25506
rect 22206 25454 22258 25506
rect 23102 25454 23154 25506
rect 25006 25454 25058 25506
rect 25678 25454 25730 25506
rect 29150 25454 29202 25506
rect 37662 25454 37714 25506
rect 14254 25342 14306 25394
rect 15486 25342 15538 25394
rect 15934 25342 15986 25394
rect 23326 25342 23378 25394
rect 23438 25342 23490 25394
rect 28142 25342 28194 25394
rect 28254 25342 28306 25394
rect 14366 25230 14418 25282
rect 14590 25230 14642 25282
rect 15262 25230 15314 25282
rect 20750 25230 20802 25282
rect 21310 25230 21362 25282
rect 22542 25230 22594 25282
rect 22878 25230 22930 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 21422 24894 21474 24946
rect 22878 24894 22930 24946
rect 26686 24894 26738 24946
rect 27470 24894 27522 24946
rect 28366 24894 28418 24946
rect 29038 24894 29090 24946
rect 29150 24894 29202 24946
rect 13694 24782 13746 24834
rect 14926 24782 14978 24834
rect 18846 24782 18898 24834
rect 25454 24782 25506 24834
rect 27582 24782 27634 24834
rect 14366 24670 14418 24722
rect 14814 24670 14866 24722
rect 15038 24670 15090 24722
rect 15262 24670 15314 24722
rect 18062 24670 18114 24722
rect 22542 24670 22594 24722
rect 25678 24670 25730 24722
rect 25902 24670 25954 24722
rect 26238 24670 26290 24722
rect 26462 24670 26514 24722
rect 26910 24670 26962 24722
rect 27246 24670 27298 24722
rect 27694 24670 27746 24722
rect 27806 24670 27858 24722
rect 28702 24670 28754 24722
rect 28926 24670 28978 24722
rect 29262 24670 29314 24722
rect 11566 24558 11618 24610
rect 20974 24558 21026 24610
rect 25790 24558 25842 24610
rect 26798 24558 26850 24610
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 19630 24110 19682 24162
rect 1934 23998 1986 24050
rect 9998 23998 10050 24050
rect 12126 23998 12178 24050
rect 13582 23998 13634 24050
rect 26462 23998 26514 24050
rect 4286 23886 4338 23938
rect 12910 23886 12962 23938
rect 14702 23886 14754 23938
rect 26574 23886 26626 23938
rect 26798 23886 26850 23938
rect 28142 23886 28194 23938
rect 13806 23774 13858 23826
rect 19630 23774 19682 23826
rect 19742 23774 19794 23826
rect 26350 23774 26402 23826
rect 28478 23774 28530 23826
rect 13582 23662 13634 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 14366 23326 14418 23378
rect 15598 23326 15650 23378
rect 16718 23326 16770 23378
rect 20750 23326 20802 23378
rect 14030 23214 14082 23266
rect 15934 23214 15986 23266
rect 16494 23214 16546 23266
rect 20414 23214 20466 23266
rect 21198 23214 21250 23266
rect 21982 23214 22034 23266
rect 23102 23214 23154 23266
rect 26462 23214 26514 23266
rect 14254 23102 14306 23154
rect 14478 23102 14530 23154
rect 14702 23102 14754 23154
rect 15486 23102 15538 23154
rect 15710 23102 15762 23154
rect 16382 23102 16434 23154
rect 22990 23102 23042 23154
rect 23326 23102 23378 23154
rect 26126 23102 26178 23154
rect 13134 22990 13186 23042
rect 22094 22990 22146 23042
rect 21310 22878 21362 22930
rect 21758 22878 21810 22930
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 19294 22542 19346 22594
rect 16158 22430 16210 22482
rect 23438 22430 23490 22482
rect 25566 22430 25618 22482
rect 26014 22430 26066 22482
rect 32062 22430 32114 22482
rect 40014 22430 40066 22482
rect 14590 22318 14642 22370
rect 14926 22318 14978 22370
rect 15150 22318 15202 22370
rect 19406 22318 19458 22370
rect 20638 22318 20690 22370
rect 21758 22318 21810 22370
rect 22766 22318 22818 22370
rect 28254 22318 28306 22370
rect 28702 22318 28754 22370
rect 29150 22318 29202 22370
rect 37662 22318 37714 22370
rect 15486 22206 15538 22258
rect 15822 22206 15874 22258
rect 16494 22206 16546 22258
rect 16942 22206 16994 22258
rect 17390 22206 17442 22258
rect 28142 22206 28194 22258
rect 29934 22206 29986 22258
rect 14814 22094 14866 22146
rect 16270 22094 16322 22146
rect 16830 22094 16882 22146
rect 17726 22094 17778 22146
rect 19294 22094 19346 22146
rect 20414 22094 20466 22146
rect 21982 22094 22034 22146
rect 28030 22094 28082 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 15822 21758 15874 21810
rect 23102 21758 23154 21810
rect 25566 21758 25618 21810
rect 26238 21758 26290 21810
rect 29710 21758 29762 21810
rect 29934 21758 29986 21810
rect 13246 21646 13298 21698
rect 24222 21646 24274 21698
rect 26126 21646 26178 21698
rect 26350 21646 26402 21698
rect 27134 21646 27186 21698
rect 13918 21534 13970 21586
rect 15150 21534 15202 21586
rect 15598 21534 15650 21586
rect 22654 21534 22706 21586
rect 22878 21534 22930 21586
rect 23326 21534 23378 21586
rect 23550 21534 23602 21586
rect 23886 21534 23938 21586
rect 25454 21534 25506 21586
rect 26910 21534 26962 21586
rect 27582 21534 27634 21586
rect 30046 21534 30098 21586
rect 37662 21534 37714 21586
rect 11118 21422 11170 21474
rect 17614 21422 17666 21474
rect 27022 21422 27074 21474
rect 28814 21422 28866 21474
rect 40014 21422 40066 21474
rect 14254 21310 14306 21362
rect 14702 21310 14754 21362
rect 14926 21310 14978 21362
rect 25566 21310 25618 21362
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 16270 20974 16322 21026
rect 17950 20974 18002 21026
rect 18622 20974 18674 21026
rect 18286 20862 18338 20914
rect 20302 20862 20354 20914
rect 22430 20862 22482 20914
rect 40014 20862 40066 20914
rect 15710 20750 15762 20802
rect 16606 20750 16658 20802
rect 16830 20750 16882 20802
rect 17614 20750 17666 20802
rect 18958 20750 19010 20802
rect 19406 20750 19458 20802
rect 20078 20750 20130 20802
rect 20414 20750 20466 20802
rect 21982 20750 22034 20802
rect 22094 20750 22146 20802
rect 22318 20750 22370 20802
rect 22542 20750 22594 20802
rect 23326 20750 23378 20802
rect 29038 20750 29090 20802
rect 29374 20750 29426 20802
rect 37662 20750 37714 20802
rect 17166 20638 17218 20690
rect 18174 20638 18226 20690
rect 19182 20638 19234 20690
rect 21310 20638 21362 20690
rect 21646 20638 21698 20690
rect 22878 20638 22930 20690
rect 25454 20638 25506 20690
rect 14254 20526 14306 20578
rect 15934 20526 15986 20578
rect 17054 20526 17106 20578
rect 17390 20526 17442 20578
rect 21422 20526 21474 20578
rect 22990 20526 23042 20578
rect 29262 20526 29314 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 16494 20190 16546 20242
rect 18062 20190 18114 20242
rect 18398 20190 18450 20242
rect 25342 20190 25394 20242
rect 25566 20190 25618 20242
rect 25790 20190 25842 20242
rect 25902 20190 25954 20242
rect 13694 20078 13746 20130
rect 16718 20078 16770 20130
rect 17726 20078 17778 20130
rect 18734 20078 18786 20130
rect 18958 20078 19010 20130
rect 23326 20078 23378 20130
rect 27582 20078 27634 20130
rect 30046 20078 30098 20130
rect 30158 20078 30210 20130
rect 4286 19966 4338 20018
rect 13470 19966 13522 20018
rect 13806 19966 13858 20018
rect 17390 19966 17442 20018
rect 18846 19966 18898 20018
rect 19742 19966 19794 20018
rect 25230 19966 25282 20018
rect 26014 19966 26066 20018
rect 26350 19966 26402 20018
rect 26910 19966 26962 20018
rect 37662 19966 37714 20018
rect 13134 19854 13186 19906
rect 16606 19854 16658 19906
rect 29710 19854 29762 19906
rect 30718 19854 30770 19906
rect 1934 19742 1986 19794
rect 30158 19742 30210 19794
rect 40014 19742 40066 19794
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 15262 19406 15314 19458
rect 17614 19406 17666 19458
rect 23438 19406 23490 19458
rect 23774 19406 23826 19458
rect 9998 19294 10050 19346
rect 16046 19294 16098 19346
rect 17726 19294 17778 19346
rect 32062 19294 32114 19346
rect 12910 19182 12962 19234
rect 13470 19182 13522 19234
rect 13806 19182 13858 19234
rect 14030 19182 14082 19234
rect 15374 19182 15426 19234
rect 16270 19182 16322 19234
rect 20302 19182 20354 19234
rect 20526 19182 20578 19234
rect 20862 19182 20914 19234
rect 21198 19182 21250 19234
rect 21534 19182 21586 19234
rect 22430 19182 22482 19234
rect 22878 19182 22930 19234
rect 24110 19182 24162 19234
rect 25678 19182 25730 19234
rect 28702 19182 28754 19234
rect 29262 19182 29314 19234
rect 12126 19070 12178 19122
rect 13582 19070 13634 19122
rect 18286 19070 18338 19122
rect 18958 19070 19010 19122
rect 19070 19070 19122 19122
rect 19966 19070 20018 19122
rect 20078 19070 20130 19122
rect 20638 19070 20690 19122
rect 21758 19070 21810 19122
rect 22318 19070 22370 19122
rect 23662 19070 23714 19122
rect 24446 19070 24498 19122
rect 28142 19070 28194 19122
rect 29934 19070 29986 19122
rect 15262 18958 15314 19010
rect 16606 18958 16658 19010
rect 16942 18958 16994 19010
rect 17278 18958 17330 19010
rect 17950 18958 18002 19010
rect 18174 18958 18226 19010
rect 19294 18958 19346 19010
rect 19742 18958 19794 19010
rect 21870 18958 21922 19010
rect 24782 18958 24834 19010
rect 25118 18958 25170 19010
rect 25342 18958 25394 19010
rect 25566 18958 25618 19010
rect 28030 18958 28082 19010
rect 28254 18958 28306 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 16830 18622 16882 18674
rect 22766 18622 22818 18674
rect 24222 18622 24274 18674
rect 28814 18622 28866 18674
rect 13358 18510 13410 18562
rect 13470 18510 13522 18562
rect 18622 18510 18674 18562
rect 21758 18510 21810 18562
rect 22990 18510 23042 18562
rect 23886 18510 23938 18562
rect 23998 18510 24050 18562
rect 26238 18510 26290 18562
rect 27358 18510 27410 18562
rect 27470 18510 27522 18562
rect 4286 18398 4338 18450
rect 13694 18398 13746 18450
rect 13806 18398 13858 18450
rect 14142 18398 14194 18450
rect 16606 18398 16658 18450
rect 17726 18398 17778 18450
rect 17950 18398 18002 18450
rect 18398 18398 18450 18450
rect 21534 18398 21586 18450
rect 22542 18398 22594 18450
rect 23214 18398 23266 18450
rect 25790 18398 25842 18450
rect 26014 18398 26066 18450
rect 26462 18398 26514 18450
rect 27694 18398 27746 18450
rect 14590 18286 14642 18338
rect 15038 18286 15090 18338
rect 21982 18286 22034 18338
rect 25454 18286 25506 18338
rect 1934 18174 1986 18226
rect 14478 18174 14530 18226
rect 17390 18174 17442 18226
rect 22654 18174 22706 18226
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 15150 17838 15202 17890
rect 22430 17838 22482 17890
rect 9998 17726 10050 17778
rect 12126 17726 12178 17778
rect 22206 17726 22258 17778
rect 23662 17726 23714 17778
rect 27246 17726 27298 17778
rect 40014 17726 40066 17778
rect 12910 17614 12962 17666
rect 15486 17614 15538 17666
rect 15710 17614 15762 17666
rect 16382 17614 16434 17666
rect 17614 17614 17666 17666
rect 21422 17614 21474 17666
rect 23550 17614 23602 17666
rect 23998 17614 24050 17666
rect 24334 17614 24386 17666
rect 26126 17614 26178 17666
rect 26462 17614 26514 17666
rect 27582 17614 27634 17666
rect 28366 17614 28418 17666
rect 37662 17614 37714 17666
rect 21646 17502 21698 17554
rect 26798 17502 26850 17554
rect 26910 17502 26962 17554
rect 27918 17502 27970 17554
rect 13582 17390 13634 17442
rect 16046 17390 16098 17442
rect 17838 17390 17890 17442
rect 22766 17390 22818 17442
rect 23774 17390 23826 17442
rect 24894 17390 24946 17442
rect 25230 17390 25282 17442
rect 25790 17390 25842 17442
rect 26686 17390 26738 17442
rect 27694 17390 27746 17442
rect 27806 17390 27858 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 21758 17054 21810 17106
rect 26686 17054 26738 17106
rect 14478 16942 14530 16994
rect 27806 16942 27858 16994
rect 13806 16830 13858 16882
rect 17502 16830 17554 16882
rect 17838 16830 17890 16882
rect 21422 16830 21474 16882
rect 27022 16830 27074 16882
rect 37662 16830 37714 16882
rect 16606 16718 16658 16770
rect 18062 16718 18114 16770
rect 29934 16718 29986 16770
rect 40014 16718 40066 16770
rect 18174 16606 18226 16658
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 20414 16270 20466 16322
rect 21310 16270 21362 16322
rect 21646 16270 21698 16322
rect 27246 16158 27298 16210
rect 28142 16158 28194 16210
rect 18286 16046 18338 16098
rect 18958 16046 19010 16098
rect 19854 16046 19906 16098
rect 20078 16046 20130 16098
rect 20638 16046 20690 16098
rect 21310 16046 21362 16098
rect 22766 16046 22818 16098
rect 26910 16046 26962 16098
rect 27694 16046 27746 16098
rect 18510 15934 18562 15986
rect 27246 15934 27298 15986
rect 18622 15822 18674 15874
rect 19966 15822 20018 15874
rect 22430 15822 22482 15874
rect 27134 15822 27186 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 27022 15486 27074 15538
rect 19070 15374 19122 15426
rect 22318 15374 22370 15426
rect 26238 15374 26290 15426
rect 28702 15374 28754 15426
rect 18398 15262 18450 15314
rect 21646 15262 21698 15314
rect 25342 15262 25394 15314
rect 26350 15262 26402 15314
rect 26686 15262 26738 15314
rect 26910 15262 26962 15314
rect 27246 15262 27298 15314
rect 28030 15262 28082 15314
rect 21198 15150 21250 15202
rect 24446 15150 24498 15202
rect 30830 15150 30882 15202
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 18174 14590 18226 14642
rect 20302 14590 20354 14642
rect 20862 14590 20914 14642
rect 21422 14590 21474 14642
rect 26462 14590 26514 14642
rect 28590 14590 28642 14642
rect 29262 14590 29314 14642
rect 40014 14590 40066 14642
rect 17502 14478 17554 14530
rect 23886 14478 23938 14530
rect 24222 14478 24274 14530
rect 24558 14478 24610 14530
rect 25006 14478 25058 14530
rect 25342 14478 25394 14530
rect 25678 14478 25730 14530
rect 37662 14478 37714 14530
rect 24222 14254 24274 14306
rect 25230 14254 25282 14306
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 26462 13918 26514 13970
rect 27246 13918 27298 13970
rect 27470 13918 27522 13970
rect 26126 13806 26178 13858
rect 26798 13806 26850 13858
rect 27582 13806 27634 13858
rect 25790 13694 25842 13746
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 23774 13022 23826 13074
rect 25902 13022 25954 13074
rect 26462 13022 26514 13074
rect 22990 12910 23042 12962
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 25790 4286 25842 4338
rect 28702 4286 28754 4338
rect 26798 4062 26850 4114
rect 29710 4062 29762 4114
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 22430 3614 22482 3666
rect 25566 3614 25618 3666
rect 29374 3614 29426 3666
rect 21422 3502 21474 3554
rect 24558 3502 24610 3554
rect 28590 3502 28642 3554
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
<< metal2 >>
rect 18816 41200 18928 42000
rect 20160 41200 20272 42000
rect 22176 41200 22288 42000
rect 22848 41200 22960 42000
rect 23520 41200 23632 42000
rect 24192 41200 24304 42000
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 18844 38162 18900 41200
rect 18844 38110 18846 38162
rect 18898 38110 18900 38162
rect 18844 38098 18900 38110
rect 18060 38050 18116 38062
rect 18060 37998 18062 38050
rect 18114 37998 18116 38050
rect 18060 37044 18116 37998
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 20188 37492 20244 41200
rect 22204 38162 22260 41200
rect 22876 38276 22932 41200
rect 22876 38210 22932 38220
rect 22204 38110 22206 38162
rect 22258 38110 22260 38162
rect 22204 38098 22260 38110
rect 20188 37426 20244 37436
rect 21420 37492 21476 37502
rect 21420 37398 21476 37436
rect 20412 37266 20468 37278
rect 20412 37214 20414 37266
rect 20466 37214 20468 37266
rect 18060 36978 18116 36988
rect 18844 37044 18900 37054
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 17388 27858 17444 27870
rect 17388 27806 17390 27858
rect 17442 27806 17444 27858
rect 4172 27636 4228 27646
rect 1932 26066 1988 26078
rect 1932 26014 1934 26066
rect 1986 26014 1988 26066
rect 1932 25620 1988 26014
rect 1932 25554 1988 25564
rect 2044 25618 2100 25630
rect 2044 25566 2046 25618
rect 2098 25566 2100 25618
rect 2044 24948 2100 25566
rect 2044 24882 2100 24892
rect 1932 24050 1988 24062
rect 1932 23998 1934 24050
rect 1986 23998 1988 24050
rect 1932 23604 1988 23998
rect 1932 23538 1988 23548
rect 1932 19796 1988 19806
rect 1932 19702 1988 19740
rect 4172 19012 4228 27580
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 16044 27076 16100 27086
rect 4284 26292 4340 26302
rect 4284 26198 4340 26236
rect 12796 26292 12852 26302
rect 12796 26178 12852 26236
rect 15708 26292 15764 26302
rect 15708 26290 15876 26292
rect 15708 26238 15710 26290
rect 15762 26238 15876 26290
rect 15708 26236 15876 26238
rect 15708 26226 15764 26236
rect 12796 26126 12798 26178
rect 12850 26126 12852 26178
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 4284 25506 4340 25518
rect 4284 25454 4286 25506
rect 4338 25454 4340 25506
rect 4284 25284 4340 25454
rect 12796 25396 12852 26126
rect 14924 26180 14980 26190
rect 15820 26180 15876 26236
rect 16044 26180 16100 27020
rect 17388 27076 17444 27806
rect 18172 27748 18228 27758
rect 18172 27654 18228 27692
rect 18844 27188 18900 36988
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 20412 31948 20468 37214
rect 23548 36708 23604 41200
rect 23996 38052 24052 38062
rect 23996 38050 24164 38052
rect 23996 37998 23998 38050
rect 24050 37998 24164 38050
rect 23996 37996 24164 37998
rect 23996 37986 24052 37996
rect 23548 36642 23604 36652
rect 23772 36482 23828 36494
rect 23772 36430 23774 36482
rect 23826 36430 23828 36482
rect 23772 31948 23828 36430
rect 20300 31892 20468 31948
rect 23660 31892 23828 31948
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 20076 27748 20132 27758
rect 20076 27298 20132 27692
rect 20076 27246 20078 27298
rect 20130 27246 20132 27298
rect 20076 27234 20132 27246
rect 20300 27746 20356 31892
rect 23436 28642 23492 28654
rect 23436 28590 23438 28642
rect 23490 28590 23492 28642
rect 23436 28532 23492 28590
rect 21308 27858 21364 27870
rect 21308 27806 21310 27858
rect 21362 27806 21364 27858
rect 20300 27694 20302 27746
rect 20354 27694 20356 27746
rect 17388 27010 17444 27020
rect 18620 27186 18900 27188
rect 18620 27134 18846 27186
rect 18898 27134 18900 27186
rect 18620 27132 18900 27134
rect 16716 26962 16772 26974
rect 16716 26910 16718 26962
rect 16770 26910 16772 26962
rect 16156 26180 16212 26190
rect 14924 26178 15204 26180
rect 14924 26126 14926 26178
rect 14978 26126 15204 26178
rect 14924 26124 15204 26126
rect 14924 26114 14980 26124
rect 12796 25330 12852 25340
rect 14252 25620 14308 25630
rect 14252 25394 14308 25564
rect 14252 25342 14254 25394
rect 14306 25342 14308 25394
rect 4284 25218 4340 25228
rect 11564 25284 11620 25294
rect 11564 24610 11620 25228
rect 13692 24836 13748 24846
rect 13692 24742 13748 24780
rect 11564 24558 11566 24610
rect 11618 24558 11620 24610
rect 11564 24546 11620 24558
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 9996 24050 10052 24062
rect 9996 23998 9998 24050
rect 10050 23998 10052 24050
rect 4284 23940 4340 23950
rect 4284 23846 4340 23884
rect 9996 23716 10052 23998
rect 12124 24052 12180 24062
rect 12124 23958 12180 23996
rect 13580 24052 13636 24062
rect 13580 23958 13636 23996
rect 9996 23650 10052 23660
rect 12908 23940 12964 23950
rect 12908 23044 12964 23884
rect 13804 23828 13860 23838
rect 13804 23734 13860 23772
rect 13580 23714 13636 23726
rect 13580 23662 13582 23714
rect 13634 23662 13636 23714
rect 13580 23380 13636 23662
rect 13580 23314 13636 23324
rect 14028 23716 14084 23726
rect 14028 23266 14084 23660
rect 14028 23214 14030 23266
rect 14082 23214 14084 23266
rect 14028 23202 14084 23214
rect 14252 23154 14308 25342
rect 15036 25506 15092 25518
rect 15036 25454 15038 25506
rect 15090 25454 15092 25506
rect 14364 25284 14420 25294
rect 14364 25190 14420 25228
rect 14588 25284 14644 25294
rect 14588 25282 14868 25284
rect 14588 25230 14590 25282
rect 14642 25230 14868 25282
rect 14588 25228 14868 25230
rect 14588 25218 14644 25228
rect 14476 25172 14532 25182
rect 14364 24724 14420 24734
rect 14476 24724 14532 25116
rect 14812 25060 14868 25228
rect 15036 25172 15092 25454
rect 15148 25284 15204 26124
rect 15820 26178 16212 26180
rect 15820 26126 16158 26178
rect 16210 26126 16212 26178
rect 15820 26124 16212 26126
rect 15260 25564 15764 25620
rect 15260 25506 15316 25564
rect 15260 25454 15262 25506
rect 15314 25454 15316 25506
rect 15260 25442 15316 25454
rect 15708 25506 15764 25564
rect 15708 25454 15710 25506
rect 15762 25454 15764 25506
rect 15708 25442 15764 25454
rect 15484 25394 15540 25406
rect 15484 25342 15486 25394
rect 15538 25342 15540 25394
rect 15260 25284 15316 25294
rect 15148 25282 15316 25284
rect 15148 25230 15262 25282
rect 15314 25230 15316 25282
rect 15148 25228 15316 25230
rect 15260 25218 15316 25228
rect 15036 25116 15204 25172
rect 14812 25004 15092 25060
rect 14924 24836 14980 24846
rect 14924 24742 14980 24780
rect 14364 24722 14532 24724
rect 14364 24670 14366 24722
rect 14418 24670 14532 24722
rect 14364 24668 14532 24670
rect 14812 24722 14868 24734
rect 14812 24670 14814 24722
rect 14866 24670 14868 24722
rect 14364 23940 14420 24668
rect 14364 23874 14420 23884
rect 14700 23940 14756 23950
rect 14700 23846 14756 23884
rect 14364 23380 14420 23390
rect 14364 23286 14420 23324
rect 14252 23102 14254 23154
rect 14306 23102 14308 23154
rect 13132 23044 13188 23054
rect 12908 23042 13188 23044
rect 12908 22990 13134 23042
rect 13186 22990 13188 23042
rect 12908 22988 13188 22990
rect 13132 22932 13188 22988
rect 13132 22876 13524 22932
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 13244 22148 13300 22158
rect 13244 21698 13300 22092
rect 13244 21646 13246 21698
rect 13298 21646 13300 21698
rect 13244 21634 13300 21646
rect 11116 21476 11172 21486
rect 11116 21382 11172 21420
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 13468 20580 13524 22876
rect 14252 22484 14308 23102
rect 14252 22418 14308 22428
rect 14476 23154 14532 23166
rect 14476 23102 14478 23154
rect 14530 23102 14532 23154
rect 14476 22372 14532 23102
rect 14700 23156 14756 23166
rect 14476 22306 14532 22316
rect 14588 22372 14644 22382
rect 14700 22372 14756 23100
rect 14588 22370 14756 22372
rect 14588 22318 14590 22370
rect 14642 22318 14756 22370
rect 14588 22316 14756 22318
rect 14588 22306 14644 22316
rect 14812 22146 14868 24670
rect 15036 24722 15092 25004
rect 15036 24670 15038 24722
rect 15090 24670 15092 24722
rect 15036 24658 15092 24670
rect 15148 24724 15204 25116
rect 15484 24836 15540 25342
rect 15820 25284 15876 26124
rect 16156 26114 16212 26124
rect 16716 26180 16772 26910
rect 18620 26514 18676 27132
rect 18844 27122 18900 27132
rect 19740 27076 19796 27086
rect 19740 27074 20132 27076
rect 19740 27022 19742 27074
rect 19794 27022 20132 27074
rect 19740 27020 20132 27022
rect 19740 27010 19796 27020
rect 19404 26962 19460 26974
rect 19404 26910 19406 26962
rect 19458 26910 19460 26962
rect 19404 26908 19460 26910
rect 18620 26462 18622 26514
rect 18674 26462 18676 26514
rect 18620 26450 18676 26462
rect 18732 26852 19460 26908
rect 19516 26964 19572 26974
rect 19516 26870 19572 26908
rect 20076 26962 20132 27020
rect 20076 26910 20078 26962
rect 20130 26910 20132 26962
rect 20076 26898 20132 26910
rect 20188 26962 20244 26974
rect 20188 26910 20190 26962
rect 20242 26910 20244 26962
rect 17500 26404 17556 26414
rect 17500 26310 17556 26348
rect 18396 26404 18452 26414
rect 18396 26310 18452 26348
rect 18732 26402 18788 26852
rect 19404 26786 19460 26796
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 18732 26350 18734 26402
rect 18786 26350 18788 26402
rect 18732 26338 18788 26350
rect 16716 26114 16772 26124
rect 17388 26290 17444 26302
rect 17388 26238 17390 26290
rect 17442 26238 17444 26290
rect 16044 25508 16100 25518
rect 16044 25414 16100 25452
rect 15932 25396 15988 25406
rect 15932 25302 15988 25340
rect 15820 25218 15876 25228
rect 15596 24836 15652 24846
rect 15484 24780 15596 24836
rect 15260 24724 15316 24734
rect 15148 24722 15316 24724
rect 15148 24670 15262 24722
rect 15314 24670 15316 24722
rect 15148 24668 15316 24670
rect 15148 24052 15204 24668
rect 15260 24658 15316 24668
rect 15036 23996 15204 24052
rect 15036 23828 15092 23996
rect 14924 22372 14980 22382
rect 14924 22278 14980 22316
rect 15036 22148 15092 23772
rect 15596 23378 15652 24780
rect 15596 23326 15598 23378
rect 15650 23326 15652 23378
rect 15596 23314 15652 23326
rect 16716 24612 16772 24622
rect 16716 23378 16772 24556
rect 17388 24612 17444 26238
rect 17500 26180 17556 26190
rect 17500 26066 17556 26124
rect 17500 26014 17502 26066
rect 17554 26014 17556 26066
rect 17500 26002 17556 26014
rect 19180 26180 19236 26190
rect 18844 25508 18900 25518
rect 18060 25284 18116 25294
rect 18060 24722 18116 25228
rect 18844 24834 18900 25452
rect 19180 25284 19236 26124
rect 20076 26180 20132 26190
rect 20076 26086 20132 26124
rect 19628 25844 19684 25854
rect 19180 25218 19236 25228
rect 19516 25788 19628 25844
rect 18844 24782 18846 24834
rect 18898 24782 18900 24834
rect 18844 24770 18900 24782
rect 18060 24670 18062 24722
rect 18114 24670 18116 24722
rect 18060 24658 18116 24670
rect 17388 24546 17444 24556
rect 19516 23828 19572 25788
rect 19628 25778 19684 25788
rect 20188 25844 20244 26910
rect 20300 26964 20356 27694
rect 20300 26898 20356 26908
rect 20860 27746 20916 27758
rect 20860 27694 20862 27746
rect 20914 27694 20916 27746
rect 20412 26292 20468 26302
rect 20860 26292 20916 27694
rect 21308 26852 21364 27806
rect 21980 27748 22036 27758
rect 21644 27746 22036 27748
rect 21644 27694 21982 27746
rect 22034 27694 22036 27746
rect 21644 27692 22036 27694
rect 21644 27298 21700 27692
rect 21980 27682 22036 27692
rect 21644 27246 21646 27298
rect 21698 27246 21700 27298
rect 21644 27234 21700 27246
rect 22540 27076 22596 27086
rect 21756 26964 21812 26974
rect 22316 26964 22372 26974
rect 21756 26962 22372 26964
rect 21756 26910 21758 26962
rect 21810 26910 22318 26962
rect 22370 26910 22372 26962
rect 21756 26908 22372 26910
rect 21756 26898 21812 26908
rect 22316 26898 22372 26908
rect 22540 26962 22596 27020
rect 23436 27076 23492 28476
rect 23660 28530 23716 31892
rect 23660 28478 23662 28530
rect 23714 28478 23716 28530
rect 23660 28466 23716 28478
rect 24108 28532 24164 37996
rect 24220 37492 24276 41200
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 25564 38276 25620 38286
rect 25564 38182 25620 38220
rect 24220 37426 24276 37436
rect 24556 38050 24612 38062
rect 24556 37998 24558 38050
rect 24610 37998 24612 38050
rect 24108 27746 24164 28476
rect 24108 27694 24110 27746
rect 24162 27694 24164 27746
rect 24108 27682 24164 27694
rect 23436 26982 23492 27020
rect 22540 26910 22542 26962
rect 22594 26910 22596 26962
rect 22540 26898 22596 26910
rect 22652 26962 22708 26974
rect 22652 26910 22654 26962
rect 22706 26910 22708 26962
rect 21644 26852 21700 26862
rect 21308 26786 21364 26796
rect 21532 26850 21700 26852
rect 21532 26798 21646 26850
rect 21698 26798 21700 26850
rect 21532 26796 21700 26798
rect 20412 26290 20916 26292
rect 20412 26238 20414 26290
rect 20466 26238 20916 26290
rect 20412 26236 20916 26238
rect 20412 26180 20468 26236
rect 20412 26114 20468 26124
rect 20860 25956 20916 26236
rect 21196 26180 21252 26190
rect 21196 26178 21364 26180
rect 21196 26126 21198 26178
rect 21250 26126 21364 26178
rect 21196 26124 21364 26126
rect 21196 26114 21252 26124
rect 20860 25890 20916 25900
rect 21196 25956 21252 25966
rect 20188 25778 20244 25788
rect 19628 25508 19684 25518
rect 19628 24162 19684 25452
rect 20748 25284 20804 25294
rect 20860 25284 20916 25294
rect 20748 25282 20860 25284
rect 20748 25230 20750 25282
rect 20802 25230 20860 25282
rect 20748 25228 20860 25230
rect 20748 25218 20804 25228
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 19628 24110 19630 24162
rect 19682 24110 19684 24162
rect 19628 24098 19684 24110
rect 19628 23828 19684 23838
rect 16716 23326 16718 23378
rect 16770 23326 16772 23378
rect 16716 23314 16772 23326
rect 19292 23826 19684 23828
rect 19292 23774 19630 23826
rect 19682 23774 19684 23826
rect 19292 23772 19684 23774
rect 15932 23266 15988 23278
rect 15932 23214 15934 23266
rect 15986 23214 15988 23266
rect 15484 23156 15540 23166
rect 14812 22094 14814 22146
rect 14866 22094 14868 22146
rect 14812 22082 14868 22094
rect 14924 22092 15092 22148
rect 15148 23154 15540 23156
rect 15148 23102 15486 23154
rect 15538 23102 15540 23154
rect 15148 23100 15540 23102
rect 15148 22370 15204 23100
rect 15484 23090 15540 23100
rect 15708 23156 15764 23166
rect 15148 22318 15150 22370
rect 15202 22318 15204 22370
rect 14700 21812 14756 21822
rect 13468 20188 13524 20524
rect 13916 21588 13972 21598
rect 13916 20580 13972 21532
rect 14252 21364 14308 21374
rect 14252 21362 14420 21364
rect 14252 21310 14254 21362
rect 14306 21310 14420 21362
rect 14252 21308 14420 21310
rect 14252 21298 14308 21308
rect 13916 20514 13972 20524
rect 14252 20580 14308 20590
rect 14252 20486 14308 20524
rect 14364 20188 14420 21308
rect 14700 21362 14756 21756
rect 14700 21310 14702 21362
rect 14754 21310 14756 21362
rect 14700 21028 14756 21310
rect 14924 21364 14980 22092
rect 15148 21812 15204 22318
rect 15484 22260 15540 22270
rect 15708 22260 15764 23100
rect 15148 21746 15204 21756
rect 15260 22258 15764 22260
rect 15260 22206 15486 22258
rect 15538 22206 15764 22258
rect 15260 22204 15764 22206
rect 15820 22258 15876 22270
rect 15820 22206 15822 22258
rect 15874 22206 15876 22258
rect 15148 21588 15204 21598
rect 15260 21588 15316 22204
rect 15484 22194 15540 22204
rect 15820 22036 15876 22206
rect 15708 21980 15876 22036
rect 15932 22260 15988 23214
rect 16492 23266 16548 23278
rect 16492 23214 16494 23266
rect 16546 23214 16548 23266
rect 16380 23156 16436 23166
rect 15708 21812 15764 21980
rect 15708 21746 15764 21756
rect 15820 21812 15876 21822
rect 15932 21812 15988 22204
rect 15820 21810 15988 21812
rect 15820 21758 15822 21810
rect 15874 21758 15988 21810
rect 15820 21756 15988 21758
rect 16044 23154 16436 23156
rect 16044 23102 16382 23154
rect 16434 23102 16436 23154
rect 16044 23100 16436 23102
rect 15820 21746 15876 21756
rect 15148 21586 15316 21588
rect 15148 21534 15150 21586
rect 15202 21534 15316 21586
rect 15148 21532 15316 21534
rect 15596 21588 15652 21598
rect 16044 21588 16100 23100
rect 16380 23090 16436 23100
rect 16156 22484 16212 22494
rect 16492 22484 16548 23214
rect 19292 22596 19348 23772
rect 19628 23762 19684 23772
rect 19740 23828 19796 23838
rect 19740 23826 20132 23828
rect 19740 23774 19742 23826
rect 19794 23774 20132 23826
rect 19740 23772 20132 23774
rect 19740 23762 19796 23772
rect 20076 23716 20132 23772
rect 20076 23660 20244 23716
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 19292 22594 19572 22596
rect 19292 22542 19294 22594
rect 19346 22542 19572 22594
rect 19292 22540 19572 22542
rect 19292 22530 19348 22540
rect 16156 22390 16212 22428
rect 16380 22428 16548 22484
rect 16268 22146 16324 22158
rect 16268 22094 16270 22146
rect 16322 22094 16324 22146
rect 16268 21812 16324 22094
rect 16380 22148 16436 22428
rect 17388 22372 17444 22382
rect 19404 22372 19460 22382
rect 16380 22082 16436 22092
rect 16492 22258 16548 22270
rect 16492 22206 16494 22258
rect 16546 22206 16548 22258
rect 16268 21746 16324 21756
rect 15596 21586 15764 21588
rect 15596 21534 15598 21586
rect 15650 21534 15764 21586
rect 15596 21532 15764 21534
rect 16044 21532 16324 21588
rect 15148 21522 15204 21532
rect 15596 21522 15652 21532
rect 14924 21270 14980 21308
rect 15708 21476 15764 21532
rect 14700 20962 14756 20972
rect 9996 20132 10052 20142
rect 4284 20020 4340 20030
rect 4284 19926 4340 19964
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 9996 19346 10052 20076
rect 9996 19294 9998 19346
rect 10050 19294 10052 19346
rect 9996 19282 10052 19294
rect 13132 20132 13524 20188
rect 13692 20132 13748 20142
rect 13132 19906 13188 20132
rect 13692 20038 13748 20076
rect 14028 20132 14420 20188
rect 15708 20802 15764 21420
rect 16268 21028 16324 21532
rect 16268 20934 16324 20972
rect 16492 20916 16548 22206
rect 16940 22260 16996 22270
rect 16996 22204 17220 22260
rect 16940 22166 16996 22204
rect 16828 22148 16884 22158
rect 16828 22054 16884 22092
rect 15708 20750 15710 20802
rect 15762 20750 15764 20802
rect 13132 19854 13134 19906
rect 13186 19854 13188 19906
rect 12908 19236 12964 19246
rect 13132 19236 13188 19854
rect 13468 20018 13524 20030
rect 13468 19966 13470 20018
rect 13522 19966 13524 20018
rect 12908 19234 13188 19236
rect 12908 19182 12910 19234
rect 12962 19182 13188 19234
rect 12908 19180 13188 19182
rect 13356 19460 13412 19470
rect 12124 19124 12180 19134
rect 12124 19030 12180 19068
rect 4172 18946 4228 18956
rect 12124 18564 12180 18574
rect 4284 18452 4340 18462
rect 4284 18358 4340 18396
rect 9996 18340 10052 18350
rect 1932 18228 1988 18238
rect 1932 18134 1988 18172
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 9996 17778 10052 18284
rect 9996 17726 9998 17778
rect 10050 17726 10052 17778
rect 9996 17714 10052 17726
rect 12124 17778 12180 18508
rect 12124 17726 12126 17778
rect 12178 17726 12180 17778
rect 12124 17714 12180 17726
rect 12908 17668 12964 19180
rect 13356 18562 13412 19404
rect 13468 19234 13524 19966
rect 13804 20018 13860 20030
rect 13804 19966 13806 20018
rect 13858 19966 13860 20018
rect 13804 19460 13860 19966
rect 13804 19394 13860 19404
rect 13468 19182 13470 19234
rect 13522 19182 13524 19234
rect 13468 19170 13524 19182
rect 13804 19236 13860 19246
rect 14028 19236 14084 20132
rect 15260 19460 15316 19470
rect 15260 19366 15316 19404
rect 15708 19348 15764 20750
rect 16380 20860 16548 20916
rect 15932 20580 15988 20590
rect 15932 20486 15988 20524
rect 16380 20132 16436 20860
rect 16604 20804 16660 20814
rect 16604 20710 16660 20748
rect 16828 20802 16884 20814
rect 16828 20750 16830 20802
rect 16882 20750 16884 20802
rect 16492 20692 16548 20702
rect 16492 20242 16548 20636
rect 16492 20190 16494 20242
rect 16546 20190 16548 20242
rect 16492 20178 16548 20190
rect 16380 20066 16436 20076
rect 16716 20132 16772 20142
rect 16828 20132 16884 20750
rect 17164 20692 17220 22204
rect 17388 22258 17444 22316
rect 17388 22206 17390 22258
rect 17442 22206 17444 22258
rect 17388 22194 17444 22206
rect 19180 22370 19460 22372
rect 19180 22318 19406 22370
rect 19458 22318 19460 22370
rect 19180 22316 19460 22318
rect 17724 22148 17780 22158
rect 17780 22092 18004 22148
rect 17724 22054 17780 22092
rect 17612 21476 17668 21486
rect 17612 21382 17668 21420
rect 17948 21028 18004 22092
rect 18396 21588 18452 21598
rect 17948 21026 18116 21028
rect 17948 20974 17950 21026
rect 18002 20974 18116 21026
rect 17948 20972 18116 20974
rect 17948 20962 18004 20972
rect 17164 20598 17220 20636
rect 17276 20804 17332 20814
rect 17612 20804 17668 20814
rect 17332 20802 17668 20804
rect 17332 20750 17614 20802
rect 17666 20750 17668 20802
rect 17332 20748 17668 20750
rect 16716 20130 16884 20132
rect 16716 20078 16718 20130
rect 16770 20078 16884 20130
rect 16716 20076 16884 20078
rect 16716 20066 16772 20076
rect 16604 19906 16660 19918
rect 16604 19854 16606 19906
rect 16658 19854 16660 19906
rect 16044 19348 16100 19358
rect 15708 19346 16100 19348
rect 15708 19294 16046 19346
rect 16098 19294 16100 19346
rect 15708 19292 16100 19294
rect 16044 19282 16100 19292
rect 13804 19142 13860 19180
rect 13916 19234 14084 19236
rect 13916 19182 14030 19234
rect 14082 19182 14084 19234
rect 13916 19180 14084 19182
rect 13580 19124 13636 19134
rect 13580 19030 13636 19068
rect 13916 18900 13972 19180
rect 14028 19170 14084 19180
rect 15372 19236 15428 19246
rect 15372 19142 15428 19180
rect 16268 19234 16324 19246
rect 16268 19182 16270 19234
rect 16322 19182 16324 19234
rect 13804 18844 13972 18900
rect 15260 19010 15316 19022
rect 15260 18958 15262 19010
rect 15314 18958 15316 19010
rect 13356 18510 13358 18562
rect 13410 18510 13412 18562
rect 13356 18498 13412 18510
rect 13468 18564 13524 18574
rect 13468 18470 13524 18508
rect 13692 18450 13748 18462
rect 13692 18398 13694 18450
rect 13746 18398 13748 18450
rect 13692 18004 13748 18398
rect 13804 18450 13860 18844
rect 13804 18398 13806 18450
rect 13858 18398 13860 18450
rect 13804 18386 13860 18398
rect 14140 18452 14196 18462
rect 14140 18358 14196 18396
rect 15036 18452 15092 18462
rect 14588 18340 14644 18350
rect 14588 18246 14644 18284
rect 15036 18338 15092 18396
rect 15036 18286 15038 18338
rect 15090 18286 15092 18338
rect 14476 18228 14532 18238
rect 13916 18226 14532 18228
rect 13916 18174 14478 18226
rect 14530 18174 14532 18226
rect 13916 18172 14532 18174
rect 13916 18004 13972 18172
rect 14476 18162 14532 18172
rect 15036 18116 15092 18286
rect 15148 18116 15204 18126
rect 15036 18060 15148 18116
rect 13692 17948 13972 18004
rect 15148 17890 15204 18060
rect 15148 17838 15150 17890
rect 15202 17838 15204 17890
rect 15148 17826 15204 17838
rect 12908 17574 12964 17612
rect 13580 17668 13636 17678
rect 13580 17442 13636 17612
rect 15260 17668 15316 18958
rect 16268 18452 16324 19182
rect 16604 19236 16660 19854
rect 16604 19170 16660 19180
rect 16828 19348 16884 20076
rect 16604 19010 16660 19022
rect 16604 18958 16606 19010
rect 16658 18958 16660 19010
rect 16604 18676 16660 18958
rect 16604 18610 16660 18620
rect 16828 18674 16884 19292
rect 17052 20578 17108 20590
rect 17052 20526 17054 20578
rect 17106 20526 17108 20578
rect 17052 19124 17108 20526
rect 17276 20020 17332 20748
rect 17612 20738 17668 20748
rect 17388 20580 17444 20590
rect 18060 20580 18116 20972
rect 18284 20916 18340 20926
rect 18284 20822 18340 20860
rect 18172 20804 18228 20814
rect 18172 20690 18228 20748
rect 18172 20638 18174 20690
rect 18226 20638 18228 20690
rect 18172 20626 18228 20638
rect 17388 20578 17556 20580
rect 17388 20526 17390 20578
rect 17442 20526 17556 20578
rect 17388 20524 17556 20526
rect 17388 20514 17444 20524
rect 17500 20356 17556 20524
rect 18060 20468 18116 20524
rect 18060 20412 18228 20468
rect 17500 20300 18116 20356
rect 17388 20020 17444 20030
rect 17276 19964 17388 20020
rect 17388 19926 17444 19964
rect 17612 19458 17668 20300
rect 18060 20242 18116 20300
rect 18060 20190 18062 20242
rect 18114 20190 18116 20242
rect 18060 20178 18116 20190
rect 17724 20132 17780 20142
rect 17780 20076 17892 20132
rect 17724 20038 17780 20076
rect 17612 19406 17614 19458
rect 17666 19406 17668 19458
rect 17612 19394 17668 19406
rect 17724 19348 17780 19358
rect 17724 19254 17780 19292
rect 17836 19124 17892 20076
rect 18172 19908 18228 20412
rect 18396 20242 18452 21532
rect 18620 21364 18676 21374
rect 18620 21026 18676 21308
rect 18620 20974 18622 21026
rect 18674 20974 18676 21026
rect 18620 20962 18676 20974
rect 18396 20190 18398 20242
rect 18450 20190 18452 20242
rect 18396 20178 18452 20190
rect 18732 20804 18788 20814
rect 18732 20130 18788 20748
rect 18956 20802 19012 20814
rect 18956 20750 18958 20802
rect 19010 20750 19012 20802
rect 18956 20468 19012 20750
rect 19180 20692 19236 22316
rect 19404 22306 19460 22316
rect 19292 22148 19348 22158
rect 19292 22054 19348 22092
rect 19404 21812 19460 21822
rect 19404 20802 19460 21756
rect 19404 20750 19406 20802
rect 19458 20750 19460 20802
rect 19404 20738 19460 20750
rect 19180 20690 19348 20692
rect 19180 20638 19182 20690
rect 19234 20638 19348 20690
rect 19180 20636 19348 20638
rect 19180 20626 19236 20636
rect 18956 20402 19012 20412
rect 18732 20078 18734 20130
rect 18786 20078 18788 20130
rect 18732 20066 18788 20078
rect 18956 20132 19012 20142
rect 18956 20038 19012 20076
rect 18844 20020 18900 20030
rect 18844 19926 18900 19964
rect 17052 19058 17108 19068
rect 17500 19068 17892 19124
rect 18060 19852 18228 19908
rect 16828 18622 16830 18674
rect 16882 18622 16884 18674
rect 16828 18610 16884 18622
rect 16940 19010 16996 19022
rect 16940 18958 16942 19010
rect 16994 18958 16996 19010
rect 16604 18452 16660 18462
rect 16268 18450 16660 18452
rect 16268 18398 16606 18450
rect 16658 18398 16660 18450
rect 16268 18396 16660 18398
rect 16604 18340 16660 18396
rect 16940 18340 16996 18958
rect 17276 19010 17332 19022
rect 17276 18958 17278 19010
rect 17330 18958 17332 19010
rect 17276 18900 17332 18958
rect 17276 18834 17332 18844
rect 16604 18284 16996 18340
rect 16380 18228 16436 18238
rect 15260 17602 15316 17612
rect 15484 17666 15540 17678
rect 15484 17614 15486 17666
rect 15538 17614 15540 17666
rect 13580 17390 13582 17442
rect 13634 17390 13636 17442
rect 13580 16884 13636 17390
rect 15484 17444 15540 17614
rect 15708 17668 15764 17678
rect 15708 17574 15764 17612
rect 16380 17666 16436 18172
rect 16380 17614 16382 17666
rect 16434 17614 16436 17666
rect 16380 17602 16436 17614
rect 16044 17444 16100 17454
rect 15484 17442 16100 17444
rect 15484 17390 16046 17442
rect 16098 17390 16100 17442
rect 15484 17388 16100 17390
rect 14476 16996 14532 17006
rect 14476 16902 14532 16940
rect 15484 16996 15540 17388
rect 16044 17378 16100 17388
rect 15484 16930 15540 16940
rect 13804 16884 13860 16894
rect 13580 16828 13804 16884
rect 13804 16790 13860 16828
rect 16604 16770 16660 18284
rect 17388 18228 17444 18238
rect 17388 18134 17444 18172
rect 17500 17444 17556 19068
rect 17948 19012 18004 19022
rect 17836 19010 18004 19012
rect 17836 18958 17950 19010
rect 18002 18958 18004 19010
rect 17836 18956 18004 18958
rect 18060 19012 18116 19852
rect 18284 19684 18340 19694
rect 18284 19122 18340 19628
rect 19292 19460 19348 20636
rect 19404 20468 19460 20478
rect 19404 19796 19460 20412
rect 19404 19730 19460 19740
rect 19404 19460 19460 19470
rect 19292 19404 19404 19460
rect 19404 19394 19460 19404
rect 18284 19070 18286 19122
rect 18338 19070 18340 19122
rect 18172 19012 18228 19022
rect 18060 19010 18228 19012
rect 18060 18958 18174 19010
rect 18226 18958 18228 19010
rect 18060 18956 18228 18958
rect 17724 18452 17780 18462
rect 17836 18452 17892 18956
rect 17948 18946 18004 18956
rect 18172 18946 18228 18956
rect 18284 18900 18340 19070
rect 18284 18834 18340 18844
rect 18396 19348 18452 19358
rect 17724 18450 17892 18452
rect 17724 18398 17726 18450
rect 17778 18398 17892 18450
rect 17724 18396 17892 18398
rect 17948 18676 18004 18686
rect 17948 18450 18004 18620
rect 17948 18398 17950 18450
rect 18002 18398 18004 18450
rect 17612 17668 17668 17678
rect 17724 17668 17780 18396
rect 17948 18386 18004 18398
rect 18396 18450 18452 19292
rect 19516 19236 19572 22540
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 20076 20802 20132 20814
rect 20076 20750 20078 20802
rect 20130 20750 20132 20802
rect 20076 20580 20132 20750
rect 20076 20514 20132 20524
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 19068 19180 19572 19236
rect 19740 20018 19796 20030
rect 19740 19966 19742 20018
rect 19794 19966 19796 20018
rect 18956 19124 19012 19134
rect 18956 19030 19012 19068
rect 19068 19122 19124 19180
rect 19068 19070 19070 19122
rect 19122 19070 19124 19122
rect 19068 19058 19124 19070
rect 19628 19124 19684 19134
rect 19292 19010 19348 19022
rect 19292 18958 19294 19010
rect 19346 18958 19348 19010
rect 18396 18398 18398 18450
rect 18450 18398 18452 18450
rect 18396 18386 18452 18398
rect 18620 18562 18676 18574
rect 18620 18510 18622 18562
rect 18674 18510 18676 18562
rect 18620 18228 18676 18510
rect 18620 18162 18676 18172
rect 19292 17780 19348 18958
rect 19292 17714 19348 17724
rect 17612 17666 17780 17668
rect 17612 17614 17614 17666
rect 17666 17614 17780 17666
rect 17612 17612 17780 17614
rect 17612 17602 17668 17612
rect 17724 17444 17780 17454
rect 17500 17388 17724 17444
rect 16604 16718 16606 16770
rect 16658 16718 16660 16770
rect 16604 16706 16660 16718
rect 17500 16884 17556 16894
rect 17724 16884 17780 17388
rect 17836 17442 17892 17454
rect 17836 17390 17838 17442
rect 17890 17390 17892 17442
rect 17836 17220 17892 17390
rect 17836 17164 18228 17220
rect 17836 16884 17892 16894
rect 17724 16882 17892 16884
rect 17724 16830 17838 16882
rect 17890 16830 17892 16882
rect 17724 16828 17892 16830
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 17500 14644 17556 16828
rect 17836 16818 17892 16828
rect 18060 16770 18116 16782
rect 18060 16718 18062 16770
rect 18114 16718 18116 16770
rect 18060 16100 18116 16718
rect 18172 16660 18228 17164
rect 19628 16772 19684 19068
rect 19740 19012 19796 19966
rect 20076 19908 20132 19918
rect 19964 19124 20020 19134
rect 19964 19030 20020 19068
rect 20076 19122 20132 19852
rect 20188 19236 20244 23660
rect 20748 23380 20804 23418
rect 20748 23314 20804 23324
rect 20412 23268 20468 23278
rect 20412 23266 20692 23268
rect 20412 23214 20414 23266
rect 20466 23214 20692 23266
rect 20412 23212 20692 23214
rect 20412 23202 20468 23212
rect 20636 22372 20692 23212
rect 20860 23156 20916 25228
rect 21196 24948 21252 25900
rect 21308 25282 21364 26124
rect 21308 25230 21310 25282
rect 21362 25230 21364 25282
rect 21308 25218 21364 25230
rect 21420 25506 21476 25518
rect 21420 25454 21422 25506
rect 21474 25454 21476 25506
rect 21420 25284 21476 25454
rect 21420 25218 21476 25228
rect 21420 24948 21476 24958
rect 21196 24946 21476 24948
rect 21196 24894 21422 24946
rect 21474 24894 21476 24946
rect 21196 24892 21476 24894
rect 21420 24882 21476 24892
rect 20972 24610 21028 24622
rect 20972 24558 20974 24610
rect 21026 24558 21028 24610
rect 20972 23380 21028 24558
rect 21028 23324 21252 23380
rect 20972 23314 21028 23324
rect 21196 23266 21252 23324
rect 21196 23214 21198 23266
rect 21250 23214 21252 23266
rect 21196 23202 21252 23214
rect 20300 22370 20692 22372
rect 20300 22318 20638 22370
rect 20690 22318 20692 22370
rect 20300 22316 20692 22318
rect 20300 21364 20356 22316
rect 20636 22306 20692 22316
rect 20748 23100 20916 23156
rect 20412 22148 20468 22158
rect 20412 22146 20692 22148
rect 20412 22094 20414 22146
rect 20466 22094 20692 22146
rect 20412 22092 20692 22094
rect 20412 22082 20468 22092
rect 20300 21308 20468 21364
rect 20300 20914 20356 20926
rect 20300 20862 20302 20914
rect 20354 20862 20356 20914
rect 20300 19684 20356 20862
rect 20412 20804 20468 21308
rect 20412 20710 20468 20748
rect 20636 19908 20692 22092
rect 20636 19842 20692 19852
rect 20300 19618 20356 19628
rect 20524 19796 20580 19806
rect 20524 19460 20580 19740
rect 20524 19404 20692 19460
rect 20300 19236 20356 19246
rect 20188 19234 20356 19236
rect 20188 19182 20302 19234
rect 20354 19182 20356 19234
rect 20188 19180 20356 19182
rect 20300 19170 20356 19180
rect 20524 19236 20580 19246
rect 20524 19142 20580 19180
rect 20076 19070 20078 19122
rect 20130 19070 20132 19122
rect 20076 19058 20132 19070
rect 20636 19122 20692 19404
rect 20636 19070 20638 19122
rect 20690 19070 20692 19122
rect 19740 18946 19796 18956
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 20636 18676 20692 19070
rect 20636 18610 20692 18620
rect 20748 18116 20804 23100
rect 21308 22932 21364 22942
rect 21308 22838 21364 22876
rect 21532 21476 21588 26796
rect 21644 26786 21700 26796
rect 21980 26740 22036 26750
rect 21644 25508 21700 25518
rect 21644 25414 21700 25452
rect 21980 25506 22036 26684
rect 22652 26740 22708 26910
rect 23660 26964 23716 26974
rect 23660 26870 23716 26908
rect 22652 26674 22708 26684
rect 23324 26180 23380 26190
rect 21980 25454 21982 25506
rect 22034 25454 22036 25506
rect 21980 25284 22036 25454
rect 22204 25508 22260 25518
rect 23100 25508 23156 25518
rect 22204 25506 23156 25508
rect 22204 25454 22206 25506
rect 22258 25454 23102 25506
rect 23154 25454 23156 25506
rect 22204 25452 23156 25454
rect 22204 25442 22260 25452
rect 23100 25442 23156 25452
rect 23324 25394 23380 26124
rect 24556 26180 24612 37998
rect 26236 37492 26292 37502
rect 26236 37398 26292 37436
rect 25340 37266 25396 37278
rect 25340 37214 25342 37266
rect 25394 37214 25396 37266
rect 24780 36708 24836 36718
rect 24780 36614 24836 36652
rect 25340 26964 25396 37214
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 25340 26898 25396 26908
rect 25452 27746 25508 27758
rect 25452 27694 25454 27746
rect 25506 27694 25508 27746
rect 25452 26852 25508 27694
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 40012 27186 40068 27198
rect 40012 27134 40014 27186
rect 40066 27134 40068 27186
rect 25452 26292 25508 26796
rect 37884 27074 37940 27086
rect 37884 27022 37886 27074
rect 37938 27022 37940 27074
rect 25564 26292 25620 26302
rect 25452 26290 25620 26292
rect 25452 26238 25566 26290
rect 25618 26238 25620 26290
rect 25452 26236 25620 26238
rect 24556 26114 24612 26124
rect 25004 25506 25060 25518
rect 25004 25454 25006 25506
rect 25058 25454 25060 25506
rect 23324 25342 23326 25394
rect 23378 25342 23380 25394
rect 23324 25330 23380 25342
rect 23436 25394 23492 25406
rect 23436 25342 23438 25394
rect 23490 25342 23492 25394
rect 22540 25284 22596 25294
rect 22876 25284 22932 25294
rect 21980 25282 22596 25284
rect 21980 25230 22542 25282
rect 22594 25230 22596 25282
rect 21980 25228 22596 25230
rect 22540 25218 22596 25228
rect 22764 25282 22932 25284
rect 22764 25230 22878 25282
rect 22930 25230 22932 25282
rect 22764 25228 22932 25230
rect 22540 24724 22596 24734
rect 22764 24724 22820 25228
rect 22876 25218 22932 25228
rect 22876 24948 22932 24958
rect 22876 24854 22932 24892
rect 23436 24948 23492 25342
rect 25004 25284 25060 25454
rect 25004 25218 25060 25228
rect 25564 25284 25620 26236
rect 32060 26292 32116 26302
rect 26348 26178 26404 26190
rect 26348 26126 26350 26178
rect 26402 26126 26404 26178
rect 25676 25508 25732 25518
rect 25676 25506 26180 25508
rect 25676 25454 25678 25506
rect 25730 25454 26180 25506
rect 25676 25452 26180 25454
rect 25676 25442 25732 25452
rect 25564 25218 25620 25228
rect 26012 25284 26068 25294
rect 23436 24882 23492 24892
rect 25452 24836 25508 24846
rect 25452 24742 25508 24780
rect 22540 24722 22820 24724
rect 22540 24670 22542 24722
rect 22594 24670 22820 24722
rect 22540 24668 22820 24670
rect 25676 24722 25732 24734
rect 25676 24670 25678 24722
rect 25730 24670 25732 24722
rect 21980 23266 22036 23278
rect 21980 23214 21982 23266
rect 22034 23214 22036 23266
rect 21756 22932 21812 22942
rect 21756 22370 21812 22876
rect 21980 22820 22036 23214
rect 22092 23044 22148 23054
rect 22540 23044 22596 24668
rect 25676 24500 25732 24670
rect 25900 24724 25956 24734
rect 25788 24612 25844 24622
rect 25788 24518 25844 24556
rect 23100 23268 23156 23278
rect 23100 23266 23268 23268
rect 23100 23214 23102 23266
rect 23154 23214 23268 23266
rect 23100 23212 23268 23214
rect 23100 23202 23156 23212
rect 22988 23156 23044 23166
rect 22092 23042 22596 23044
rect 22092 22990 22094 23042
rect 22146 22990 22596 23042
rect 22092 22988 22596 22990
rect 22652 23154 23044 23156
rect 22652 23102 22990 23154
rect 23042 23102 23044 23154
rect 22652 23100 23044 23102
rect 22092 22978 22148 22988
rect 21980 22764 22260 22820
rect 21756 22318 21758 22370
rect 21810 22318 21812 22370
rect 21756 22306 21812 22318
rect 21980 22146 22036 22158
rect 21980 22094 21982 22146
rect 22034 22094 22036 22146
rect 21980 21700 22036 22094
rect 21980 21634 22036 21644
rect 20860 21420 21588 21476
rect 20860 19234 20916 21420
rect 20860 19182 20862 19234
rect 20914 19182 20916 19234
rect 20860 18452 20916 19182
rect 21196 20916 21252 20926
rect 21196 19234 21252 20860
rect 22092 20916 22148 20926
rect 21980 20802 22036 20814
rect 21980 20750 21982 20802
rect 22034 20750 22036 20802
rect 21308 20690 21364 20702
rect 21308 20638 21310 20690
rect 21362 20638 21364 20690
rect 21308 19684 21364 20638
rect 21644 20692 21700 20702
rect 21980 20692 22036 20750
rect 22092 20802 22148 20860
rect 22092 20750 22094 20802
rect 22146 20750 22148 20802
rect 22092 20738 22148 20750
rect 21644 20690 21980 20692
rect 21644 20638 21646 20690
rect 21698 20638 21980 20690
rect 21644 20636 21980 20638
rect 21644 20626 21700 20636
rect 21980 20626 22036 20636
rect 21420 20578 21476 20590
rect 21420 20526 21422 20578
rect 21474 20526 21476 20578
rect 21420 20468 21476 20526
rect 22204 20580 22260 22764
rect 22652 22036 22708 23100
rect 22988 23090 23044 23100
rect 22764 22484 22820 22494
rect 22764 22370 22820 22428
rect 22764 22318 22766 22370
rect 22818 22318 22820 22370
rect 22764 22306 22820 22318
rect 22428 21980 22708 22036
rect 22316 21812 22372 21822
rect 22316 20802 22372 21756
rect 22428 20914 22484 21980
rect 23212 21924 23268 23212
rect 23324 23154 23380 23166
rect 23324 23102 23326 23154
rect 23378 23102 23380 23154
rect 23324 22484 23380 23102
rect 25676 22708 25732 24444
rect 25340 22652 25732 22708
rect 23436 22484 23492 22494
rect 23324 22482 23492 22484
rect 23324 22430 23438 22482
rect 23490 22430 23492 22482
rect 23324 22428 23492 22430
rect 23436 22418 23492 22428
rect 23100 21812 23156 21822
rect 22428 20862 22430 20914
rect 22482 20862 22484 20914
rect 22428 20850 22484 20862
rect 22540 21810 23156 21812
rect 22540 21758 23102 21810
rect 23154 21758 23156 21810
rect 22540 21756 23156 21758
rect 22316 20750 22318 20802
rect 22370 20750 22372 20802
rect 22316 20738 22372 20750
rect 22540 20802 22596 21756
rect 23100 21746 23156 21756
rect 22540 20750 22542 20802
rect 22594 20750 22596 20802
rect 22540 20738 22596 20750
rect 22652 21586 22708 21598
rect 22652 21534 22654 21586
rect 22706 21534 22708 21586
rect 22652 20804 22708 21534
rect 22876 21588 22932 21598
rect 22876 21494 22932 21532
rect 22652 20738 22708 20748
rect 22204 20514 22260 20524
rect 22876 20690 22932 20702
rect 22876 20638 22878 20690
rect 22930 20638 22932 20690
rect 21420 20132 21476 20412
rect 22876 20468 22932 20638
rect 22988 20580 23044 20590
rect 22988 20486 23044 20524
rect 22876 20402 22932 20412
rect 21476 20076 21812 20132
rect 21420 20066 21476 20076
rect 21364 19628 21588 19684
rect 21308 19618 21364 19628
rect 21196 19182 21198 19234
rect 21250 19182 21252 19234
rect 21196 19170 21252 19182
rect 21532 19234 21588 19628
rect 21532 19182 21534 19234
rect 21586 19182 21588 19234
rect 21532 19170 21588 19182
rect 21756 19124 21812 20076
rect 22428 19234 22484 19246
rect 22428 19182 22430 19234
rect 22482 19182 22484 19234
rect 21644 19122 21812 19124
rect 21644 19070 21758 19122
rect 21810 19070 21812 19122
rect 21644 19068 21812 19070
rect 21644 19012 21700 19068
rect 21756 19058 21812 19068
rect 22316 19122 22372 19134
rect 22316 19070 22318 19122
rect 22370 19070 22372 19122
rect 20860 18386 20916 18396
rect 21420 18956 21700 19012
rect 21868 19012 21924 19022
rect 20748 18050 20804 18060
rect 21420 18004 21476 18956
rect 21868 18918 21924 18956
rect 21532 18676 21588 18686
rect 21532 18450 21588 18620
rect 21868 18676 21924 18686
rect 21532 18398 21534 18450
rect 21586 18398 21588 18450
rect 21532 18386 21588 18398
rect 21756 18562 21812 18574
rect 21756 18510 21758 18562
rect 21810 18510 21812 18562
rect 21756 18228 21812 18510
rect 21756 18162 21812 18172
rect 21868 18004 21924 18620
rect 22316 18564 22372 19070
rect 22428 18676 22484 19182
rect 22876 19234 22932 19246
rect 22876 19182 22878 19234
rect 22930 19182 22932 19234
rect 22428 18610 22484 18620
rect 22764 19012 22820 19022
rect 22764 18674 22820 18956
rect 22764 18622 22766 18674
rect 22818 18622 22820 18674
rect 22764 18610 22820 18622
rect 22316 18498 22372 18508
rect 22876 18564 22932 19182
rect 22876 18498 22932 18508
rect 22988 18562 23044 18574
rect 22988 18510 22990 18562
rect 23042 18510 23044 18562
rect 22540 18452 22596 18462
rect 22540 18358 22596 18396
rect 22988 18452 23044 18510
rect 22988 18386 23044 18396
rect 23212 18450 23268 21868
rect 25340 21812 25396 22652
rect 25564 22484 25620 22494
rect 25116 21756 25396 21812
rect 25452 22482 25620 22484
rect 25452 22430 25566 22482
rect 25618 22430 25620 22482
rect 25452 22428 25620 22430
rect 25452 21812 25508 22428
rect 25564 22418 25620 22428
rect 23548 21700 23604 21710
rect 23324 21586 23380 21598
rect 23324 21534 23326 21586
rect 23378 21534 23380 21586
rect 23324 21476 23380 21534
rect 23324 21410 23380 21420
rect 23548 21586 23604 21644
rect 24220 21698 24276 21710
rect 24220 21646 24222 21698
rect 24274 21646 24276 21698
rect 23548 21534 23550 21586
rect 23602 21534 23604 21586
rect 23324 20804 23380 20814
rect 23324 20130 23380 20748
rect 23324 20078 23326 20130
rect 23378 20078 23380 20130
rect 23324 20066 23380 20078
rect 23436 20692 23492 20702
rect 23436 19458 23492 20636
rect 23436 19406 23438 19458
rect 23490 19406 23492 19458
rect 23436 19394 23492 19406
rect 23548 19236 23604 21534
rect 23884 21586 23940 21598
rect 23884 21534 23886 21586
rect 23938 21534 23940 21586
rect 23884 20580 23940 21534
rect 24220 21476 24276 21646
rect 24276 21420 24612 21476
rect 24220 21410 24276 21420
rect 23884 20514 23940 20524
rect 23436 19180 23604 19236
rect 23660 19908 23716 19918
rect 23660 19236 23716 19852
rect 23772 19460 23828 19470
rect 23772 19366 23828 19404
rect 24108 19236 24164 19246
rect 23660 19234 24164 19236
rect 23660 19182 24110 19234
rect 24162 19182 24164 19234
rect 23660 19180 24164 19182
rect 23436 18676 23492 19180
rect 23660 19122 23716 19180
rect 24108 19170 24164 19180
rect 24444 19124 24500 19134
rect 23660 19070 23662 19122
rect 23714 19070 23716 19122
rect 23660 19058 23716 19070
rect 24332 19068 24444 19124
rect 23436 18610 23492 18620
rect 23884 18676 23940 18686
rect 23884 18562 23940 18620
rect 24220 18676 24276 18686
rect 24220 18582 24276 18620
rect 23884 18510 23886 18562
rect 23938 18510 23940 18562
rect 23884 18498 23940 18510
rect 23996 18564 24052 18574
rect 23212 18398 23214 18450
rect 23266 18398 23268 18450
rect 21980 18340 22036 18350
rect 21980 18246 22036 18284
rect 23212 18340 23268 18398
rect 23212 18274 23268 18284
rect 23660 18452 23716 18462
rect 22652 18228 22708 18238
rect 21420 17948 21700 18004
rect 20412 17892 20468 17902
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 19628 16716 19908 16772
rect 18172 16658 18452 16660
rect 18172 16606 18174 16658
rect 18226 16606 18452 16658
rect 18172 16604 18452 16606
rect 18172 16594 18228 16604
rect 18284 16100 18340 16110
rect 18060 16098 18340 16100
rect 18060 16046 18286 16098
rect 18338 16046 18340 16098
rect 18060 16044 18340 16046
rect 18284 16034 18340 16044
rect 18396 16100 18452 16604
rect 18396 16034 18452 16044
rect 18956 16100 19012 16110
rect 18956 16006 19012 16044
rect 19852 16100 19908 16716
rect 20412 16322 20468 17836
rect 21420 17666 21476 17678
rect 21420 17614 21422 17666
rect 21474 17614 21476 17666
rect 21420 16882 21476 17614
rect 21644 17554 21700 17948
rect 21644 17502 21646 17554
rect 21698 17502 21700 17554
rect 21644 17490 21700 17502
rect 21756 17948 21924 18004
rect 22428 18226 22708 18228
rect 22428 18174 22654 18226
rect 22706 18174 22708 18226
rect 22428 18172 22708 18174
rect 21756 17332 21812 17948
rect 22428 17890 22484 18172
rect 22652 18162 22708 18172
rect 23548 18228 23604 18238
rect 22428 17838 22430 17890
rect 22482 17838 22484 17890
rect 22428 17826 22484 17838
rect 22204 17780 22260 17790
rect 22204 17686 22260 17724
rect 23548 17666 23604 18172
rect 23660 17778 23716 18396
rect 23996 18004 24052 18508
rect 23660 17726 23662 17778
rect 23714 17726 23716 17778
rect 23660 17714 23716 17726
rect 23772 17948 24052 18004
rect 23548 17614 23550 17666
rect 23602 17614 23604 17666
rect 23548 17602 23604 17614
rect 21420 16830 21422 16882
rect 21474 16830 21476 16882
rect 21420 16548 21476 16830
rect 20412 16270 20414 16322
rect 20466 16270 20468 16322
rect 20412 16258 20468 16270
rect 20524 16492 21476 16548
rect 21644 17276 21812 17332
rect 22764 17442 22820 17454
rect 22764 17390 22766 17442
rect 22818 17390 22820 17442
rect 19852 16006 19908 16044
rect 20076 16100 20132 16110
rect 20076 16006 20132 16044
rect 18508 15988 18564 15998
rect 18508 15894 18564 15932
rect 18620 15874 18676 15886
rect 18620 15822 18622 15874
rect 18674 15822 18676 15874
rect 18620 15540 18676 15822
rect 17500 14530 17556 14588
rect 18172 15484 18676 15540
rect 19068 15876 19124 15886
rect 18172 14642 18228 15484
rect 19068 15426 19124 15820
rect 19964 15876 20020 15914
rect 19964 15810 20020 15820
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 19068 15374 19070 15426
rect 19122 15374 19124 15426
rect 19068 15362 19124 15374
rect 18172 14590 18174 14642
rect 18226 14590 18228 14642
rect 18172 14578 18228 14590
rect 18396 15314 18452 15326
rect 18396 15262 18398 15314
rect 18450 15262 18452 15314
rect 18396 14644 18452 15262
rect 18396 14578 18452 14588
rect 20300 14644 20356 14654
rect 20524 14644 20580 16492
rect 21308 16324 21364 16334
rect 20636 16322 21364 16324
rect 20636 16270 21310 16322
rect 21362 16270 21364 16322
rect 20636 16268 21364 16270
rect 20636 16098 20692 16268
rect 21308 16258 21364 16268
rect 21644 16322 21700 17276
rect 21756 17108 21812 17118
rect 21756 17014 21812 17052
rect 21644 16270 21646 16322
rect 21698 16270 21700 16322
rect 21644 16258 21700 16270
rect 21308 16100 21364 16110
rect 20636 16046 20638 16098
rect 20690 16046 20692 16098
rect 20636 16034 20692 16046
rect 21196 16098 21364 16100
rect 21196 16046 21310 16098
rect 21362 16046 21364 16098
rect 21196 16044 21364 16046
rect 21196 15202 21252 16044
rect 21308 16034 21364 16044
rect 22764 16098 22820 17390
rect 23772 17442 23828 17948
rect 24332 17892 24388 19068
rect 24444 19030 24500 19068
rect 24108 17836 24388 17892
rect 23996 17668 24052 17678
rect 24108 17668 24164 17836
rect 23996 17666 24164 17668
rect 23996 17614 23998 17666
rect 24050 17614 24164 17666
rect 23996 17612 24164 17614
rect 24332 17668 24388 17678
rect 24332 17666 24500 17668
rect 24332 17614 24334 17666
rect 24386 17614 24500 17666
rect 24332 17612 24500 17614
rect 23996 17602 24052 17612
rect 24332 17602 24388 17612
rect 23772 17390 23774 17442
rect 23826 17390 23828 17442
rect 23772 17108 23828 17390
rect 23772 17042 23828 17052
rect 22764 16046 22766 16098
rect 22818 16046 22820 16098
rect 22764 16034 22820 16046
rect 23884 16772 23940 16782
rect 23884 16100 23940 16716
rect 22428 15876 22484 15886
rect 22316 15874 22484 15876
rect 22316 15822 22430 15874
rect 22482 15822 22484 15874
rect 22316 15820 22484 15822
rect 22316 15426 22372 15820
rect 22428 15810 22484 15820
rect 22316 15374 22318 15426
rect 22370 15374 22372 15426
rect 22316 15362 22372 15374
rect 21644 15316 21700 15326
rect 21644 15222 21700 15260
rect 22988 15316 23044 15326
rect 21196 15150 21198 15202
rect 21250 15150 21252 15202
rect 20300 14642 20580 14644
rect 20300 14590 20302 14642
rect 20354 14590 20580 14642
rect 20300 14588 20580 14590
rect 20860 14644 20916 14654
rect 20300 14578 20356 14588
rect 20860 14550 20916 14588
rect 17500 14478 17502 14530
rect 17554 14478 17556 14530
rect 17500 14466 17556 14478
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 21196 8428 21252 15150
rect 21420 14644 21476 14654
rect 21420 14550 21476 14588
rect 22988 12962 23044 15260
rect 23884 14530 23940 16044
rect 23884 14478 23886 14530
rect 23938 14478 23940 14530
rect 23884 14466 23940 14478
rect 24220 15428 24276 15438
rect 24220 14530 24276 15372
rect 24220 14478 24222 14530
rect 24274 14478 24276 14530
rect 24220 14466 24276 14478
rect 24444 15202 24500 17612
rect 24556 16772 24612 21420
rect 24780 19012 24836 19022
rect 24780 18918 24836 18956
rect 25116 19010 25172 21756
rect 25452 21746 25508 21756
rect 25564 22260 25620 22270
rect 25564 21810 25620 22204
rect 25564 21758 25566 21810
rect 25618 21758 25620 21810
rect 25564 21746 25620 21758
rect 25788 21700 25844 21710
rect 25676 21644 25788 21700
rect 25452 21588 25508 21598
rect 25452 21494 25508 21532
rect 25564 21364 25620 21374
rect 25564 21270 25620 21308
rect 25452 20690 25508 20702
rect 25452 20638 25454 20690
rect 25506 20638 25508 20690
rect 25340 20580 25396 20590
rect 25340 20242 25396 20524
rect 25340 20190 25342 20242
rect 25394 20190 25396 20242
rect 25340 20178 25396 20190
rect 25452 20244 25508 20638
rect 25228 20018 25284 20030
rect 25228 19966 25230 20018
rect 25282 19966 25284 20018
rect 25228 19908 25284 19966
rect 25228 19842 25284 19852
rect 25340 19012 25396 19022
rect 25116 18958 25118 19010
rect 25170 18958 25172 19010
rect 24892 17442 24948 17454
rect 24892 17390 24894 17442
rect 24946 17390 24948 17442
rect 24892 17108 24948 17390
rect 24892 17042 24948 17052
rect 24556 16706 24612 16716
rect 25116 15428 25172 18958
rect 25228 19010 25396 19012
rect 25228 18958 25342 19010
rect 25394 18958 25396 19010
rect 25228 18956 25396 18958
rect 25228 18452 25284 18956
rect 25340 18946 25396 18956
rect 25452 18788 25508 20188
rect 25564 20244 25620 20254
rect 25676 20244 25732 21644
rect 25788 21634 25844 21644
rect 25564 20242 25732 20244
rect 25564 20190 25566 20242
rect 25618 20190 25732 20242
rect 25564 20188 25732 20190
rect 25564 20178 25620 20188
rect 25676 19234 25732 20188
rect 25788 21476 25844 21486
rect 25788 20242 25844 21420
rect 25788 20190 25790 20242
rect 25842 20190 25844 20242
rect 25788 20178 25844 20190
rect 25900 20242 25956 24668
rect 26012 22484 26068 25228
rect 26124 24052 26180 25452
rect 26348 24836 26404 26126
rect 28476 26178 28532 26190
rect 28476 26126 28478 26178
rect 28530 26126 28532 26178
rect 28252 25732 28308 25742
rect 27916 25730 28308 25732
rect 27916 25678 28254 25730
rect 28306 25678 28308 25730
rect 27916 25676 28308 25678
rect 27804 25618 27860 25630
rect 27804 25566 27806 25618
rect 27858 25566 27860 25618
rect 27020 25508 27076 25518
rect 26908 25452 27020 25508
rect 26908 25172 26964 25452
rect 27020 25442 27076 25452
rect 27804 25508 27860 25566
rect 27804 25442 27860 25452
rect 26684 25116 26964 25172
rect 26684 24946 26740 25116
rect 27916 25060 27972 25676
rect 28252 25666 28308 25676
rect 28476 25508 28532 26126
rect 28252 25452 28532 25508
rect 28924 26178 28980 26190
rect 28924 26126 28926 26178
rect 28978 26126 28980 26178
rect 27468 25004 27972 25060
rect 28140 25394 28196 25406
rect 28140 25342 28142 25394
rect 28194 25342 28196 25394
rect 26684 24894 26686 24946
rect 26738 24894 26740 24946
rect 26684 24882 26740 24894
rect 26908 24948 26964 24958
rect 26348 24770 26404 24780
rect 26236 24724 26292 24734
rect 26236 24630 26292 24668
rect 26460 24722 26516 24734
rect 26460 24670 26462 24722
rect 26514 24670 26516 24722
rect 26236 24500 26292 24510
rect 26460 24500 26516 24670
rect 26908 24724 26964 24892
rect 27468 24946 27524 25004
rect 27468 24894 27470 24946
rect 27522 24894 27524 24946
rect 27468 24882 27524 24894
rect 27580 24836 27636 24846
rect 27580 24742 27636 24780
rect 26908 24630 26964 24668
rect 27244 24722 27300 24734
rect 27244 24670 27246 24722
rect 27298 24670 27300 24722
rect 26292 24444 26516 24500
rect 26796 24610 26852 24622
rect 26796 24558 26798 24610
rect 26850 24558 26852 24610
rect 26236 24434 26292 24444
rect 26460 24052 26516 24062
rect 26124 24050 26516 24052
rect 26124 23998 26462 24050
rect 26514 23998 26516 24050
rect 26124 23996 26516 23998
rect 26460 23986 26516 23996
rect 26572 23938 26628 23950
rect 26572 23886 26574 23938
rect 26626 23886 26628 23938
rect 26348 23828 26404 23838
rect 26236 23772 26348 23828
rect 26012 22390 26068 22428
rect 26124 23154 26180 23166
rect 26124 23102 26126 23154
rect 26178 23102 26180 23154
rect 26124 22372 26180 23102
rect 26124 22306 26180 22316
rect 26236 21810 26292 23772
rect 26348 23734 26404 23772
rect 26460 23268 26516 23278
rect 26572 23268 26628 23886
rect 26796 23938 26852 24558
rect 27244 24612 27300 24670
rect 27244 24546 27300 24556
rect 27692 24722 27748 24734
rect 27692 24670 27694 24722
rect 27746 24670 27748 24722
rect 27692 24612 27748 24670
rect 26796 23886 26798 23938
rect 26850 23886 26852 23938
rect 26796 23874 26852 23886
rect 26460 23266 26628 23268
rect 26460 23214 26462 23266
rect 26514 23214 26628 23266
rect 26460 23212 26628 23214
rect 26460 22372 26516 23212
rect 26460 22306 26516 22316
rect 26796 22484 26852 22494
rect 26236 21758 26238 21810
rect 26290 21758 26292 21810
rect 26236 21746 26292 21758
rect 26124 21698 26180 21710
rect 26124 21646 26126 21698
rect 26178 21646 26180 21698
rect 26124 21476 26180 21646
rect 26348 21700 26404 21710
rect 26348 21606 26404 21644
rect 26124 21410 26180 21420
rect 25900 20190 25902 20242
rect 25954 20190 25956 20242
rect 25900 20178 25956 20190
rect 26460 21364 26516 21374
rect 26012 20020 26068 20030
rect 25676 19182 25678 19234
rect 25730 19182 25732 19234
rect 25676 19170 25732 19182
rect 25900 20018 26068 20020
rect 25900 19966 26014 20018
rect 26066 19966 26068 20018
rect 25900 19964 26068 19966
rect 25228 17892 25284 18396
rect 25228 17826 25284 17836
rect 25340 18732 25508 18788
rect 25564 19012 25620 19022
rect 25228 17444 25284 17454
rect 25228 17350 25284 17388
rect 25116 15362 25172 15372
rect 25228 15876 25284 15886
rect 24444 15150 24446 15202
rect 24498 15150 24500 15202
rect 24220 14306 24276 14318
rect 24220 14254 24222 14306
rect 24274 14254 24276 14306
rect 24220 13636 24276 14254
rect 23772 13580 24276 13636
rect 23772 13074 23828 13580
rect 23772 13022 23774 13074
rect 23826 13022 23828 13074
rect 23772 13010 23828 13022
rect 22988 12910 22990 12962
rect 23042 12910 23044 12962
rect 22988 12898 23044 12910
rect 24444 8428 24500 15150
rect 25228 15204 25284 15820
rect 25340 15316 25396 18732
rect 25564 18676 25620 18956
rect 25564 18610 25620 18620
rect 25788 18450 25844 18462
rect 25788 18398 25790 18450
rect 25842 18398 25844 18450
rect 25452 18340 25508 18350
rect 25788 18340 25844 18398
rect 25452 18338 25844 18340
rect 25452 18286 25454 18338
rect 25506 18286 25844 18338
rect 25452 18284 25844 18286
rect 25452 18116 25508 18284
rect 25452 18050 25508 18060
rect 25788 17442 25844 17454
rect 25788 17390 25790 17442
rect 25842 17390 25844 17442
rect 25788 15876 25844 17390
rect 25900 17444 25956 19964
rect 26012 19954 26068 19964
rect 26348 20018 26404 20030
rect 26348 19966 26350 20018
rect 26402 19966 26404 20018
rect 26348 19124 26404 19966
rect 26236 18564 26292 18574
rect 26236 18470 26292 18508
rect 26012 18452 26068 18462
rect 26012 18358 26068 18396
rect 26124 17668 26180 17678
rect 26348 17668 26404 19068
rect 26460 18450 26516 21308
rect 26796 20244 26852 22428
rect 27692 22372 27748 24556
rect 27804 24722 27860 24734
rect 27804 24670 27806 24722
rect 27858 24670 27860 24722
rect 27804 24500 27860 24670
rect 27804 23940 27860 24444
rect 27804 23874 27860 23884
rect 28140 24724 28196 25342
rect 28252 25396 28308 25452
rect 28252 25302 28308 25340
rect 28364 25284 28420 25294
rect 28364 24946 28420 25228
rect 28364 24894 28366 24946
rect 28418 24894 28420 24946
rect 28364 24882 28420 24894
rect 28924 24948 28980 26126
rect 29484 26180 29540 26190
rect 29932 26180 29988 26190
rect 29484 26178 29988 26180
rect 29484 26126 29486 26178
rect 29538 26126 29934 26178
rect 29986 26126 29988 26178
rect 29484 26124 29988 26126
rect 29036 26068 29092 26078
rect 29260 26068 29316 26078
rect 29036 26066 29316 26068
rect 29036 26014 29038 26066
rect 29090 26014 29262 26066
rect 29314 26014 29316 26066
rect 29036 26012 29316 26014
rect 29036 26002 29092 26012
rect 29260 26002 29316 26012
rect 29148 25508 29204 25518
rect 29484 25508 29540 26124
rect 29932 26114 29988 26124
rect 30044 26066 30100 26078
rect 30044 26014 30046 26066
rect 30098 26014 30100 26066
rect 29148 25506 29540 25508
rect 29148 25454 29150 25506
rect 29202 25454 29540 25506
rect 29148 25452 29540 25454
rect 29596 25620 29652 25630
rect 29148 25284 29204 25452
rect 29148 25218 29204 25228
rect 29596 25060 29652 25564
rect 29932 25620 29988 25630
rect 30044 25620 30100 26014
rect 29932 25618 30100 25620
rect 29932 25566 29934 25618
rect 29986 25566 30100 25618
rect 29932 25564 30100 25566
rect 32060 25620 32116 26236
rect 37660 26292 37716 26302
rect 37660 26198 37716 26236
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 29932 25554 29988 25564
rect 32060 25526 32116 25564
rect 37660 25508 37716 25518
rect 37660 25414 37716 25452
rect 37884 25284 37940 27022
rect 40012 26292 40068 27134
rect 40012 26226 40068 26236
rect 39900 26178 39956 26190
rect 39900 26126 39902 26178
rect 39954 26126 39956 26178
rect 39900 25620 39956 26126
rect 39900 25554 39956 25564
rect 40012 25618 40068 25630
rect 40012 25566 40014 25618
rect 40066 25566 40068 25618
rect 37884 25218 37940 25228
rect 29148 25004 29652 25060
rect 29036 24948 29092 24958
rect 28924 24946 29092 24948
rect 28924 24894 29038 24946
rect 29090 24894 29092 24946
rect 28924 24892 29092 24894
rect 29036 24882 29092 24892
rect 29148 24946 29204 25004
rect 29148 24894 29150 24946
rect 29202 24894 29204 24946
rect 29148 24882 29204 24894
rect 40012 24948 40068 25566
rect 40012 24882 40068 24892
rect 28140 23938 28196 24668
rect 28140 23886 28142 23938
rect 28194 23886 28196 23938
rect 28140 23874 28196 23886
rect 28476 24724 28532 24734
rect 28476 23826 28532 24668
rect 28700 24722 28756 24734
rect 28700 24670 28702 24722
rect 28754 24670 28756 24722
rect 28700 24612 28756 24670
rect 28700 24546 28756 24556
rect 28924 24722 28980 24734
rect 28924 24670 28926 24722
rect 28978 24670 28980 24722
rect 28924 24500 28980 24670
rect 29260 24724 29316 24734
rect 29260 24630 29316 24668
rect 29820 24724 29876 24734
rect 28924 24434 28980 24444
rect 28476 23774 28478 23826
rect 28530 23774 28532 23826
rect 28476 23762 28532 23774
rect 29036 22540 29764 22596
rect 27692 22306 27748 22316
rect 28252 22372 28308 22382
rect 28252 22278 28308 22316
rect 28700 22372 28756 22382
rect 29036 22372 29092 22540
rect 28700 22370 29092 22372
rect 28700 22318 28702 22370
rect 28754 22318 29092 22370
rect 28700 22316 29092 22318
rect 29148 22370 29204 22382
rect 29148 22318 29150 22370
rect 29202 22318 29204 22370
rect 28700 22306 28756 22316
rect 28140 22260 28196 22270
rect 28140 22166 28196 22204
rect 28028 22146 28084 22158
rect 28028 22094 28030 22146
rect 28082 22094 28084 22146
rect 28028 21924 28084 22094
rect 27132 21700 27188 21710
rect 27132 21606 27188 21644
rect 26908 21588 26964 21598
rect 26908 21494 26964 21532
rect 27580 21586 27636 21598
rect 27580 21534 27582 21586
rect 27634 21534 27636 21586
rect 26796 20020 26852 20188
rect 27020 21474 27076 21486
rect 27020 21422 27022 21474
rect 27074 21422 27076 21474
rect 27020 20188 27076 21422
rect 27580 21028 27636 21534
rect 27580 20962 27636 20972
rect 27020 20132 27636 20188
rect 27580 20130 27636 20132
rect 27580 20078 27582 20130
rect 27634 20078 27636 20130
rect 27580 20066 27636 20078
rect 26908 20020 26964 20030
rect 26796 19964 26908 20020
rect 26964 19964 27076 20020
rect 26908 19926 26964 19964
rect 26460 18398 26462 18450
rect 26514 18398 26516 18450
rect 26460 18386 26516 18398
rect 26908 19236 26964 19246
rect 26124 17666 26348 17668
rect 26124 17614 26126 17666
rect 26178 17614 26348 17666
rect 26124 17612 26348 17614
rect 26124 17602 26180 17612
rect 26348 17574 26404 17612
rect 26460 17780 26516 17790
rect 26460 17666 26516 17724
rect 26460 17614 26462 17666
rect 26514 17614 26516 17666
rect 26460 17602 26516 17614
rect 26796 17554 26852 17566
rect 26796 17502 26798 17554
rect 26850 17502 26852 17554
rect 26012 17444 26068 17454
rect 26684 17444 26740 17454
rect 25900 17388 26012 17444
rect 26012 17378 26068 17388
rect 26572 17442 26740 17444
rect 26572 17390 26686 17442
rect 26738 17390 26740 17442
rect 26572 17388 26740 17390
rect 26572 15988 26628 17388
rect 26684 17378 26740 17388
rect 26796 17332 26852 17502
rect 26908 17554 26964 19180
rect 26908 17502 26910 17554
rect 26962 17502 26964 17554
rect 26908 17490 26964 17502
rect 26908 17332 26964 17342
rect 26796 17276 26908 17332
rect 26908 17266 26964 17276
rect 26684 17108 26740 17118
rect 27020 17108 27076 19964
rect 28028 19236 28084 21868
rect 28812 21476 28868 21486
rect 29148 21476 29204 22318
rect 29708 21810 29764 22540
rect 29708 21758 29710 21810
rect 29762 21758 29764 21810
rect 29708 21746 29764 21758
rect 29820 21588 29876 24668
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 30156 22484 30212 22494
rect 30044 22428 30156 22484
rect 29932 22260 29988 22270
rect 29932 22166 29988 22204
rect 29932 21812 29988 21822
rect 30044 21812 30100 22428
rect 30156 22418 30212 22428
rect 32060 22484 32116 22494
rect 32060 22390 32116 22428
rect 37660 22484 37716 22494
rect 37660 22370 37716 22428
rect 37660 22318 37662 22370
rect 37714 22318 37716 22370
rect 37660 22306 37716 22318
rect 40012 22482 40068 22494
rect 40012 22430 40014 22482
rect 40066 22430 40068 22482
rect 40012 22260 40068 22430
rect 40012 22194 40068 22204
rect 29932 21810 30100 21812
rect 29932 21758 29934 21810
rect 29986 21758 30100 21810
rect 29932 21756 30100 21758
rect 29932 21746 29988 21756
rect 30044 21588 30100 21598
rect 29820 21586 30100 21588
rect 29820 21534 30046 21586
rect 30098 21534 30100 21586
rect 29820 21532 30100 21534
rect 28812 21474 29204 21476
rect 28812 21422 28814 21474
rect 28866 21422 29204 21474
rect 28812 21420 29204 21422
rect 28812 20188 28868 21420
rect 29036 21028 29092 21038
rect 29036 20802 29092 20972
rect 29036 20750 29038 20802
rect 29090 20750 29092 20802
rect 29036 20738 29092 20750
rect 29372 20804 29428 20814
rect 30044 20804 30100 21532
rect 37660 21588 37716 21598
rect 37660 21494 37716 21532
rect 40012 21588 40068 21598
rect 40012 21474 40068 21532
rect 40012 21422 40014 21474
rect 40066 21422 40068 21474
rect 40012 21410 40068 21422
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 40012 20916 40068 20926
rect 40012 20822 40068 20860
rect 29372 20802 30100 20804
rect 29372 20750 29374 20802
rect 29426 20750 30100 20802
rect 29372 20748 30100 20750
rect 29372 20738 29428 20748
rect 29260 20580 29316 20590
rect 29260 20486 29316 20524
rect 29708 20580 29764 20590
rect 28812 20132 29316 20188
rect 28812 20020 28868 20132
rect 28028 19170 28084 19180
rect 28700 19796 28756 19806
rect 28700 19234 28756 19740
rect 28700 19182 28702 19234
rect 28754 19182 28756 19234
rect 28700 19170 28756 19182
rect 28140 19124 28196 19134
rect 28140 19030 28196 19068
rect 28028 19010 28084 19022
rect 28028 18958 28030 19010
rect 28082 18958 28084 19010
rect 28028 18788 28084 18958
rect 28252 19012 28308 19022
rect 28252 18918 28308 18956
rect 28028 18722 28084 18732
rect 28812 18674 28868 19964
rect 29260 19908 29316 20132
rect 29260 19234 29316 19852
rect 29708 19906 29764 20524
rect 30044 20130 30100 20748
rect 37660 20804 37716 20814
rect 37660 20710 37716 20748
rect 30044 20078 30046 20130
rect 30098 20078 30100 20130
rect 30044 20066 30100 20078
rect 30156 20132 30212 20142
rect 30156 20038 30212 20076
rect 32060 20020 32116 20030
rect 29708 19854 29710 19906
rect 29762 19854 29764 19906
rect 29708 19842 29764 19854
rect 30716 19908 30772 19918
rect 30716 19814 30772 19852
rect 30156 19796 30212 19806
rect 30156 19702 30212 19740
rect 32060 19346 32116 19964
rect 37660 20020 37716 20030
rect 37660 19926 37716 19964
rect 40012 19794 40068 19806
rect 40012 19742 40014 19794
rect 40066 19742 40068 19794
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 40012 19572 40068 19742
rect 40012 19506 40068 19516
rect 32060 19294 32062 19346
rect 32114 19294 32116 19346
rect 32060 19282 32116 19294
rect 29260 19182 29262 19234
rect 29314 19182 29316 19234
rect 29260 19170 29316 19182
rect 29932 19124 29988 19134
rect 29932 19030 29988 19068
rect 28812 18622 28814 18674
rect 28866 18622 28868 18674
rect 28812 18610 28868 18622
rect 27356 18564 27412 18574
rect 27356 18470 27412 18508
rect 27468 18562 27524 18574
rect 27468 18510 27470 18562
rect 27522 18510 27524 18562
rect 27468 18004 27524 18510
rect 27692 18452 27748 18462
rect 27692 18450 28532 18452
rect 27692 18398 27694 18450
rect 27746 18398 28532 18450
rect 27692 18396 28532 18398
rect 27692 18386 27748 18396
rect 27132 17948 27524 18004
rect 27580 18228 27636 18238
rect 27132 17220 27188 17948
rect 27244 17780 27300 17790
rect 27244 17778 27412 17780
rect 27244 17726 27246 17778
rect 27298 17726 27412 17778
rect 27244 17724 27412 17726
rect 27244 17714 27300 17724
rect 27132 17164 27300 17220
rect 26684 17106 27076 17108
rect 26684 17054 26686 17106
rect 26738 17054 27076 17106
rect 26684 17052 27076 17054
rect 26684 17042 26740 17052
rect 27020 16884 27076 17052
rect 27020 16790 27076 16828
rect 27132 16996 27188 17006
rect 26908 16100 26964 16110
rect 27132 16100 27188 16940
rect 27244 16210 27300 17164
rect 27356 17108 27412 17724
rect 27356 17042 27412 17052
rect 27580 17666 27636 18172
rect 27580 17614 27582 17666
rect 27634 17614 27636 17666
rect 27580 16996 27636 17614
rect 28364 17668 28420 17678
rect 28364 17574 28420 17612
rect 27916 17556 27972 17566
rect 27916 17462 27972 17500
rect 27692 17442 27748 17454
rect 27692 17390 27694 17442
rect 27746 17390 27748 17442
rect 27692 17332 27748 17390
rect 27692 17266 27748 17276
rect 27804 17444 27860 17454
rect 27804 17220 27860 17388
rect 27804 17164 27972 17220
rect 27692 17108 27748 17118
rect 27692 16996 27748 17052
rect 27804 16996 27860 17006
rect 27692 16994 27860 16996
rect 27692 16942 27806 16994
rect 27858 16942 27860 16994
rect 27692 16940 27860 16942
rect 27580 16930 27636 16940
rect 27804 16930 27860 16940
rect 27244 16158 27246 16210
rect 27298 16158 27300 16210
rect 27244 16146 27300 16158
rect 26908 16098 27188 16100
rect 26908 16046 26910 16098
rect 26962 16046 27188 16098
rect 26908 16044 27188 16046
rect 27692 16100 27748 16110
rect 26908 16034 26964 16044
rect 27692 16006 27748 16044
rect 26572 15922 26628 15932
rect 27244 15988 27300 15998
rect 27244 15894 27300 15932
rect 25788 15810 25844 15820
rect 27132 15874 27188 15886
rect 27132 15822 27134 15874
rect 27186 15822 27188 15874
rect 27132 15764 27188 15822
rect 27916 15764 27972 17164
rect 27132 15708 27972 15764
rect 28140 16884 28196 16894
rect 28140 16210 28196 16828
rect 28140 16158 28142 16210
rect 28194 16158 28196 16210
rect 27020 15540 27076 15550
rect 26796 15538 27076 15540
rect 26796 15486 27022 15538
rect 27074 15486 27076 15538
rect 26796 15484 27076 15486
rect 26236 15428 26292 15438
rect 26236 15334 26292 15372
rect 26348 15316 26404 15326
rect 26684 15316 26740 15326
rect 25396 15260 25732 15316
rect 25340 15222 25396 15260
rect 24556 14532 24612 14542
rect 25004 14532 25060 14542
rect 24556 14530 25060 14532
rect 24556 14478 24558 14530
rect 24610 14478 25006 14530
rect 25058 14478 25060 14530
rect 24556 14476 25060 14478
rect 25228 14532 25284 15148
rect 25676 14644 25732 15260
rect 26348 15314 26740 15316
rect 26348 15262 26350 15314
rect 26402 15262 26686 15314
rect 26738 15262 26740 15314
rect 26348 15260 26740 15262
rect 26348 15250 26404 15260
rect 26684 15250 26740 15260
rect 26796 14868 26852 15484
rect 27020 15474 27076 15484
rect 26908 15314 26964 15326
rect 26908 15262 26910 15314
rect 26962 15262 26964 15314
rect 26908 15204 26964 15262
rect 26908 15138 26964 15148
rect 27244 15314 27300 15326
rect 27244 15262 27246 15314
rect 27298 15262 27300 15314
rect 25340 14532 25396 14542
rect 25228 14530 25396 14532
rect 25228 14478 25342 14530
rect 25394 14478 25396 14530
rect 25228 14476 25396 14478
rect 24556 14466 24612 14476
rect 25004 14466 25060 14476
rect 25340 14466 25396 14476
rect 25676 14530 25732 14588
rect 26460 14812 26852 14868
rect 26460 14642 26516 14812
rect 26460 14590 26462 14642
rect 26514 14590 26516 14642
rect 26460 14578 26516 14590
rect 25676 14478 25678 14530
rect 25730 14478 25732 14530
rect 25228 14306 25284 14318
rect 25228 14254 25230 14306
rect 25282 14254 25284 14306
rect 25228 12852 25284 14254
rect 25676 13076 25732 14478
rect 26012 14028 26516 14084
rect 25676 13010 25732 13020
rect 25788 13748 25844 13758
rect 26012 13748 26068 14028
rect 26460 13970 26516 14028
rect 26460 13918 26462 13970
rect 26514 13918 26516 13970
rect 26460 13906 26516 13918
rect 27244 13970 27300 15262
rect 27244 13918 27246 13970
rect 27298 13918 27300 13970
rect 27244 13906 27300 13918
rect 27468 14420 27524 14430
rect 27468 13970 27524 14364
rect 27468 13918 27470 13970
rect 27522 13918 27524 13970
rect 27468 13906 27524 13918
rect 25788 13746 26068 13748
rect 25788 13694 25790 13746
rect 25842 13694 26068 13746
rect 25788 13692 26068 13694
rect 26124 13858 26180 13870
rect 26124 13806 26126 13858
rect 26178 13806 26180 13858
rect 25788 13076 25844 13692
rect 25900 13076 25956 13086
rect 25788 13074 25956 13076
rect 25788 13022 25902 13074
rect 25954 13022 25956 13074
rect 25788 13020 25956 13022
rect 25788 12852 25844 13020
rect 25900 13010 25956 13020
rect 25228 12796 25844 12852
rect 21196 8372 21476 8428
rect 24444 8372 24612 8428
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 21420 3554 21476 8372
rect 21420 3502 21422 3554
rect 21474 3502 21476 3554
rect 21420 3490 21476 3502
rect 21532 3668 21588 3678
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 21532 800 21588 3612
rect 22428 3668 22484 3678
rect 22428 3574 22484 3612
rect 24220 3668 24276 3678
rect 24220 800 24276 3612
rect 24556 3554 24612 8372
rect 25788 4338 25844 12796
rect 25788 4286 25790 4338
rect 25842 4286 25844 4338
rect 25788 4274 25844 4286
rect 25564 3668 25620 3678
rect 25564 3574 25620 3612
rect 24556 3502 24558 3554
rect 24610 3502 24612 3554
rect 24556 3490 24612 3502
rect 26124 3556 26180 13806
rect 26796 13860 26852 13870
rect 26796 13766 26852 13804
rect 27580 13858 27636 15708
rect 28028 15316 28084 15326
rect 28140 15316 28196 16158
rect 28476 15428 28532 18396
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 40012 17778 40068 17790
rect 40012 17726 40014 17778
rect 40066 17726 40068 17778
rect 29932 17668 29988 17678
rect 29932 16770 29988 17612
rect 37660 17668 37716 17678
rect 37660 17574 37716 17612
rect 40012 17556 40068 17726
rect 40012 17490 40068 17500
rect 29932 16718 29934 16770
rect 29986 16718 29988 16770
rect 29932 16706 29988 16718
rect 37660 16882 37716 16894
rect 37660 16830 37662 16882
rect 37714 16830 37716 16882
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 30828 16100 30884 16110
rect 28700 15428 28756 15438
rect 28476 15426 28756 15428
rect 28476 15374 28702 15426
rect 28754 15374 28756 15426
rect 28476 15372 28756 15374
rect 28700 15362 28756 15372
rect 28028 15314 28196 15316
rect 28028 15262 28030 15314
rect 28082 15262 28196 15314
rect 28028 15260 28196 15262
rect 28028 15250 28084 15260
rect 30828 15204 30884 16044
rect 30828 15110 30884 15148
rect 37660 15204 37716 16830
rect 40012 16884 40068 16894
rect 40012 16770 40068 16828
rect 40012 16718 40014 16770
rect 40066 16718 40068 16770
rect 40012 16706 40068 16718
rect 37660 15138 37716 15148
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 28588 14642 28644 14654
rect 28588 14590 28590 14642
rect 28642 14590 28644 14642
rect 28588 14420 28644 14590
rect 29260 14644 29316 14654
rect 29260 14550 29316 14588
rect 40012 14642 40068 14654
rect 40012 14590 40014 14642
rect 40066 14590 40068 14642
rect 37660 14532 37716 14542
rect 37660 14438 37716 14476
rect 28588 14354 28644 14364
rect 40012 14196 40068 14590
rect 40012 14130 40068 14140
rect 27580 13806 27582 13858
rect 27634 13806 27636 13858
rect 27580 13794 27636 13806
rect 28700 13860 28756 13870
rect 26460 13076 26516 13086
rect 26460 12982 26516 13020
rect 28700 4338 28756 13804
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 28700 4286 28702 4338
rect 28754 4286 28756 4338
rect 28700 4274 28756 4286
rect 26796 4114 26852 4126
rect 27132 4116 27188 4126
rect 26796 4062 26798 4114
rect 26850 4062 26852 4114
rect 26124 3490 26180 3500
rect 26236 3668 26292 3678
rect 25564 3444 25620 3454
rect 25564 800 25620 3388
rect 26236 800 26292 3612
rect 26796 3444 26852 4062
rect 26796 3378 26852 3388
rect 26908 4060 27132 4116
rect 26908 800 26964 4060
rect 27132 4050 27188 4060
rect 29708 4116 29764 4126
rect 29708 4022 29764 4060
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 29372 3668 29428 3678
rect 29372 3574 29428 3612
rect 28588 3556 28644 3566
rect 28588 3462 28644 3500
rect 21504 0 21616 800
rect 24192 0 24304 800
rect 25536 0 25648 800
rect 26208 0 26320 800
rect 26880 0 26992 800
<< via2 >>
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 22876 38220 22932 38276
rect 20188 37436 20244 37492
rect 21420 37490 21476 37492
rect 21420 37438 21422 37490
rect 21422 37438 21474 37490
rect 21474 37438 21476 37490
rect 21420 37436 21476 37438
rect 18060 36988 18116 37044
rect 18844 36988 18900 37044
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 4172 27580 4228 27636
rect 1932 25564 1988 25620
rect 2044 24892 2100 24948
rect 1932 23548 1988 23604
rect 1932 19794 1988 19796
rect 1932 19742 1934 19794
rect 1934 19742 1986 19794
rect 1986 19742 1988 19794
rect 1932 19740 1988 19742
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 16044 27074 16100 27076
rect 16044 27022 16046 27074
rect 16046 27022 16098 27074
rect 16098 27022 16100 27074
rect 16044 27020 16100 27022
rect 4284 26290 4340 26292
rect 4284 26238 4286 26290
rect 4286 26238 4338 26290
rect 4338 26238 4340 26290
rect 4284 26236 4340 26238
rect 12796 26236 12852 26292
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 18172 27746 18228 27748
rect 18172 27694 18174 27746
rect 18174 27694 18226 27746
rect 18226 27694 18228 27746
rect 18172 27692 18228 27694
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 23548 36652 23604 36708
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 20076 27692 20132 27748
rect 23436 28476 23492 28532
rect 17388 27020 17444 27076
rect 12796 25340 12852 25396
rect 14252 25564 14308 25620
rect 4284 25228 4340 25284
rect 11564 25228 11620 25284
rect 13692 24834 13748 24836
rect 13692 24782 13694 24834
rect 13694 24782 13746 24834
rect 13746 24782 13748 24834
rect 13692 24780 13748 24782
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 4284 23938 4340 23940
rect 4284 23886 4286 23938
rect 4286 23886 4338 23938
rect 4338 23886 4340 23938
rect 4284 23884 4340 23886
rect 12124 24050 12180 24052
rect 12124 23998 12126 24050
rect 12126 23998 12178 24050
rect 12178 23998 12180 24050
rect 12124 23996 12180 23998
rect 13580 24050 13636 24052
rect 13580 23998 13582 24050
rect 13582 23998 13634 24050
rect 13634 23998 13636 24050
rect 13580 23996 13636 23998
rect 9996 23660 10052 23716
rect 12908 23938 12964 23940
rect 12908 23886 12910 23938
rect 12910 23886 12962 23938
rect 12962 23886 12964 23938
rect 12908 23884 12964 23886
rect 13804 23826 13860 23828
rect 13804 23774 13806 23826
rect 13806 23774 13858 23826
rect 13858 23774 13860 23826
rect 13804 23772 13860 23774
rect 13580 23324 13636 23380
rect 14028 23660 14084 23716
rect 14364 25282 14420 25284
rect 14364 25230 14366 25282
rect 14366 25230 14418 25282
rect 14418 25230 14420 25282
rect 14364 25228 14420 25230
rect 14476 25116 14532 25172
rect 14924 24834 14980 24836
rect 14924 24782 14926 24834
rect 14926 24782 14978 24834
rect 14978 24782 14980 24834
rect 14924 24780 14980 24782
rect 14364 23884 14420 23940
rect 14700 23938 14756 23940
rect 14700 23886 14702 23938
rect 14702 23886 14754 23938
rect 14754 23886 14756 23938
rect 14700 23884 14756 23886
rect 14364 23378 14420 23380
rect 14364 23326 14366 23378
rect 14366 23326 14418 23378
rect 14418 23326 14420 23378
rect 14364 23324 14420 23326
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 13244 22092 13300 22148
rect 11116 21474 11172 21476
rect 11116 21422 11118 21474
rect 11118 21422 11170 21474
rect 11170 21422 11172 21474
rect 11116 21420 11172 21422
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 14252 22428 14308 22484
rect 14700 23154 14756 23156
rect 14700 23102 14702 23154
rect 14702 23102 14754 23154
rect 14754 23102 14756 23154
rect 14700 23100 14756 23102
rect 14476 22316 14532 22372
rect 19516 26962 19572 26964
rect 19516 26910 19518 26962
rect 19518 26910 19570 26962
rect 19570 26910 19572 26962
rect 19516 26908 19572 26910
rect 17500 26402 17556 26404
rect 17500 26350 17502 26402
rect 17502 26350 17554 26402
rect 17554 26350 17556 26402
rect 17500 26348 17556 26350
rect 18396 26402 18452 26404
rect 18396 26350 18398 26402
rect 18398 26350 18450 26402
rect 18450 26350 18452 26402
rect 18396 26348 18452 26350
rect 19404 26796 19460 26852
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 16716 26124 16772 26180
rect 16044 25506 16100 25508
rect 16044 25454 16046 25506
rect 16046 25454 16098 25506
rect 16098 25454 16100 25506
rect 16044 25452 16100 25454
rect 15932 25394 15988 25396
rect 15932 25342 15934 25394
rect 15934 25342 15986 25394
rect 15986 25342 15988 25394
rect 15932 25340 15988 25342
rect 15820 25228 15876 25284
rect 15596 24780 15652 24836
rect 15036 23772 15092 23828
rect 14924 22370 14980 22372
rect 14924 22318 14926 22370
rect 14926 22318 14978 22370
rect 14978 22318 14980 22370
rect 14924 22316 14980 22318
rect 16716 24556 16772 24612
rect 17500 26124 17556 26180
rect 19180 26178 19236 26180
rect 19180 26126 19182 26178
rect 19182 26126 19234 26178
rect 19234 26126 19236 26178
rect 19180 26124 19236 26126
rect 18844 25452 18900 25508
rect 18060 25228 18116 25284
rect 20076 26178 20132 26180
rect 20076 26126 20078 26178
rect 20078 26126 20130 26178
rect 20130 26126 20132 26178
rect 20076 26124 20132 26126
rect 19180 25228 19236 25284
rect 19628 25788 19684 25844
rect 17388 24556 17444 24612
rect 20300 26908 20356 26964
rect 22540 27020 22596 27076
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 25564 38274 25620 38276
rect 25564 38222 25566 38274
rect 25566 38222 25618 38274
rect 25618 38222 25620 38274
rect 25564 38220 25620 38222
rect 24220 37436 24276 37492
rect 24108 28476 24164 28532
rect 23436 27074 23492 27076
rect 23436 27022 23438 27074
rect 23438 27022 23490 27074
rect 23490 27022 23492 27074
rect 23436 27020 23492 27022
rect 21308 26796 21364 26852
rect 20412 26124 20468 26180
rect 20860 25900 20916 25956
rect 21196 25900 21252 25956
rect 20188 25788 20244 25844
rect 19628 25452 19684 25508
rect 20860 25228 20916 25284
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 15708 23154 15764 23156
rect 15708 23102 15710 23154
rect 15710 23102 15762 23154
rect 15762 23102 15764 23154
rect 15708 23100 15764 23102
rect 14700 21756 14756 21812
rect 13468 20524 13524 20580
rect 13916 21586 13972 21588
rect 13916 21534 13918 21586
rect 13918 21534 13970 21586
rect 13970 21534 13972 21586
rect 13916 21532 13972 21534
rect 13916 20524 13972 20580
rect 14252 20578 14308 20580
rect 14252 20526 14254 20578
rect 14254 20526 14306 20578
rect 14306 20526 14308 20578
rect 14252 20524 14308 20526
rect 15148 21756 15204 21812
rect 15932 22204 15988 22260
rect 15708 21756 15764 21812
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 16156 22482 16212 22484
rect 16156 22430 16158 22482
rect 16158 22430 16210 22482
rect 16210 22430 16212 22482
rect 16156 22428 16212 22430
rect 17388 22316 17444 22372
rect 16380 22092 16436 22148
rect 16268 21756 16324 21812
rect 14924 21362 14980 21364
rect 14924 21310 14926 21362
rect 14926 21310 14978 21362
rect 14978 21310 14980 21362
rect 14924 21308 14980 21310
rect 15708 21420 15764 21476
rect 14700 20972 14756 21028
rect 9996 20076 10052 20132
rect 4284 20018 4340 20020
rect 4284 19966 4286 20018
rect 4286 19966 4338 20018
rect 4338 19966 4340 20018
rect 4284 19964 4340 19966
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 13692 20130 13748 20132
rect 13692 20078 13694 20130
rect 13694 20078 13746 20130
rect 13746 20078 13748 20130
rect 13692 20076 13748 20078
rect 16268 21026 16324 21028
rect 16268 20974 16270 21026
rect 16270 20974 16322 21026
rect 16322 20974 16324 21026
rect 16268 20972 16324 20974
rect 16940 22258 16996 22260
rect 16940 22206 16942 22258
rect 16942 22206 16994 22258
rect 16994 22206 16996 22258
rect 16940 22204 16996 22206
rect 16828 22146 16884 22148
rect 16828 22094 16830 22146
rect 16830 22094 16882 22146
rect 16882 22094 16884 22146
rect 16828 22092 16884 22094
rect 13356 19404 13412 19460
rect 12124 19122 12180 19124
rect 12124 19070 12126 19122
rect 12126 19070 12178 19122
rect 12178 19070 12180 19122
rect 12124 19068 12180 19070
rect 4172 18956 4228 19012
rect 12124 18508 12180 18564
rect 4284 18450 4340 18452
rect 4284 18398 4286 18450
rect 4286 18398 4338 18450
rect 4338 18398 4340 18450
rect 4284 18396 4340 18398
rect 9996 18284 10052 18340
rect 1932 18226 1988 18228
rect 1932 18174 1934 18226
rect 1934 18174 1986 18226
rect 1986 18174 1988 18226
rect 1932 18172 1988 18174
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 13804 19404 13860 19460
rect 15260 19458 15316 19460
rect 15260 19406 15262 19458
rect 15262 19406 15314 19458
rect 15314 19406 15316 19458
rect 15260 19404 15316 19406
rect 15932 20578 15988 20580
rect 15932 20526 15934 20578
rect 15934 20526 15986 20578
rect 15986 20526 15988 20578
rect 15932 20524 15988 20526
rect 16604 20802 16660 20804
rect 16604 20750 16606 20802
rect 16606 20750 16658 20802
rect 16658 20750 16660 20802
rect 16604 20748 16660 20750
rect 16492 20636 16548 20692
rect 16380 20076 16436 20132
rect 17724 22146 17780 22148
rect 17724 22094 17726 22146
rect 17726 22094 17778 22146
rect 17778 22094 17780 22146
rect 17724 22092 17780 22094
rect 17612 21474 17668 21476
rect 17612 21422 17614 21474
rect 17614 21422 17666 21474
rect 17666 21422 17668 21474
rect 17612 21420 17668 21422
rect 18396 21532 18452 21588
rect 17164 20690 17220 20692
rect 17164 20638 17166 20690
rect 17166 20638 17218 20690
rect 17218 20638 17220 20690
rect 17164 20636 17220 20638
rect 17276 20748 17332 20804
rect 13804 19234 13860 19236
rect 13804 19182 13806 19234
rect 13806 19182 13858 19234
rect 13858 19182 13860 19234
rect 13804 19180 13860 19182
rect 13580 19122 13636 19124
rect 13580 19070 13582 19122
rect 13582 19070 13634 19122
rect 13634 19070 13636 19122
rect 13580 19068 13636 19070
rect 15372 19234 15428 19236
rect 15372 19182 15374 19234
rect 15374 19182 15426 19234
rect 15426 19182 15428 19234
rect 15372 19180 15428 19182
rect 13468 18562 13524 18564
rect 13468 18510 13470 18562
rect 13470 18510 13522 18562
rect 13522 18510 13524 18562
rect 13468 18508 13524 18510
rect 14140 18450 14196 18452
rect 14140 18398 14142 18450
rect 14142 18398 14194 18450
rect 14194 18398 14196 18450
rect 14140 18396 14196 18398
rect 15036 18396 15092 18452
rect 14588 18338 14644 18340
rect 14588 18286 14590 18338
rect 14590 18286 14642 18338
rect 14642 18286 14644 18338
rect 14588 18284 14644 18286
rect 15148 18060 15204 18116
rect 12908 17666 12964 17668
rect 12908 17614 12910 17666
rect 12910 17614 12962 17666
rect 12962 17614 12964 17666
rect 12908 17612 12964 17614
rect 13580 17612 13636 17668
rect 16604 19180 16660 19236
rect 16828 19292 16884 19348
rect 16604 18620 16660 18676
rect 18284 20914 18340 20916
rect 18284 20862 18286 20914
rect 18286 20862 18338 20914
rect 18338 20862 18340 20914
rect 18284 20860 18340 20862
rect 18172 20748 18228 20804
rect 18060 20524 18116 20580
rect 17388 20018 17444 20020
rect 17388 19966 17390 20018
rect 17390 19966 17442 20018
rect 17442 19966 17444 20018
rect 17388 19964 17444 19966
rect 17724 20130 17780 20132
rect 17724 20078 17726 20130
rect 17726 20078 17778 20130
rect 17778 20078 17780 20130
rect 17724 20076 17780 20078
rect 17724 19346 17780 19348
rect 17724 19294 17726 19346
rect 17726 19294 17778 19346
rect 17778 19294 17780 19346
rect 17724 19292 17780 19294
rect 18620 21308 18676 21364
rect 18732 20748 18788 20804
rect 19292 22146 19348 22148
rect 19292 22094 19294 22146
rect 19294 22094 19346 22146
rect 19346 22094 19348 22146
rect 19292 22092 19348 22094
rect 19404 21756 19460 21812
rect 18956 20412 19012 20468
rect 18956 20130 19012 20132
rect 18956 20078 18958 20130
rect 18958 20078 19010 20130
rect 19010 20078 19012 20130
rect 18956 20076 19012 20078
rect 18844 20018 18900 20020
rect 18844 19966 18846 20018
rect 18846 19966 18898 20018
rect 18898 19966 18900 20018
rect 18844 19964 18900 19966
rect 17052 19068 17108 19124
rect 17276 18844 17332 18900
rect 16380 18172 16436 18228
rect 15260 17612 15316 17668
rect 15708 17666 15764 17668
rect 15708 17614 15710 17666
rect 15710 17614 15762 17666
rect 15762 17614 15764 17666
rect 15708 17612 15764 17614
rect 14476 16994 14532 16996
rect 14476 16942 14478 16994
rect 14478 16942 14530 16994
rect 14530 16942 14532 16994
rect 14476 16940 14532 16942
rect 15484 16940 15540 16996
rect 13804 16882 13860 16884
rect 13804 16830 13806 16882
rect 13806 16830 13858 16882
rect 13858 16830 13860 16882
rect 13804 16828 13860 16830
rect 17388 18226 17444 18228
rect 17388 18174 17390 18226
rect 17390 18174 17442 18226
rect 17442 18174 17444 18226
rect 17388 18172 17444 18174
rect 18284 19628 18340 19684
rect 19404 20412 19460 20468
rect 19404 19740 19460 19796
rect 19404 19404 19460 19460
rect 18284 18844 18340 18900
rect 18396 19292 18452 19348
rect 17948 18620 18004 18676
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 20076 20524 20132 20580
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 18956 19122 19012 19124
rect 18956 19070 18958 19122
rect 18958 19070 19010 19122
rect 19010 19070 19012 19122
rect 18956 19068 19012 19070
rect 19628 19068 19684 19124
rect 18620 18172 18676 18228
rect 19292 17724 19348 17780
rect 17724 17388 17780 17444
rect 17500 16882 17556 16884
rect 17500 16830 17502 16882
rect 17502 16830 17554 16882
rect 17554 16830 17556 16882
rect 17500 16828 17556 16830
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 20076 19852 20132 19908
rect 19964 19122 20020 19124
rect 19964 19070 19966 19122
rect 19966 19070 20018 19122
rect 20018 19070 20020 19122
rect 19964 19068 20020 19070
rect 20748 23378 20804 23380
rect 20748 23326 20750 23378
rect 20750 23326 20802 23378
rect 20802 23326 20804 23378
rect 20748 23324 20804 23326
rect 21420 25228 21476 25284
rect 20972 23324 21028 23380
rect 20412 20802 20468 20804
rect 20412 20750 20414 20802
rect 20414 20750 20466 20802
rect 20466 20750 20468 20802
rect 20412 20748 20468 20750
rect 20636 19852 20692 19908
rect 20300 19628 20356 19684
rect 20524 19740 20580 19796
rect 20524 19234 20580 19236
rect 20524 19182 20526 19234
rect 20526 19182 20578 19234
rect 20578 19182 20580 19234
rect 20524 19180 20580 19182
rect 19740 19010 19796 19012
rect 19740 18958 19742 19010
rect 19742 18958 19794 19010
rect 19794 18958 19796 19010
rect 19740 18956 19796 18958
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 20636 18620 20692 18676
rect 21308 22930 21364 22932
rect 21308 22878 21310 22930
rect 21310 22878 21362 22930
rect 21362 22878 21364 22930
rect 21308 22876 21364 22878
rect 21980 26684 22036 26740
rect 21644 25506 21700 25508
rect 21644 25454 21646 25506
rect 21646 25454 21698 25506
rect 21698 25454 21700 25506
rect 21644 25452 21700 25454
rect 23660 26962 23716 26964
rect 23660 26910 23662 26962
rect 23662 26910 23714 26962
rect 23714 26910 23716 26962
rect 23660 26908 23716 26910
rect 22652 26684 22708 26740
rect 23324 26178 23380 26180
rect 23324 26126 23326 26178
rect 23326 26126 23378 26178
rect 23378 26126 23380 26178
rect 23324 26124 23380 26126
rect 26236 37490 26292 37492
rect 26236 37438 26238 37490
rect 26238 37438 26290 37490
rect 26290 37438 26292 37490
rect 26236 37436 26292 37438
rect 24780 36706 24836 36708
rect 24780 36654 24782 36706
rect 24782 36654 24834 36706
rect 24834 36654 24836 36706
rect 24780 36652 24836 36654
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 25340 26908 25396 26964
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 25452 26796 25508 26852
rect 24556 26124 24612 26180
rect 22876 24946 22932 24948
rect 22876 24894 22878 24946
rect 22878 24894 22930 24946
rect 22930 24894 22932 24946
rect 22876 24892 22932 24894
rect 25004 25228 25060 25284
rect 32060 26236 32116 26292
rect 25564 25228 25620 25284
rect 26012 25228 26068 25284
rect 23436 24892 23492 24948
rect 25452 24834 25508 24836
rect 25452 24782 25454 24834
rect 25454 24782 25506 24834
rect 25506 24782 25508 24834
rect 25452 24780 25508 24782
rect 21756 22930 21812 22932
rect 21756 22878 21758 22930
rect 21758 22878 21810 22930
rect 21810 22878 21812 22930
rect 21756 22876 21812 22878
rect 25900 24722 25956 24724
rect 25900 24670 25902 24722
rect 25902 24670 25954 24722
rect 25954 24670 25956 24722
rect 25900 24668 25956 24670
rect 25788 24610 25844 24612
rect 25788 24558 25790 24610
rect 25790 24558 25842 24610
rect 25842 24558 25844 24610
rect 25788 24556 25844 24558
rect 25676 24444 25732 24500
rect 21980 21644 22036 21700
rect 21196 20860 21252 20916
rect 22092 20860 22148 20916
rect 21980 20636 22036 20692
rect 22764 22428 22820 22484
rect 22316 21756 22372 21812
rect 23212 21868 23268 21924
rect 22876 21586 22932 21588
rect 22876 21534 22878 21586
rect 22878 21534 22930 21586
rect 22930 21534 22932 21586
rect 22876 21532 22932 21534
rect 22652 20748 22708 20804
rect 22204 20524 22260 20580
rect 21420 20412 21476 20468
rect 22988 20578 23044 20580
rect 22988 20526 22990 20578
rect 22990 20526 23042 20578
rect 23042 20526 23044 20578
rect 22988 20524 23044 20526
rect 22876 20412 22932 20468
rect 21420 20076 21476 20132
rect 21308 19628 21364 19684
rect 20860 18396 20916 18452
rect 21868 19010 21924 19012
rect 21868 18958 21870 19010
rect 21870 18958 21922 19010
rect 21922 18958 21924 19010
rect 21868 18956 21924 18958
rect 20748 18060 20804 18116
rect 21532 18620 21588 18676
rect 21868 18620 21924 18676
rect 21756 18172 21812 18228
rect 22428 18620 22484 18676
rect 22764 18956 22820 19012
rect 22316 18508 22372 18564
rect 22876 18508 22932 18564
rect 22540 18450 22596 18452
rect 22540 18398 22542 18450
rect 22542 18398 22594 18450
rect 22594 18398 22596 18450
rect 22540 18396 22596 18398
rect 22988 18396 23044 18452
rect 25452 21756 25508 21812
rect 23548 21644 23604 21700
rect 23324 21420 23380 21476
rect 23324 20802 23380 20804
rect 23324 20750 23326 20802
rect 23326 20750 23378 20802
rect 23378 20750 23380 20802
rect 23324 20748 23380 20750
rect 23436 20636 23492 20692
rect 24220 21420 24276 21476
rect 23884 20524 23940 20580
rect 23660 19852 23716 19908
rect 23772 19458 23828 19460
rect 23772 19406 23774 19458
rect 23774 19406 23826 19458
rect 23826 19406 23828 19458
rect 23772 19404 23828 19406
rect 24444 19122 24500 19124
rect 24444 19070 24446 19122
rect 24446 19070 24498 19122
rect 24498 19070 24500 19122
rect 24444 19068 24500 19070
rect 23436 18620 23492 18676
rect 23884 18620 23940 18676
rect 24220 18674 24276 18676
rect 24220 18622 24222 18674
rect 24222 18622 24274 18674
rect 24274 18622 24276 18674
rect 24220 18620 24276 18622
rect 23996 18562 24052 18564
rect 23996 18510 23998 18562
rect 23998 18510 24050 18562
rect 24050 18510 24052 18562
rect 23996 18508 24052 18510
rect 21980 18338 22036 18340
rect 21980 18286 21982 18338
rect 21982 18286 22034 18338
rect 22034 18286 22036 18338
rect 21980 18284 22036 18286
rect 23212 18284 23268 18340
rect 23660 18396 23716 18452
rect 20412 17836 20468 17892
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 18396 16044 18452 16100
rect 18956 16098 19012 16100
rect 18956 16046 18958 16098
rect 18958 16046 19010 16098
rect 19010 16046 19012 16098
rect 18956 16044 19012 16046
rect 23548 18172 23604 18228
rect 22204 17778 22260 17780
rect 22204 17726 22206 17778
rect 22206 17726 22258 17778
rect 22258 17726 22260 17778
rect 22204 17724 22260 17726
rect 19852 16098 19908 16100
rect 19852 16046 19854 16098
rect 19854 16046 19906 16098
rect 19906 16046 19908 16098
rect 19852 16044 19908 16046
rect 20076 16098 20132 16100
rect 20076 16046 20078 16098
rect 20078 16046 20130 16098
rect 20130 16046 20132 16098
rect 20076 16044 20132 16046
rect 18508 15986 18564 15988
rect 18508 15934 18510 15986
rect 18510 15934 18562 15986
rect 18562 15934 18564 15986
rect 18508 15932 18564 15934
rect 17500 14588 17556 14644
rect 19068 15820 19124 15876
rect 19964 15874 20020 15876
rect 19964 15822 19966 15874
rect 19966 15822 20018 15874
rect 20018 15822 20020 15874
rect 19964 15820 20020 15822
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 18396 14588 18452 14644
rect 21756 17106 21812 17108
rect 21756 17054 21758 17106
rect 21758 17054 21810 17106
rect 21810 17054 21812 17106
rect 21756 17052 21812 17054
rect 23772 17052 23828 17108
rect 23884 16716 23940 16772
rect 23884 16044 23940 16100
rect 21644 15314 21700 15316
rect 21644 15262 21646 15314
rect 21646 15262 21698 15314
rect 21698 15262 21700 15314
rect 21644 15260 21700 15262
rect 22988 15260 23044 15316
rect 20860 14642 20916 14644
rect 20860 14590 20862 14642
rect 20862 14590 20914 14642
rect 20914 14590 20916 14642
rect 20860 14588 20916 14590
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 21420 14642 21476 14644
rect 21420 14590 21422 14642
rect 21422 14590 21474 14642
rect 21474 14590 21476 14642
rect 21420 14588 21476 14590
rect 24220 15372 24276 15428
rect 24780 19010 24836 19012
rect 24780 18958 24782 19010
rect 24782 18958 24834 19010
rect 24834 18958 24836 19010
rect 24780 18956 24836 18958
rect 25564 22204 25620 22260
rect 25788 21644 25844 21700
rect 25452 21586 25508 21588
rect 25452 21534 25454 21586
rect 25454 21534 25506 21586
rect 25506 21534 25508 21586
rect 25452 21532 25508 21534
rect 25564 21362 25620 21364
rect 25564 21310 25566 21362
rect 25566 21310 25618 21362
rect 25618 21310 25620 21362
rect 25564 21308 25620 21310
rect 25340 20524 25396 20580
rect 25452 20188 25508 20244
rect 25228 19852 25284 19908
rect 24892 17052 24948 17108
rect 24556 16716 24612 16772
rect 25788 21420 25844 21476
rect 27020 25452 27076 25508
rect 27804 25452 27860 25508
rect 26908 24892 26964 24948
rect 26348 24780 26404 24836
rect 26236 24722 26292 24724
rect 26236 24670 26238 24722
rect 26238 24670 26290 24722
rect 26290 24670 26292 24722
rect 26236 24668 26292 24670
rect 27580 24834 27636 24836
rect 27580 24782 27582 24834
rect 27582 24782 27634 24834
rect 27634 24782 27636 24834
rect 27580 24780 27636 24782
rect 26908 24722 26964 24724
rect 26908 24670 26910 24722
rect 26910 24670 26962 24722
rect 26962 24670 26964 24722
rect 26908 24668 26964 24670
rect 26236 24444 26292 24500
rect 26348 23826 26404 23828
rect 26348 23774 26350 23826
rect 26350 23774 26402 23826
rect 26402 23774 26404 23826
rect 26348 23772 26404 23774
rect 26012 22482 26068 22484
rect 26012 22430 26014 22482
rect 26014 22430 26066 22482
rect 26066 22430 26068 22482
rect 26012 22428 26068 22430
rect 26124 22316 26180 22372
rect 27244 24556 27300 24612
rect 27692 24556 27748 24612
rect 26460 22316 26516 22372
rect 26796 22428 26852 22484
rect 26348 21698 26404 21700
rect 26348 21646 26350 21698
rect 26350 21646 26402 21698
rect 26402 21646 26404 21698
rect 26348 21644 26404 21646
rect 26124 21420 26180 21476
rect 26460 21308 26516 21364
rect 25228 18396 25284 18452
rect 25228 17836 25284 17892
rect 25564 19010 25620 19012
rect 25564 18958 25566 19010
rect 25566 18958 25618 19010
rect 25618 18958 25620 19010
rect 25564 18956 25620 18958
rect 25228 17442 25284 17444
rect 25228 17390 25230 17442
rect 25230 17390 25282 17442
rect 25282 17390 25284 17442
rect 25228 17388 25284 17390
rect 25116 15372 25172 15428
rect 25228 15820 25284 15876
rect 25564 18620 25620 18676
rect 25452 18060 25508 18116
rect 26348 19068 26404 19124
rect 26236 18562 26292 18564
rect 26236 18510 26238 18562
rect 26238 18510 26290 18562
rect 26290 18510 26292 18562
rect 26236 18508 26292 18510
rect 26012 18450 26068 18452
rect 26012 18398 26014 18450
rect 26014 18398 26066 18450
rect 26066 18398 26068 18450
rect 26012 18396 26068 18398
rect 27804 24444 27860 24500
rect 27804 23884 27860 23940
rect 28252 25394 28308 25396
rect 28252 25342 28254 25394
rect 28254 25342 28306 25394
rect 28306 25342 28308 25394
rect 28252 25340 28308 25342
rect 28364 25228 28420 25284
rect 29596 25564 29652 25620
rect 29148 25228 29204 25284
rect 37660 26290 37716 26292
rect 37660 26238 37662 26290
rect 37662 26238 37714 26290
rect 37714 26238 37716 26290
rect 37660 26236 37716 26238
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 32060 25618 32116 25620
rect 32060 25566 32062 25618
rect 32062 25566 32114 25618
rect 32114 25566 32116 25618
rect 32060 25564 32116 25566
rect 37660 25506 37716 25508
rect 37660 25454 37662 25506
rect 37662 25454 37714 25506
rect 37714 25454 37716 25506
rect 37660 25452 37716 25454
rect 40012 26236 40068 26292
rect 39900 25564 39956 25620
rect 37884 25228 37940 25284
rect 40012 24892 40068 24948
rect 28140 24668 28196 24724
rect 28476 24668 28532 24724
rect 28700 24556 28756 24612
rect 29260 24722 29316 24724
rect 29260 24670 29262 24722
rect 29262 24670 29314 24722
rect 29314 24670 29316 24722
rect 29260 24668 29316 24670
rect 29820 24668 29876 24724
rect 28924 24444 28980 24500
rect 27692 22316 27748 22372
rect 28252 22370 28308 22372
rect 28252 22318 28254 22370
rect 28254 22318 28306 22370
rect 28306 22318 28308 22370
rect 28252 22316 28308 22318
rect 28140 22258 28196 22260
rect 28140 22206 28142 22258
rect 28142 22206 28194 22258
rect 28194 22206 28196 22258
rect 28140 22204 28196 22206
rect 28028 21868 28084 21924
rect 27132 21698 27188 21700
rect 27132 21646 27134 21698
rect 27134 21646 27186 21698
rect 27186 21646 27188 21698
rect 27132 21644 27188 21646
rect 26908 21586 26964 21588
rect 26908 21534 26910 21586
rect 26910 21534 26962 21586
rect 26962 21534 26964 21586
rect 26908 21532 26964 21534
rect 26796 20188 26852 20244
rect 27580 20972 27636 21028
rect 26908 20018 26964 20020
rect 26908 19966 26910 20018
rect 26910 19966 26962 20018
rect 26962 19966 26964 20018
rect 26908 19964 26964 19966
rect 26908 19180 26964 19236
rect 26348 17612 26404 17668
rect 26460 17724 26516 17780
rect 26012 17388 26068 17444
rect 26908 17276 26964 17332
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 30156 22428 30212 22484
rect 29932 22258 29988 22260
rect 29932 22206 29934 22258
rect 29934 22206 29986 22258
rect 29986 22206 29988 22258
rect 29932 22204 29988 22206
rect 32060 22482 32116 22484
rect 32060 22430 32062 22482
rect 32062 22430 32114 22482
rect 32114 22430 32116 22482
rect 32060 22428 32116 22430
rect 37660 22428 37716 22484
rect 40012 22204 40068 22260
rect 29036 20972 29092 21028
rect 37660 21586 37716 21588
rect 37660 21534 37662 21586
rect 37662 21534 37714 21586
rect 37714 21534 37716 21586
rect 37660 21532 37716 21534
rect 40012 21532 40068 21588
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 40012 20914 40068 20916
rect 40012 20862 40014 20914
rect 40014 20862 40066 20914
rect 40066 20862 40068 20914
rect 40012 20860 40068 20862
rect 29260 20578 29316 20580
rect 29260 20526 29262 20578
rect 29262 20526 29314 20578
rect 29314 20526 29316 20578
rect 29260 20524 29316 20526
rect 29708 20524 29764 20580
rect 28812 19964 28868 20020
rect 28028 19180 28084 19236
rect 28700 19740 28756 19796
rect 28140 19122 28196 19124
rect 28140 19070 28142 19122
rect 28142 19070 28194 19122
rect 28194 19070 28196 19122
rect 28140 19068 28196 19070
rect 28252 19010 28308 19012
rect 28252 18958 28254 19010
rect 28254 18958 28306 19010
rect 28306 18958 28308 19010
rect 28252 18956 28308 18958
rect 28028 18732 28084 18788
rect 29260 19852 29316 19908
rect 37660 20802 37716 20804
rect 37660 20750 37662 20802
rect 37662 20750 37714 20802
rect 37714 20750 37716 20802
rect 37660 20748 37716 20750
rect 30156 20130 30212 20132
rect 30156 20078 30158 20130
rect 30158 20078 30210 20130
rect 30210 20078 30212 20130
rect 30156 20076 30212 20078
rect 32060 19964 32116 20020
rect 30716 19906 30772 19908
rect 30716 19854 30718 19906
rect 30718 19854 30770 19906
rect 30770 19854 30772 19906
rect 30716 19852 30772 19854
rect 30156 19794 30212 19796
rect 30156 19742 30158 19794
rect 30158 19742 30210 19794
rect 30210 19742 30212 19794
rect 30156 19740 30212 19742
rect 37660 20018 37716 20020
rect 37660 19966 37662 20018
rect 37662 19966 37714 20018
rect 37714 19966 37716 20018
rect 37660 19964 37716 19966
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 40012 19516 40068 19572
rect 29932 19122 29988 19124
rect 29932 19070 29934 19122
rect 29934 19070 29986 19122
rect 29986 19070 29988 19122
rect 29932 19068 29988 19070
rect 27356 18562 27412 18564
rect 27356 18510 27358 18562
rect 27358 18510 27410 18562
rect 27410 18510 27412 18562
rect 27356 18508 27412 18510
rect 27580 18172 27636 18228
rect 27020 16882 27076 16884
rect 27020 16830 27022 16882
rect 27022 16830 27074 16882
rect 27074 16830 27076 16882
rect 27020 16828 27076 16830
rect 27132 16940 27188 16996
rect 27356 17052 27412 17108
rect 28364 17666 28420 17668
rect 28364 17614 28366 17666
rect 28366 17614 28418 17666
rect 28418 17614 28420 17666
rect 28364 17612 28420 17614
rect 27916 17554 27972 17556
rect 27916 17502 27918 17554
rect 27918 17502 27970 17554
rect 27970 17502 27972 17554
rect 27916 17500 27972 17502
rect 27692 17276 27748 17332
rect 27804 17442 27860 17444
rect 27804 17390 27806 17442
rect 27806 17390 27858 17442
rect 27858 17390 27860 17442
rect 27804 17388 27860 17390
rect 27580 16940 27636 16996
rect 27692 17052 27748 17108
rect 27692 16098 27748 16100
rect 27692 16046 27694 16098
rect 27694 16046 27746 16098
rect 27746 16046 27748 16098
rect 27692 16044 27748 16046
rect 26572 15932 26628 15988
rect 27244 15986 27300 15988
rect 27244 15934 27246 15986
rect 27246 15934 27298 15986
rect 27298 15934 27300 15986
rect 27244 15932 27300 15934
rect 25788 15820 25844 15876
rect 28140 16828 28196 16884
rect 26236 15426 26292 15428
rect 26236 15374 26238 15426
rect 26238 15374 26290 15426
rect 26290 15374 26292 15426
rect 26236 15372 26292 15374
rect 25340 15314 25396 15316
rect 25340 15262 25342 15314
rect 25342 15262 25394 15314
rect 25394 15262 25396 15314
rect 25340 15260 25396 15262
rect 25228 15148 25284 15204
rect 26908 15148 26964 15204
rect 25676 14588 25732 14644
rect 25676 13020 25732 13076
rect 27468 14364 27524 14420
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 21532 3612 21588 3668
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 22428 3666 22484 3668
rect 22428 3614 22430 3666
rect 22430 3614 22482 3666
rect 22482 3614 22484 3666
rect 22428 3612 22484 3614
rect 24220 3612 24276 3668
rect 25564 3666 25620 3668
rect 25564 3614 25566 3666
rect 25566 3614 25618 3666
rect 25618 3614 25620 3666
rect 25564 3612 25620 3614
rect 26796 13858 26852 13860
rect 26796 13806 26798 13858
rect 26798 13806 26850 13858
rect 26850 13806 26852 13858
rect 26796 13804 26852 13806
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 29932 17612 29988 17668
rect 37660 17666 37716 17668
rect 37660 17614 37662 17666
rect 37662 17614 37714 17666
rect 37714 17614 37716 17666
rect 37660 17612 37716 17614
rect 40012 17500 40068 17556
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 30828 16044 30884 16100
rect 30828 15202 30884 15204
rect 30828 15150 30830 15202
rect 30830 15150 30882 15202
rect 30882 15150 30884 15202
rect 30828 15148 30884 15150
rect 40012 16828 40068 16884
rect 37660 15148 37716 15204
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 29260 14642 29316 14644
rect 29260 14590 29262 14642
rect 29262 14590 29314 14642
rect 29314 14590 29316 14642
rect 29260 14588 29316 14590
rect 37660 14530 37716 14532
rect 37660 14478 37662 14530
rect 37662 14478 37714 14530
rect 37714 14478 37716 14530
rect 37660 14476 37716 14478
rect 28588 14364 28644 14420
rect 40012 14140 40068 14196
rect 28700 13804 28756 13860
rect 26460 13074 26516 13076
rect 26460 13022 26462 13074
rect 26462 13022 26514 13074
rect 26514 13022 26516 13074
rect 26460 13020 26516 13022
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 26124 3500 26180 3556
rect 26236 3612 26292 3668
rect 25564 3388 25620 3444
rect 26796 3388 26852 3444
rect 27132 4060 27188 4116
rect 29708 4114 29764 4116
rect 29708 4062 29710 4114
rect 29710 4062 29762 4114
rect 29762 4062 29764 4114
rect 29708 4060 29764 4062
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 29372 3666 29428 3668
rect 29372 3614 29374 3666
rect 29374 3614 29426 3666
rect 29426 3614 29428 3666
rect 29372 3612 29428 3614
rect 28588 3554 28644 3556
rect 28588 3502 28590 3554
rect 28590 3502 28642 3554
rect 28642 3502 28644 3554
rect 28588 3500 28644 3502
<< metal3 >>
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 22866 38220 22876 38276
rect 22932 38220 25564 38276
rect 25620 38220 25630 38276
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 20178 37436 20188 37492
rect 20244 37436 21420 37492
rect 21476 37436 21486 37492
rect 24210 37436 24220 37492
rect 24276 37436 26236 37492
rect 26292 37436 26302 37492
rect 18050 36988 18060 37044
rect 18116 36988 18844 37044
rect 18900 36988 18910 37044
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 23538 36652 23548 36708
rect 23604 36652 24780 36708
rect 24836 36652 24846 36708
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 23426 28476 23436 28532
rect 23492 28476 24108 28532
rect 24164 28476 24174 28532
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 18162 27692 18172 27748
rect 18228 27692 20076 27748
rect 20132 27692 20142 27748
rect 0 27636 800 27664
rect 0 27580 4172 27636
rect 4228 27580 4238 27636
rect 0 27552 800 27580
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 16034 27020 16044 27076
rect 16100 27020 17388 27076
rect 17444 27020 17454 27076
rect 22530 27020 22540 27076
rect 22596 27020 23436 27076
rect 23492 27020 23502 27076
rect 19506 26908 19516 26964
rect 19572 26908 20300 26964
rect 20356 26908 20366 26964
rect 23650 26908 23660 26964
rect 23716 26908 25340 26964
rect 25396 26908 25406 26964
rect 19394 26796 19404 26852
rect 19460 26796 21140 26852
rect 21298 26796 21308 26852
rect 21364 26796 25452 26852
rect 25508 26796 25518 26852
rect 21084 26740 21140 26796
rect 21084 26684 21980 26740
rect 22036 26684 22652 26740
rect 22708 26684 22718 26740
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 17490 26348 17500 26404
rect 17556 26348 18396 26404
rect 18452 26348 18462 26404
rect 41200 26292 42000 26320
rect 4274 26236 4284 26292
rect 4340 26236 12796 26292
rect 12852 26236 12862 26292
rect 32050 26236 32060 26292
rect 32116 26236 37660 26292
rect 37716 26236 37726 26292
rect 40002 26236 40012 26292
rect 40068 26236 42000 26292
rect 41200 26208 42000 26236
rect 16706 26124 16716 26180
rect 16772 26124 17500 26180
rect 17556 26124 17566 26180
rect 19170 26124 19180 26180
rect 19236 26124 20076 26180
rect 20132 26124 20412 26180
rect 20468 26124 20478 26180
rect 23314 26124 23324 26180
rect 23380 26124 24556 26180
rect 24612 26124 24622 26180
rect 20850 25900 20860 25956
rect 20916 25900 21196 25956
rect 21252 25900 21262 25956
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 19618 25788 19628 25844
rect 19684 25788 20188 25844
rect 20244 25788 20254 25844
rect 0 25620 800 25648
rect 41200 25620 42000 25648
rect 0 25564 1932 25620
rect 1988 25564 1998 25620
rect 14242 25564 14252 25620
rect 14308 25564 15148 25620
rect 29586 25564 29596 25620
rect 29652 25564 32060 25620
rect 32116 25564 32126 25620
rect 39890 25564 39900 25620
rect 39956 25564 42000 25620
rect 0 25536 800 25564
rect 15092 25508 15148 25564
rect 41200 25536 42000 25564
rect 15092 25452 16044 25508
rect 16100 25452 16110 25508
rect 18834 25452 18844 25508
rect 18900 25452 19628 25508
rect 19684 25452 21644 25508
rect 21700 25452 21710 25508
rect 27010 25452 27020 25508
rect 27076 25452 27804 25508
rect 27860 25452 37660 25508
rect 37716 25452 37726 25508
rect 12786 25340 12796 25396
rect 12852 25340 15932 25396
rect 15988 25340 15998 25396
rect 28242 25340 28252 25396
rect 28308 25340 29540 25396
rect 29484 25284 29540 25340
rect 4274 25228 4284 25284
rect 4340 25228 11564 25284
rect 11620 25228 14364 25284
rect 14420 25228 14430 25284
rect 15092 25228 15820 25284
rect 15876 25228 18060 25284
rect 18116 25228 19180 25284
rect 19236 25228 19246 25284
rect 20850 25228 20860 25284
rect 20916 25228 21420 25284
rect 21476 25228 21486 25284
rect 24994 25228 25004 25284
rect 25060 25228 25564 25284
rect 25620 25228 26012 25284
rect 26068 25228 28364 25284
rect 28420 25228 29148 25284
rect 29204 25228 29214 25284
rect 29484 25228 37884 25284
rect 37940 25228 37950 25284
rect 15092 25172 15148 25228
rect 14466 25116 14476 25172
rect 14532 25116 15148 25172
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 0 24948 800 24976
rect 41200 24948 42000 24976
rect 0 24892 2044 24948
rect 2100 24892 2110 24948
rect 22866 24892 22876 24948
rect 22932 24892 23436 24948
rect 23492 24892 26908 24948
rect 26964 24892 26974 24948
rect 40002 24892 40012 24948
rect 40068 24892 42000 24948
rect 0 24864 800 24892
rect 41200 24864 42000 24892
rect 13682 24780 13692 24836
rect 13748 24780 14924 24836
rect 14980 24780 14990 24836
rect 15586 24780 15596 24836
rect 15652 24780 25452 24836
rect 25508 24780 25518 24836
rect 26338 24780 26348 24836
rect 26404 24780 27580 24836
rect 27636 24780 27646 24836
rect 25890 24668 25900 24724
rect 25956 24668 26236 24724
rect 26292 24668 26302 24724
rect 26898 24668 26908 24724
rect 26964 24668 28140 24724
rect 28196 24668 28206 24724
rect 28466 24668 28476 24724
rect 28532 24668 29260 24724
rect 29316 24668 29820 24724
rect 29876 24668 29886 24724
rect 16706 24556 16716 24612
rect 16772 24556 17388 24612
rect 17444 24556 17454 24612
rect 25778 24556 25788 24612
rect 25844 24556 27244 24612
rect 27300 24556 27310 24612
rect 27682 24556 27692 24612
rect 27748 24556 28700 24612
rect 28756 24556 28766 24612
rect 25666 24444 25676 24500
rect 25732 24444 26236 24500
rect 26292 24444 26302 24500
rect 27794 24444 27804 24500
rect 27860 24444 28924 24500
rect 28980 24444 28990 24500
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 12114 23996 12124 24052
rect 12180 23996 13580 24052
rect 13636 23996 13646 24052
rect 4274 23884 4284 23940
rect 4340 23884 8428 23940
rect 12898 23884 12908 23940
rect 12964 23884 14364 23940
rect 14420 23884 14700 23940
rect 14756 23884 14766 23940
rect 26852 23884 27804 23940
rect 27860 23884 27870 23940
rect 8372 23716 8428 23884
rect 26852 23828 26908 23884
rect 13794 23772 13804 23828
rect 13860 23772 15036 23828
rect 15092 23772 15102 23828
rect 26338 23772 26348 23828
rect 26404 23772 26908 23828
rect 8372 23660 9996 23716
rect 10052 23660 14028 23716
rect 14084 23660 14094 23716
rect 0 23604 800 23632
rect 0 23548 1932 23604
rect 1988 23548 1998 23604
rect 0 23520 800 23548
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 13570 23324 13580 23380
rect 13636 23324 14364 23380
rect 14420 23324 14430 23380
rect 20738 23324 20748 23380
rect 20804 23324 20972 23380
rect 21028 23324 21038 23380
rect 14690 23100 14700 23156
rect 14756 23100 15708 23156
rect 15764 23100 15774 23156
rect 21298 22876 21308 22932
rect 21364 22876 21756 22932
rect 21812 22876 21822 22932
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 14242 22428 14252 22484
rect 14308 22428 16156 22484
rect 16212 22428 16222 22484
rect 22754 22428 22764 22484
rect 22820 22428 26012 22484
rect 26068 22428 26796 22484
rect 26852 22428 26862 22484
rect 30146 22428 30156 22484
rect 30212 22428 32060 22484
rect 32116 22428 37660 22484
rect 37716 22428 37726 22484
rect 14466 22316 14476 22372
rect 14532 22316 14924 22372
rect 14980 22316 17388 22372
rect 17444 22316 26124 22372
rect 26180 22316 26190 22372
rect 26450 22316 26460 22372
rect 26516 22316 27692 22372
rect 27748 22316 28252 22372
rect 28308 22316 28318 22372
rect 25564 22260 25620 22316
rect 41200 22260 42000 22288
rect 15922 22204 15932 22260
rect 15988 22204 16940 22260
rect 16996 22204 17006 22260
rect 25554 22204 25564 22260
rect 25620 22204 25630 22260
rect 28130 22204 28140 22260
rect 28196 22204 29932 22260
rect 29988 22204 29998 22260
rect 40002 22204 40012 22260
rect 40068 22204 42000 22260
rect 41200 22176 42000 22204
rect 13234 22092 13244 22148
rect 13300 22092 16380 22148
rect 16436 22092 16828 22148
rect 16884 22092 16894 22148
rect 17714 22092 17724 22148
rect 17780 22092 19292 22148
rect 19348 22092 19358 22148
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 23202 21868 23212 21924
rect 23268 21868 28028 21924
rect 28084 21868 28094 21924
rect 14690 21756 14700 21812
rect 14756 21756 15148 21812
rect 15204 21756 15214 21812
rect 15698 21756 15708 21812
rect 15764 21756 16268 21812
rect 16324 21756 19404 21812
rect 19460 21756 19470 21812
rect 22306 21756 22316 21812
rect 22372 21756 25452 21812
rect 25508 21756 31948 21812
rect 21970 21644 21980 21700
rect 22036 21644 23548 21700
rect 23604 21644 23614 21700
rect 25778 21644 25788 21700
rect 25844 21644 26348 21700
rect 26404 21644 27132 21700
rect 27188 21644 27198 21700
rect 31892 21588 31948 21756
rect 41200 21588 42000 21616
rect 13906 21532 13916 21588
rect 13972 21532 17668 21588
rect 18386 21532 18396 21588
rect 18452 21532 22876 21588
rect 22932 21532 25452 21588
rect 25508 21532 25518 21588
rect 17612 21476 17668 21532
rect 25452 21476 25508 21532
rect 11106 21420 11116 21476
rect 11172 21420 15708 21476
rect 15764 21420 15774 21476
rect 17602 21420 17612 21476
rect 17668 21420 17678 21476
rect 23314 21420 23324 21476
rect 23380 21420 24220 21476
rect 24276 21420 24286 21476
rect 25452 21420 25788 21476
rect 25844 21420 26124 21476
rect 26180 21420 26190 21476
rect 26852 21364 26908 21588
rect 26964 21532 26974 21588
rect 31892 21532 37660 21588
rect 37716 21532 37726 21588
rect 40002 21532 40012 21588
rect 40068 21532 42000 21588
rect 41200 21504 42000 21532
rect 14914 21308 14924 21364
rect 14980 21308 18620 21364
rect 18676 21308 18686 21364
rect 25554 21308 25564 21364
rect 25620 21308 26460 21364
rect 26516 21308 26908 21364
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 14690 20972 14700 21028
rect 14756 20972 16268 21028
rect 16324 20972 16334 21028
rect 27570 20972 27580 21028
rect 27636 20972 29036 21028
rect 29092 20972 29102 21028
rect 41200 20916 42000 20944
rect 18274 20860 18284 20916
rect 18340 20860 21196 20916
rect 21252 20860 22092 20916
rect 22148 20860 22158 20916
rect 40002 20860 40012 20916
rect 40068 20860 42000 20916
rect 41200 20832 42000 20860
rect 16594 20748 16604 20804
rect 16660 20748 17276 20804
rect 17332 20748 17342 20804
rect 18162 20748 18172 20804
rect 18228 20748 18732 20804
rect 18788 20748 20412 20804
rect 20468 20748 20478 20804
rect 22642 20748 22652 20804
rect 22708 20748 23324 20804
rect 23380 20748 23390 20804
rect 31892 20748 37660 20804
rect 37716 20748 37726 20804
rect 16482 20636 16492 20692
rect 16548 20636 17164 20692
rect 17220 20636 17230 20692
rect 21970 20636 21980 20692
rect 22036 20636 23436 20692
rect 23492 20636 23502 20692
rect 31892 20580 31948 20748
rect 13458 20524 13468 20580
rect 13524 20524 13916 20580
rect 13972 20524 14252 20580
rect 14308 20524 14318 20580
rect 15922 20524 15932 20580
rect 15988 20524 18060 20580
rect 18116 20524 18126 20580
rect 20066 20524 20076 20580
rect 20132 20524 22204 20580
rect 22260 20524 22988 20580
rect 23044 20524 23884 20580
rect 23940 20524 25340 20580
rect 25396 20524 25406 20580
rect 29250 20524 29260 20580
rect 29316 20524 29708 20580
rect 29764 20524 31948 20580
rect 18946 20412 18956 20468
rect 19012 20412 19404 20468
rect 19460 20412 19470 20468
rect 21410 20412 21420 20468
rect 21476 20412 22876 20468
rect 22932 20412 22942 20468
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 25442 20188 25452 20244
rect 25508 20188 26796 20244
rect 26852 20188 26862 20244
rect 8372 20076 9996 20132
rect 10052 20076 13692 20132
rect 13748 20076 13758 20132
rect 16370 20076 16380 20132
rect 16436 20076 17724 20132
rect 17780 20076 17790 20132
rect 18946 20076 18956 20132
rect 19012 20076 21420 20132
rect 21476 20076 21486 20132
rect 30146 20076 30156 20132
rect 30212 20076 31948 20132
rect 8372 20020 8428 20076
rect 31892 20020 31948 20076
rect 4274 19964 4284 20020
rect 4340 19964 8428 20020
rect 17378 19964 17388 20020
rect 17444 19964 18844 20020
rect 18900 19964 18910 20020
rect 26898 19964 26908 20020
rect 26964 19964 28812 20020
rect 28868 19964 28878 20020
rect 31892 19964 32060 20020
rect 32116 19964 37660 20020
rect 37716 19964 37726 20020
rect 20066 19852 20076 19908
rect 20132 19852 20636 19908
rect 20692 19852 23660 19908
rect 23716 19852 25228 19908
rect 25284 19852 25294 19908
rect 29250 19852 29260 19908
rect 29316 19852 30716 19908
rect 30772 19852 30782 19908
rect 1922 19740 1932 19796
rect 1988 19740 1998 19796
rect 19394 19740 19404 19796
rect 19460 19740 20524 19796
rect 20580 19740 20590 19796
rect 28690 19740 28700 19796
rect 28756 19740 30156 19796
rect 30212 19740 30222 19796
rect 0 19572 800 19600
rect 1932 19572 1988 19740
rect 18274 19628 18284 19684
rect 18340 19628 20300 19684
rect 20356 19628 21308 19684
rect 21364 19628 21374 19684
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 41200 19572 42000 19600
rect 0 19516 1988 19572
rect 40002 19516 40012 19572
rect 40068 19516 42000 19572
rect 0 19488 800 19516
rect 41200 19488 42000 19516
rect 13346 19404 13356 19460
rect 13412 19404 13804 19460
rect 13860 19404 15260 19460
rect 15316 19404 15326 19460
rect 19394 19404 19404 19460
rect 19460 19404 23772 19460
rect 23828 19404 23838 19460
rect 16818 19292 16828 19348
rect 16884 19292 17724 19348
rect 17780 19292 18396 19348
rect 18452 19292 18462 19348
rect 13794 19180 13804 19236
rect 13860 19180 15148 19236
rect 15362 19180 15372 19236
rect 15428 19180 16604 19236
rect 16660 19180 20524 19236
rect 20580 19180 20590 19236
rect 26898 19180 26908 19236
rect 26964 19180 28028 19236
rect 28084 19180 28094 19236
rect 15092 19124 15148 19180
rect 12114 19068 12124 19124
rect 12180 19068 13580 19124
rect 13636 19068 13646 19124
rect 15092 19068 17052 19124
rect 17108 19068 18956 19124
rect 19012 19068 19022 19124
rect 19618 19068 19628 19124
rect 19684 19068 19964 19124
rect 20020 19068 20030 19124
rect 24434 19068 24444 19124
rect 24500 19068 26348 19124
rect 26404 19068 26414 19124
rect 28130 19068 28140 19124
rect 28196 19068 29932 19124
rect 29988 19068 29998 19124
rect 4162 18956 4172 19012
rect 4228 18956 19740 19012
rect 19796 18956 19806 19012
rect 21858 18956 21868 19012
rect 21924 18956 22764 19012
rect 22820 18956 24780 19012
rect 24836 18956 24846 19012
rect 25554 18956 25564 19012
rect 25620 18956 28252 19012
rect 28308 18956 28318 19012
rect 17266 18844 17276 18900
rect 17332 18844 18284 18900
rect 18340 18844 18350 18900
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 20412 18732 28028 18788
rect 28084 18732 28094 18788
rect 20412 18676 20468 18732
rect 16594 18620 16604 18676
rect 16660 18620 17948 18676
rect 18004 18620 20468 18676
rect 20626 18620 20636 18676
rect 20692 18620 21532 18676
rect 21588 18620 21598 18676
rect 21858 18620 21868 18676
rect 21924 18620 22428 18676
rect 22484 18620 23436 18676
rect 23492 18620 23884 18676
rect 23940 18620 23950 18676
rect 24210 18620 24220 18676
rect 24276 18620 25564 18676
rect 25620 18620 25630 18676
rect 21532 18564 21588 18620
rect 12114 18508 12124 18564
rect 12180 18508 13468 18564
rect 13524 18508 13534 18564
rect 21532 18508 22316 18564
rect 22372 18508 22382 18564
rect 22866 18508 22876 18564
rect 22932 18508 23996 18564
rect 24052 18508 24062 18564
rect 26226 18508 26236 18564
rect 26292 18508 27356 18564
rect 27412 18508 27422 18564
rect 4274 18396 4284 18452
rect 4340 18396 8428 18452
rect 14130 18396 14140 18452
rect 14196 18396 15036 18452
rect 15092 18396 15102 18452
rect 20850 18396 20860 18452
rect 20916 18396 22540 18452
rect 22596 18396 22606 18452
rect 22978 18396 22988 18452
rect 23044 18396 23660 18452
rect 23716 18396 23726 18452
rect 25218 18396 25228 18452
rect 25284 18396 26012 18452
rect 26068 18396 26078 18452
rect 8372 18340 8428 18396
rect 8372 18284 9996 18340
rect 10052 18284 14588 18340
rect 14644 18284 14654 18340
rect 21970 18284 21980 18340
rect 22036 18284 23212 18340
rect 23268 18284 23278 18340
rect 0 18228 800 18256
rect 0 18172 1932 18228
rect 1988 18172 1998 18228
rect 16370 18172 16380 18228
rect 16436 18172 17388 18228
rect 17444 18172 17454 18228
rect 18610 18172 18620 18228
rect 18676 18172 21756 18228
rect 21812 18172 23548 18228
rect 23604 18172 27580 18228
rect 27636 18172 27646 18228
rect 0 18144 800 18172
rect 15138 18060 15148 18116
rect 15204 18060 20748 18116
rect 20804 18060 25452 18116
rect 25508 18060 25518 18116
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 20402 17836 20412 17892
rect 20468 17836 25228 17892
rect 25284 17836 25294 17892
rect 19282 17724 19292 17780
rect 19348 17724 22204 17780
rect 22260 17724 26460 17780
rect 26516 17724 26526 17780
rect 12898 17612 12908 17668
rect 12964 17612 13580 17668
rect 13636 17612 13646 17668
rect 15250 17612 15260 17668
rect 15316 17612 15708 17668
rect 15764 17612 15774 17668
rect 26338 17612 26348 17668
rect 26404 17612 26908 17668
rect 28354 17612 28364 17668
rect 28420 17612 29932 17668
rect 29988 17612 37660 17668
rect 37716 17612 37726 17668
rect 15708 17444 15764 17612
rect 26852 17556 26908 17612
rect 41200 17556 42000 17584
rect 26852 17500 27916 17556
rect 27972 17500 27982 17556
rect 40002 17500 40012 17556
rect 40068 17500 42000 17556
rect 41200 17472 42000 17500
rect 15708 17388 17724 17444
rect 17780 17388 17790 17444
rect 25218 17388 25228 17444
rect 25284 17388 26012 17444
rect 26068 17388 27804 17444
rect 27860 17388 27870 17444
rect 26898 17276 26908 17332
rect 26964 17276 27692 17332
rect 27748 17276 27758 17332
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 21746 17052 21756 17108
rect 21812 17052 23772 17108
rect 23828 17052 24892 17108
rect 24948 17052 24958 17108
rect 27346 17052 27356 17108
rect 27412 17052 27692 17108
rect 27748 17052 27758 17108
rect 14466 16940 14476 16996
rect 14532 16940 15484 16996
rect 15540 16940 15550 16996
rect 27122 16940 27132 16996
rect 27188 16940 27580 16996
rect 27636 16940 27646 16996
rect 41200 16884 42000 16912
rect 13794 16828 13804 16884
rect 13860 16828 17500 16884
rect 17556 16828 17566 16884
rect 27010 16828 27020 16884
rect 27076 16828 28140 16884
rect 28196 16828 28206 16884
rect 40002 16828 40012 16884
rect 40068 16828 42000 16884
rect 41200 16800 42000 16828
rect 23874 16716 23884 16772
rect 23940 16716 24556 16772
rect 24612 16716 24622 16772
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 18386 16044 18396 16100
rect 18452 16044 18956 16100
rect 19012 16044 19852 16100
rect 19908 16044 19918 16100
rect 20066 16044 20076 16100
rect 20132 16044 23884 16100
rect 23940 16044 23950 16100
rect 27682 16044 27692 16100
rect 27748 16044 30828 16100
rect 30884 16044 30894 16100
rect 20076 15988 20132 16044
rect 18498 15932 18508 15988
rect 18564 15932 20132 15988
rect 26562 15932 26572 15988
rect 26628 15932 27244 15988
rect 27300 15932 27310 15988
rect 19058 15820 19068 15876
rect 19124 15820 19964 15876
rect 20020 15820 20030 15876
rect 25218 15820 25228 15876
rect 25284 15820 25788 15876
rect 25844 15820 25854 15876
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 24210 15372 24220 15428
rect 24276 15372 25116 15428
rect 25172 15372 26236 15428
rect 26292 15372 26302 15428
rect 21634 15260 21644 15316
rect 21700 15260 22988 15316
rect 23044 15260 25340 15316
rect 25396 15260 25406 15316
rect 26908 15204 26964 15932
rect 25218 15148 25228 15204
rect 25284 15148 26908 15204
rect 26964 15148 26974 15204
rect 30818 15148 30828 15204
rect 30884 15148 37660 15204
rect 37716 15148 37726 15204
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 17490 14588 17500 14644
rect 17556 14588 18396 14644
rect 18452 14588 20860 14644
rect 20916 14588 21420 14644
rect 21476 14588 21486 14644
rect 25666 14588 25676 14644
rect 25732 14588 29260 14644
rect 29316 14588 29326 14644
rect 31892 14476 37660 14532
rect 37716 14476 37726 14532
rect 31892 14420 31948 14476
rect 27458 14364 27468 14420
rect 27524 14364 28588 14420
rect 28644 14364 31948 14420
rect 41200 14196 42000 14224
rect 40002 14140 40012 14196
rect 40068 14140 42000 14196
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 41200 14112 42000 14140
rect 26786 13804 26796 13860
rect 26852 13804 28700 13860
rect 28756 13804 28766 13860
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 25666 13020 25676 13076
rect 25732 13020 26460 13076
rect 26516 13020 26526 13076
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 27122 4060 27132 4116
rect 27188 4060 29708 4116
rect 29764 4060 29774 4116
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 21522 3612 21532 3668
rect 21588 3612 22428 3668
rect 22484 3612 22494 3668
rect 24210 3612 24220 3668
rect 24276 3612 25564 3668
rect 25620 3612 25630 3668
rect 26226 3612 26236 3668
rect 26292 3612 29372 3668
rect 29428 3612 29438 3668
rect 26114 3500 26124 3556
rect 26180 3500 28588 3556
rect 28644 3500 28654 3556
rect 25554 3388 25564 3444
rect 25620 3388 26796 3444
rect 26852 3388 26862 3444
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
<< via3 >>
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
<< metal4 >>
rect 4448 38444 4768 38476
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 37660 20128 38476
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19808 34524 20128 36036
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 19808 23548 20128 25060
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 19808 21980 20128 23492
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 38444 35488 38476
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _115_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21168 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _116_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 22736 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _117_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21056 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _118_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21616 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _119_
timestamp 1698175906
transform -1 0 23072 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _120_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19264 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _121_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 15456 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _122_
timestamp 1698175906
transform -1 0 20944 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _123_
timestamp 1698175906
transform -1 0 20944 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _124_
timestamp 1698175906
transform 1 0 16800 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _125_
timestamp 1698175906
transform 1 0 21168 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _126_
timestamp 1698175906
transform 1 0 23296 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _127_
timestamp 1698175906
transform -1 0 19600 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _128_
timestamp 1698175906
transform -1 0 20384 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _129_
timestamp 1698175906
transform -1 0 17920 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _130_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19376 0 1 20384
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _131_
timestamp 1698175906
transform -1 0 16016 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _132_
timestamp 1698175906
transform 1 0 18592 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _133_
timestamp 1698175906
transform 1 0 17248 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _134_
timestamp 1698175906
transform -1 0 16688 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _135_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 13888 0 -1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _136_
timestamp 1698175906
transform 1 0 21280 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _137_
timestamp 1698175906
transform 1 0 21504 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _138_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 23296 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _139_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 19376 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _140_
timestamp 1698175906
transform -1 0 14000 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _141_
timestamp 1698175906
transform 1 0 14112 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _142_
timestamp 1698175906
transform 1 0 16352 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _143_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 17024 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _144_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 14448 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _145_
timestamp 1698175906
transform 1 0 14672 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _146_
timestamp 1698175906
transform -1 0 16240 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _147_
timestamp 1698175906
transform 1 0 15344 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _148_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 15344 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _149_
timestamp 1698175906
transform -1 0 15680 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _150_
timestamp 1698175906
transform 1 0 23744 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _151_
timestamp 1698175906
transform 1 0 15904 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _152_
timestamp 1698175906
transform 1 0 22400 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _153_
timestamp 1698175906
transform 1 0 28000 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _154_
timestamp 1698175906
transform 1 0 29904 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _155_
timestamp 1698175906
transform 1 0 27888 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _156_
timestamp 1698175906
transform -1 0 17136 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _157_
timestamp 1698175906
transform -1 0 18480 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _158_
timestamp 1698175906
transform -1 0 18144 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _159_
timestamp 1698175906
transform -1 0 16576 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _160_
timestamp 1698175906
transform 1 0 23744 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _161_
timestamp 1698175906
transform 1 0 17360 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _162_
timestamp 1698175906
transform -1 0 18368 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _163_
timestamp 1698175906
transform -1 0 19040 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _164_
timestamp 1698175906
transform 1 0 19824 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _165_
timestamp 1698175906
transform -1 0 19936 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _166_
timestamp 1698175906
transform 1 0 25088 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _167_
timestamp 1698175906
transform -1 0 25872 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _168_
timestamp 1698175906
transform -1 0 21840 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _169_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19712 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _170_
timestamp 1698175906
transform -1 0 18928 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _171_
timestamp 1698175906
transform 1 0 16240 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _172_
timestamp 1698175906
transform 1 0 17248 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _173_
timestamp 1698175906
transform -1 0 17920 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _174_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 17808 0 1 20384
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _175_
timestamp 1698175906
transform -1 0 16912 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _176_
timestamp 1698175906
transform -1 0 15568 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _177_
timestamp 1698175906
transform -1 0 14000 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _178_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 15344 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _179_
timestamp 1698175906
transform 1 0 13328 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _180_
timestamp 1698175906
transform -1 0 14784 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _181_
timestamp 1698175906
transform -1 0 15904 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _182_
timestamp 1698175906
transform 1 0 13216 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _183_
timestamp 1698175906
transform 1 0 18144 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _184_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21392 0 -1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _185_
timestamp 1698175906
transform 1 0 17920 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _186_
timestamp 1698175906
transform 1 0 22848 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _187_
timestamp 1698175906
transform 1 0 17808 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _188_
timestamp 1698175906
transform 1 0 21728 0 1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _189_
timestamp 1698175906
transform 1 0 22848 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _190_
timestamp 1698175906
transform 1 0 18816 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _191_
timestamp 1698175906
transform 1 0 23968 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _192_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 23408 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _193_
timestamp 1698175906
transform 1 0 21168 0 1 18816
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _194_
timestamp 1698175906
transform 1 0 20384 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _195_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 22400 0 -1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _196_
timestamp 1698175906
transform 1 0 22064 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _197_
timestamp 1698175906
transform -1 0 22960 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _198_
timestamp 1698175906
transform -1 0 26320 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _199_
timestamp 1698175906
transform 1 0 24752 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _200_
timestamp 1698175906
transform 1 0 27440 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _201_
timestamp 1698175906
transform 1 0 26320 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _202_
timestamp 1698175906
transform 1 0 26768 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _203_
timestamp 1698175906
transform 1 0 25312 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _204_
timestamp 1698175906
transform -1 0 26544 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _205_
timestamp 1698175906
transform 1 0 27216 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _206_
timestamp 1698175906
transform -1 0 22848 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _207_
timestamp 1698175906
transform -1 0 21952 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _208_
timestamp 1698175906
transform -1 0 27776 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _209_
timestamp 1698175906
transform 1 0 24640 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _210_
timestamp 1698175906
transform 1 0 26096 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _211_
timestamp 1698175906
transform -1 0 27440 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _212_
timestamp 1698175906
transform -1 0 25536 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _213_
timestamp 1698175906
transform -1 0 24640 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _214_
timestamp 1698175906
transform 1 0 25984 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _215_
timestamp 1698175906
transform -1 0 30240 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _216_
timestamp 1698175906
transform 1 0 27888 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _217_
timestamp 1698175906
transform -1 0 26544 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _218_
timestamp 1698175906
transform 1 0 28560 0 -1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _219_
timestamp 1698175906
transform 1 0 28784 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _220_
timestamp 1698175906
transform 1 0 28000 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _221_
timestamp 1698175906
transform 1 0 25648 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _222_
timestamp 1698175906
transform -1 0 26096 0 -1 25088
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _223_
timestamp 1698175906
transform 1 0 27104 0 -1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _224_
timestamp 1698175906
transform 1 0 26096 0 -1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _225_
timestamp 1698175906
transform 1 0 26208 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _226_
timestamp 1698175906
transform -1 0 23632 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _227_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 22400 0 1 25088
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _228_
timestamp 1698175906
transform -1 0 29568 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _229_
timestamp 1698175906
transform 1 0 26768 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _230_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17248 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _231_
timestamp 1698175906
transform -1 0 13104 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _232_
timestamp 1698175906
transform -1 0 14672 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _233_
timestamp 1698175906
transform -1 0 15904 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _234_
timestamp 1698175906
transform 1 0 29008 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _235_
timestamp 1698175906
transform -1 0 14224 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _236_
timestamp 1698175906
transform 1 0 13552 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _237_
timestamp 1698175906
transform 1 0 17248 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _238_
timestamp 1698175906
transform 1 0 17920 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _239_
timestamp 1698175906
transform 1 0 18144 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _240_
timestamp 1698175906
transform 1 0 15792 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _241_
timestamp 1698175906
transform -1 0 13104 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _242_
timestamp 1698175906
transform -1 0 13104 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _243_
timestamp 1698175906
transform 1 0 22512 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _244_
timestamp 1698175906
transform 1 0 21392 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _245_
timestamp 1698175906
transform 1 0 26880 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _246_
timestamp 1698175906
transform 1 0 27776 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _247_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21056 0 -1 28224
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _248_
timestamp 1698175906
transform 1 0 25536 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _249_
timestamp 1698175906
transform 1 0 22848 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _250_
timestamp 1698175906
transform 1 0 29008 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _251_
timestamp 1698175906
transform 1 0 29008 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _252_
timestamp 1698175906
transform 1 0 25424 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _253_
timestamp 1698175906
transform 1 0 24752 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _254_
timestamp 1698175906
transform 1 0 20272 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _255_
timestamp 1698175906
transform 1 0 26656 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _256_
timestamp 1698175906
transform 1 0 23184 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _257_
timestamp 1698175906
transform 1 0 26320 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _258_
timestamp 1698175906
transform 1 0 25648 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _259_
timestamp 1698175906
transform 1 0 23184 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__182__C dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 15008 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__204__B
timestamp 1698175906
transform 1 0 25424 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__227__A3
timestamp 1698175906
transform 1 0 20720 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__230__CLK
timestamp 1698175906
transform -1 0 20944 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__231__CLK
timestamp 1698175906
transform 1 0 13104 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__232__CLK
timestamp 1698175906
transform 1 0 14672 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__233__CLK
timestamp 1698175906
transform 1 0 16128 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__234__CLK
timestamp 1698175906
transform 1 0 28784 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__235__CLK
timestamp 1698175906
transform 1 0 14224 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__236__CLK
timestamp 1698175906
transform 1 0 17472 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__237__CLK
timestamp 1698175906
transform -1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__238__CLK
timestamp 1698175906
transform 1 0 21392 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__239__CLK
timestamp 1698175906
transform 1 0 21392 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__240__CLK
timestamp 1698175906
transform 1 0 19152 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__241__CLK
timestamp 1698175906
transform 1 0 13104 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__242__CLK
timestamp 1698175906
transform 1 0 13552 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__243__CLK
timestamp 1698175906
transform 1 0 25984 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__244__CLK
timestamp 1698175906
transform 1 0 25312 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__245__CLK
timestamp 1698175906
transform 1 0 26656 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__246__CLK
timestamp 1698175906
transform 1 0 28112 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__247__CLK
timestamp 1698175906
transform -1 0 25536 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__248__CLK
timestamp 1698175906
transform 1 0 29232 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__249__CLK
timestamp 1698175906
transform -1 0 26544 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__250__CLK
timestamp 1698175906
transform 1 0 28784 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__251__CLK
timestamp 1698175906
transform 1 0 29456 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__252__CLK
timestamp 1698175906
transform 1 0 29904 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__253__CLK
timestamp 1698175906
transform 1 0 28336 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__254__CLK
timestamp 1698175906
transform 1 0 20048 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__255__CLK
timestamp 1698175906
transform 1 0 30688 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1698175906
transform -1 0 19824 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19264 0 -1 20384
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1698175906
transform -1 0 22848 0 -1 21952
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1698175906
transform 1 0 23184 0 1 20384
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1568 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698175906
transform 1 0 5376 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698175906
transform 1 0 9184 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698175906
transform 1 0 12992 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_138
timestamp 1698175906
transform 1 0 16800 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_172 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 20608 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_176 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21056 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_232
timestamp 1698175906
transform 1 0 27328 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_236
timestamp 1698175906
transform 1 0 27776 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_266
timestamp 1698175906
transform 1 0 31136 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_270
timestamp 1698175906
transform 1 0 31584 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_274
timestamp 1698175906
transform 1 0 32032 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_308
timestamp 1698175906
transform 1 0 35840 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_342
timestamp 1698175906
transform 1 0 39648 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_346
timestamp 1698175906
transform 1 0 40096 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_348 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 40320 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1568 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698175906
transform 1 0 8736 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698175906
transform 1 0 9408 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698175906
transform 1 0 16576 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_142
timestamp 1698175906
transform 1 0 17248 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_206
timestamp 1698175906
transform 1 0 24416 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_212
timestamp 1698175906
transform 1 0 25088 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_216
timestamp 1698175906
transform 1 0 25536 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_269 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 31472 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_277
timestamp 1698175906
transform 1 0 32368 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_279
timestamp 1698175906
transform 1 0 32592 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_282
timestamp 1698175906
transform 1 0 32928 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_346
timestamp 1698175906
transform 1 0 40096 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_348
timestamp 1698175906
transform 1 0 40320 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698175906
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698175906
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698175906
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698175906
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_107
timestamp 1698175906
transform 1 0 13328 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_171
timestamp 1698175906
transform 1 0 20496 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_177
timestamp 1698175906
transform 1 0 21168 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_241
timestamp 1698175906
transform 1 0 28336 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698175906
transform 1 0 29008 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698175906
transform 1 0 36176 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_317
timestamp 1698175906
transform 1 0 36848 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698175906
transform 1 0 1568 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698175906
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698175906
transform 1 0 9408 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698175906
transform 1 0 16576 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_142
timestamp 1698175906
transform 1 0 17248 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_206
timestamp 1698175906
transform 1 0 24416 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_212
timestamp 1698175906
transform 1 0 25088 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_276
timestamp 1698175906
transform 1 0 32256 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_282
timestamp 1698175906
transform 1 0 32928 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_346
timestamp 1698175906
transform 1 0 40096 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_348
timestamp 1698175906
transform 1 0 40320 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698175906
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698175906
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698175906
transform 1 0 5488 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698175906
transform 1 0 12656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_107
timestamp 1698175906
transform 1 0 13328 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698175906
transform 1 0 20496 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_177
timestamp 1698175906
transform 1 0 21168 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_241
timestamp 1698175906
transform 1 0 28336 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698175906
transform 1 0 29008 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698175906
transform 1 0 36176 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_317
timestamp 1698175906
transform 1 0 36848 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698175906
transform 1 0 1568 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698175906
transform 1 0 8736 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698175906
transform 1 0 9408 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698175906
transform 1 0 16576 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_142
timestamp 1698175906
transform 1 0 17248 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_206
timestamp 1698175906
transform 1 0 24416 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_212
timestamp 1698175906
transform 1 0 25088 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698175906
transform 1 0 32256 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_282
timestamp 1698175906
transform 1 0 32928 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_346
timestamp 1698175906
transform 1 0 40096 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_348
timestamp 1698175906
transform 1 0 40320 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698175906
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698175906
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698175906
transform 1 0 5488 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698175906
transform 1 0 12656 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_107
timestamp 1698175906
transform 1 0 13328 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_171
timestamp 1698175906
transform 1 0 20496 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_177
timestamp 1698175906
transform 1 0 21168 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_241
timestamp 1698175906
transform 1 0 28336 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_247
timestamp 1698175906
transform 1 0 29008 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_311
timestamp 1698175906
transform 1 0 36176 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_317
timestamp 1698175906
transform 1 0 36848 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698175906
transform 1 0 1568 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698175906
transform 1 0 8736 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_72
timestamp 1698175906
transform 1 0 9408 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698175906
transform 1 0 16576 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_142
timestamp 1698175906
transform 1 0 17248 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_206
timestamp 1698175906
transform 1 0 24416 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_212
timestamp 1698175906
transform 1 0 25088 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_276
timestamp 1698175906
transform 1 0 32256 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_282
timestamp 1698175906
transform 1 0 32928 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_346
timestamp 1698175906
transform 1 0 40096 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_348
timestamp 1698175906
transform 1 0 40320 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698175906
transform 1 0 1568 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698175906
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_37
timestamp 1698175906
transform 1 0 5488 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_101
timestamp 1698175906
transform 1 0 12656 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_107
timestamp 1698175906
transform 1 0 13328 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_171
timestamp 1698175906
transform 1 0 20496 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_177
timestamp 1698175906
transform 1 0 21168 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_241
timestamp 1698175906
transform 1 0 28336 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_247
timestamp 1698175906
transform 1 0 29008 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_311
timestamp 1698175906
transform 1 0 36176 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_317
timestamp 1698175906
transform 1 0 36848 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698175906
transform 1 0 1568 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698175906
transform 1 0 8736 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_72
timestamp 1698175906
transform 1 0 9408 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_136
timestamp 1698175906
transform 1 0 16576 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_142
timestamp 1698175906
transform 1 0 17248 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_206
timestamp 1698175906
transform 1 0 24416 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_212
timestamp 1698175906
transform 1 0 25088 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_276
timestamp 1698175906
transform 1 0 32256 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_282
timestamp 1698175906
transform 1 0 32928 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_346
timestamp 1698175906
transform 1 0 40096 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_348
timestamp 1698175906
transform 1 0 40320 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698175906
transform 1 0 1568 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698175906
transform 1 0 5152 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_37
timestamp 1698175906
transform 1 0 5488 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698175906
transform 1 0 12656 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_107
timestamp 1698175906
transform 1 0 13328 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_171
timestamp 1698175906
transform 1 0 20496 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_177
timestamp 1698175906
transform 1 0 21168 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_241
timestamp 1698175906
transform 1 0 28336 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_247
timestamp 1698175906
transform 1 0 29008 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_311
timestamp 1698175906
transform 1 0 36176 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_317
timestamp 1698175906
transform 1 0 36848 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2
timestamp 1698175906
transform 1 0 1568 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698175906
transform 1 0 8736 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_72
timestamp 1698175906
transform 1 0 9408 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698175906
transform 1 0 16576 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_142
timestamp 1698175906
transform 1 0 17248 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_206
timestamp 1698175906
transform 1 0 24416 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_212
timestamp 1698175906
transform 1 0 25088 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_276
timestamp 1698175906
transform 1 0 32256 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_282
timestamp 1698175906
transform 1 0 32928 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_346
timestamp 1698175906
transform 1 0 40096 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_348
timestamp 1698175906
transform 1 0 40320 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698175906
transform 1 0 1568 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698175906
transform 1 0 5152 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_37
timestamp 1698175906
transform 1 0 5488 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698175906
transform 1 0 12656 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_107
timestamp 1698175906
transform 1 0 13328 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_171
timestamp 1698175906
transform 1 0 20496 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_177
timestamp 1698175906
transform 1 0 21168 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_185
timestamp 1698175906
transform 1 0 22064 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_189
timestamp 1698175906
transform 1 0 22512 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_191
timestamp 1698175906
transform 1 0 22736 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_221
timestamp 1698175906
transform 1 0 26096 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_225 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 26544 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_241
timestamp 1698175906
transform 1 0 28336 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_247
timestamp 1698175906
transform 1 0 29008 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_311
timestamp 1698175906
transform 1 0 36176 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_317
timestamp 1698175906
transform 1 0 36848 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_2
timestamp 1698175906
transform 1 0 1568 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_66
timestamp 1698175906
transform 1 0 8736 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_72
timestamp 1698175906
transform 1 0 9408 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_136
timestamp 1698175906
transform 1 0 16576 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_142
timestamp 1698175906
transform 1 0 17248 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_206
timestamp 1698175906
transform 1 0 24416 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_212
timestamp 1698175906
transform 1 0 25088 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_216
timestamp 1698175906
transform 1 0 25536 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_229
timestamp 1698175906
transform 1 0 26992 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_236
timestamp 1698175906
transform 1 0 27776 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_268
timestamp 1698175906
transform 1 0 31360 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_276
timestamp 1698175906
transform 1 0 32256 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_282
timestamp 1698175906
transform 1 0 32928 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_346
timestamp 1698175906
transform 1 0 40096 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_348
timestamp 1698175906
transform 1 0 40320 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698175906
transform 1 0 1568 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698175906
transform 1 0 5152 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_37
timestamp 1698175906
transform 1 0 5488 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_101
timestamp 1698175906
transform 1 0 12656 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_107
timestamp 1698175906
transform 1 0 13328 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_139
timestamp 1698175906
transform 1 0 16912 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_141
timestamp 1698175906
transform 1 0 17136 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_171
timestamp 1698175906
transform 1 0 20496 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_177
timestamp 1698175906
transform 1 0 21168 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_181
timestamp 1698175906
transform 1 0 21616 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_197
timestamp 1698175906
transform 1 0 23408 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_199
timestamp 1698175906
transform 1 0 23632 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_208
timestamp 1698175906
transform 1 0 24640 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_210
timestamp 1698175906
transform 1 0 24864 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_247
timestamp 1698175906
transform 1 0 29008 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_251
timestamp 1698175906
transform 1 0 29456 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_317
timestamp 1698175906
transform 1 0 36848 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_321
timestamp 1698175906
transform 1 0 37296 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_2
timestamp 1698175906
transform 1 0 1568 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_66
timestamp 1698175906
transform 1 0 8736 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_72
timestamp 1698175906
transform 1 0 9408 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_136
timestamp 1698175906
transform 1 0 16576 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_142
timestamp 1698175906
transform 1 0 17248 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_208
timestamp 1698175906
transform 1 0 24640 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_212
timestamp 1698175906
transform 1 0 25088 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_216
timestamp 1698175906
transform 1 0 25536 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_220
timestamp 1698175906
transform 1 0 25984 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_233
timestamp 1698175906
transform 1 0 27440 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_235
timestamp 1698175906
transform 1 0 27664 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_265
timestamp 1698175906
transform 1 0 31024 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_273
timestamp 1698175906
transform 1 0 31920 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_277
timestamp 1698175906
transform 1 0 32368 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_279
timestamp 1698175906
transform 1 0 32592 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_282
timestamp 1698175906
transform 1 0 32928 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_346
timestamp 1698175906
transform 1 0 40096 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_348
timestamp 1698175906
transform 1 0 40320 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_2
timestamp 1698175906
transform 1 0 1568 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698175906
transform 1 0 5152 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_37
timestamp 1698175906
transform 1 0 5488 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_101
timestamp 1698175906
transform 1 0 12656 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_107
timestamp 1698175906
transform 1 0 13328 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_139
timestamp 1698175906
transform 1 0 16912 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_147
timestamp 1698175906
transform 1 0 17808 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_149
timestamp 1698175906
transform 1 0 18032 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_158
timestamp 1698175906
transform 1 0 19040 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_162
timestamp 1698175906
transform 1 0 19488 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_174
timestamp 1698175906
transform 1 0 20832 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_183
timestamp 1698175906
transform 1 0 21840 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_193
timestamp 1698175906
transform 1 0 22960 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_225
timestamp 1698175906
transform 1 0 26544 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_237
timestamp 1698175906
transform 1 0 27888 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_241
timestamp 1698175906
transform 1 0 28336 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_247
timestamp 1698175906
transform 1 0 29008 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_311
timestamp 1698175906
transform 1 0 36176 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_317
timestamp 1698175906
transform 1 0 36848 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_2
timestamp 1698175906
transform 1 0 1568 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_66
timestamp 1698175906
transform 1 0 8736 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_72
timestamp 1698175906
transform 1 0 9408 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_104
timestamp 1698175906
transform 1 0 12992 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_108
timestamp 1698175906
transform 1 0 13440 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_138
timestamp 1698175906
transform 1 0 16800 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_142
timestamp 1698175906
transform 1 0 17248 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_152
timestamp 1698175906
transform 1 0 18368 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_168
timestamp 1698175906
transform 1 0 20160 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_176
timestamp 1698175906
transform 1 0 21056 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_184
timestamp 1698175906
transform 1 0 21952 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_200
timestamp 1698175906
transform 1 0 23744 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_208
timestamp 1698175906
transform 1 0 24640 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_212
timestamp 1698175906
transform 1 0 25088 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_220
timestamp 1698175906
transform 1 0 25984 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_224
timestamp 1698175906
transform 1 0 26432 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_257
timestamp 1698175906
transform 1 0 30128 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_273
timestamp 1698175906
transform 1 0 31920 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_277
timestamp 1698175906
transform 1 0 32368 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_279
timestamp 1698175906
transform 1 0 32592 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_282
timestamp 1698175906
transform 1 0 32928 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_314
timestamp 1698175906
transform 1 0 36512 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_322
timestamp 1698175906
transform 1 0 37408 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_2
timestamp 1698175906
transform 1 0 1568 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698175906
transform 1 0 5152 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_37
timestamp 1698175906
transform 1 0 5488 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_69
timestamp 1698175906
transform 1 0 9072 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_73
timestamp 1698175906
transform 1 0 9520 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_75
timestamp 1698175906
transform 1 0 9744 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_107
timestamp 1698175906
transform 1 0 13328 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_111
timestamp 1698175906
transform 1 0 13776 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_119
timestamp 1698175906
transform 1 0 14672 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_121
timestamp 1698175906
transform 1 0 14896 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_136
timestamp 1698175906
transform 1 0 16576 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_140
timestamp 1698175906
transform 1 0 17024 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_142
timestamp 1698175906
transform 1 0 17248 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_149
timestamp 1698175906
transform 1 0 18032 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_165
timestamp 1698175906
transform 1 0 19824 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_173
timestamp 1698175906
transform 1 0 20720 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_183
timestamp 1698175906
transform 1 0 21840 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_193
timestamp 1698175906
transform 1 0 22960 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_207
timestamp 1698175906
transform 1 0 24528 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_215
timestamp 1698175906
transform 1 0 25424 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_243
timestamp 1698175906
transform 1 0 28560 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_247
timestamp 1698175906
transform 1 0 29008 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_311
timestamp 1698175906
transform 1 0 36176 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_317
timestamp 1698175906
transform 1 0 36848 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_321
timestamp 1698175906
transform 1 0 37296 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_28
timestamp 1698175906
transform 1 0 4480 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_60
timestamp 1698175906
transform 1 0 8064 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_68
timestamp 1698175906
transform 1 0 8960 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_72
timestamp 1698175906
transform 1 0 9408 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_104
timestamp 1698175906
transform 1 0 12992 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_120
timestamp 1698175906
transform 1 0 14784 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_124
timestamp 1698175906
transform 1 0 15232 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_132
timestamp 1698175906
transform 1 0 16128 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_156
timestamp 1698175906
transform 1 0 18816 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_172
timestamp 1698175906
transform 1 0 20608 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_176
timestamp 1698175906
transform 1 0 21056 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_178
timestamp 1698175906
transform 1 0 21280 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_197
timestamp 1698175906
transform 1 0 23408 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_199
timestamp 1698175906
transform 1 0 23632 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_205
timestamp 1698175906
transform 1 0 24304 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_209
timestamp 1698175906
transform 1 0 24752 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_212
timestamp 1698175906
transform 1 0 25088 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_214
timestamp 1698175906
transform 1 0 25312 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_225
timestamp 1698175906
transform 1 0 26544 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_229
timestamp 1698175906
transform 1 0 26992 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_236
timestamp 1698175906
transform 1 0 27776 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_244
timestamp 1698175906
transform 1 0 28672 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_247
timestamp 1698175906
transform 1 0 29008 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_279
timestamp 1698175906
transform 1 0 32592 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_282
timestamp 1698175906
transform 1 0 32928 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_346
timestamp 1698175906
transform 1 0 40096 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_348
timestamp 1698175906
transform 1 0 40320 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_2
timestamp 1698175906
transform 1 0 1568 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698175906
transform 1 0 5152 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_37
timestamp 1698175906
transform 1 0 5488 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_69
timestamp 1698175906
transform 1 0 9072 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_73
timestamp 1698175906
transform 1 0 9520 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_75
timestamp 1698175906
transform 1 0 9744 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_115
timestamp 1698175906
transform 1 0 14224 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_119
timestamp 1698175906
transform 1 0 14672 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_121
timestamp 1698175906
transform 1 0 14896 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_127
timestamp 1698175906
transform 1 0 15568 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_129
timestamp 1698175906
transform 1 0 15792 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_153
timestamp 1698175906
transform 1 0 18480 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_155
timestamp 1698175906
transform 1 0 18704 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_161
timestamp 1698175906
transform 1 0 19376 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_184
timestamp 1698175906
transform 1 0 21952 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_219
timestamp 1698175906
transform 1 0 25872 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_235
timestamp 1698175906
transform 1 0 27664 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_276
timestamp 1698175906
transform 1 0 32256 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_308
timestamp 1698175906
transform 1 0 35840 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_312
timestamp 1698175906
transform 1 0 36288 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_314
timestamp 1698175906
transform 1 0 36512 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_317
timestamp 1698175906
transform 1 0 36848 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_28
timestamp 1698175906
transform 1 0 4480 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_60
timestamp 1698175906
transform 1 0 8064 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_68
timestamp 1698175906
transform 1 0 8960 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_72
timestamp 1698175906
transform 1 0 9408 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_104
timestamp 1698175906
transform 1 0 12992 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_107
timestamp 1698175906
transform 1 0 13328 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_113
timestamp 1698175906
transform 1 0 14000 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_129
timestamp 1698175906
transform 1 0 15792 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_139
timestamp 1698175906
transform 1 0 16912 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_225
timestamp 1698175906
transform 1 0 26544 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_260
timestamp 1698175906
transform 1 0 30464 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_264
timestamp 1698175906
transform 1 0 30912 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_282
timestamp 1698175906
transform 1 0 32928 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_314
timestamp 1698175906
transform 1 0 36512 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_322
timestamp 1698175906
transform 1 0 37408 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_2
timestamp 1698175906
transform 1 0 1568 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698175906
transform 1 0 5152 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_37
timestamp 1698175906
transform 1 0 5488 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_101
timestamp 1698175906
transform 1 0 12656 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_107
timestamp 1698175906
transform 1 0 13328 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_117
timestamp 1698175906
transform 1 0 14448 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_125
timestamp 1698175906
transform 1 0 15344 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_252
timestamp 1698175906
transform 1 0 29568 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_284
timestamp 1698175906
transform 1 0 33152 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_300
timestamp 1698175906
transform 1 0 34944 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_308
timestamp 1698175906
transform 1 0 35840 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_312
timestamp 1698175906
transform 1 0 36288 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_314
timestamp 1698175906
transform 1 0 36512 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_317
timestamp 1698175906
transform 1 0 36848 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_321
timestamp 1698175906
transform 1 0 37296 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_2
timestamp 1698175906
transform 1 0 1568 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_66
timestamp 1698175906
transform 1 0 8736 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_72
timestamp 1698175906
transform 1 0 9408 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_80
timestamp 1698175906
transform 1 0 10304 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_84
timestamp 1698175906
transform 1 0 10752 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_131
timestamp 1698175906
transform 1 0 16016 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_139
timestamp 1698175906
transform 1 0 16912 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_206
timestamp 1698175906
transform 1 0 24416 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_212
timestamp 1698175906
transform 1 0 25088 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_225
timestamp 1698175906
transform 1 0 26544 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_235
timestamp 1698175906
transform 1 0 27664 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_243
timestamp 1698175906
transform 1 0 28560 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_247
timestamp 1698175906
transform 1 0 29008 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_251
timestamp 1698175906
transform 1 0 29456 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_258
timestamp 1698175906
transform 1 0 30240 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_274
timestamp 1698175906
transform 1 0 32032 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_278
timestamp 1698175906
transform 1 0 32480 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_282
timestamp 1698175906
transform 1 0 32928 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_314
timestamp 1698175906
transform 1 0 36512 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_322
timestamp 1698175906
transform 1 0 37408 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_2
timestamp 1698175906
transform 1 0 1568 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698175906
transform 1 0 5152 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_37
timestamp 1698175906
transform 1 0 5488 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_101
timestamp 1698175906
transform 1 0 12656 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_107
timestamp 1698175906
transform 1 0 13328 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_115
timestamp 1698175906
transform 1 0 14224 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_141
timestamp 1698175906
transform 1 0 17136 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_148
timestamp 1698175906
transform 1 0 17920 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_156
timestamp 1698175906
transform 1 0 18816 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_163
timestamp 1698175906
transform 1 0 19600 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_167
timestamp 1698175906
transform 1 0 20048 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_177
timestamp 1698175906
transform 1 0 21168 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_179
timestamp 1698175906
transform 1 0 21392 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_186
timestamp 1698175906
transform 1 0 22176 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_188
timestamp 1698175906
transform 1 0 22400 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_218
timestamp 1698175906
transform 1 0 25760 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_222
timestamp 1698175906
transform 1 0 26208 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_230
timestamp 1698175906
transform 1 0 27104 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_234
timestamp 1698175906
transform 1 0 27552 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_236
timestamp 1698175906
transform 1 0 27776 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_276
timestamp 1698175906
transform 1 0 32256 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_308
timestamp 1698175906
transform 1 0 35840 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_312
timestamp 1698175906
transform 1 0 36288 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_314
timestamp 1698175906
transform 1 0 36512 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_317
timestamp 1698175906
transform 1 0 36848 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_321
timestamp 1698175906
transform 1 0 37296 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_2
timestamp 1698175906
transform 1 0 1568 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_66
timestamp 1698175906
transform 1 0 8736 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_72
timestamp 1698175906
transform 1 0 9408 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_104
timestamp 1698175906
transform 1 0 12992 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_107
timestamp 1698175906
transform 1 0 13328 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_111
timestamp 1698175906
transform 1 0 13776 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_121
timestamp 1698175906
transform 1 0 14896 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_138
timestamp 1698175906
transform 1 0 16800 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_142
timestamp 1698175906
transform 1 0 17248 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_158
timestamp 1698175906
transform 1 0 19040 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_166
timestamp 1698175906
transform 1 0 19936 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_168
timestamp 1698175906
transform 1 0 20160 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_175
timestamp 1698175906
transform 1 0 20944 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_180
timestamp 1698175906
transform 1 0 21504 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_187
timestamp 1698175906
transform 1 0 22288 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_191
timestamp 1698175906
transform 1 0 22736 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_197
timestamp 1698175906
transform 1 0 23408 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_205
timestamp 1698175906
transform 1 0 24304 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_209
timestamp 1698175906
transform 1 0 24752 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_212
timestamp 1698175906
transform 1 0 25088 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_226
timestamp 1698175906
transform 1 0 26656 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_258
timestamp 1698175906
transform 1 0 30240 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_274
timestamp 1698175906
transform 1 0 32032 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_278
timestamp 1698175906
transform 1 0 32480 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_282
timestamp 1698175906
transform 1 0 32928 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_346
timestamp 1698175906
transform 1 0 40096 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_348
timestamp 1698175906
transform 1 0 40320 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_28
timestamp 1698175906
transform 1 0 4480 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_32
timestamp 1698175906
transform 1 0 4928 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698175906
transform 1 0 5152 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_37
timestamp 1698175906
transform 1 0 5488 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_69
timestamp 1698175906
transform 1 0 9072 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_73
timestamp 1698175906
transform 1 0 9520 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_75
timestamp 1698175906
transform 1 0 9744 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_113
timestamp 1698175906
transform 1 0 14000 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_117
timestamp 1698175906
transform 1 0 14448 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_121
timestamp 1698175906
transform 1 0 14896 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_153
timestamp 1698175906
transform 1 0 18480 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_166
timestamp 1698175906
transform 1 0 19936 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_174
timestamp 1698175906
transform 1 0 20832 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_177
timestamp 1698175906
transform 1 0 21168 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_209
timestamp 1698175906
transform 1 0 24752 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_217
timestamp 1698175906
transform 1 0 25648 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_221
timestamp 1698175906
transform 1 0 26096 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_230
timestamp 1698175906
transform 1 0 27104 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_244
timestamp 1698175906
transform 1 0 28672 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_247
timestamp 1698175906
transform 1 0 29008 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_311
timestamp 1698175906
transform 1 0 36176 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_317
timestamp 1698175906
transform 1 0 36848 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_2
timestamp 1698175906
transform 1 0 1568 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_66
timestamp 1698175906
transform 1 0 8736 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_72
timestamp 1698175906
transform 1 0 9408 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_88
timestamp 1698175906
transform 1 0 11200 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_127
timestamp 1698175906
transform 1 0 15568 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_135
timestamp 1698175906
transform 1 0 16464 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_139
timestamp 1698175906
transform 1 0 16912 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_142
timestamp 1698175906
transform 1 0 17248 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_146
timestamp 1698175906
transform 1 0 17696 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_177
timestamp 1698175906
transform 1 0 21168 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_181
timestamp 1698175906
transform 1 0 21616 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_185
timestamp 1698175906
transform 1 0 22064 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_187
timestamp 1698175906
transform 1 0 22288 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_194
timestamp 1698175906
transform 1 0 23072 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_212
timestamp 1698175906
transform 1 0 25088 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_239
timestamp 1698175906
transform 1 0 28112 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_252
timestamp 1698175906
transform 1 0 29568 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_268
timestamp 1698175906
transform 1 0 31360 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_276
timestamp 1698175906
transform 1 0 32256 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_282
timestamp 1698175906
transform 1 0 32928 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_346
timestamp 1698175906
transform 1 0 40096 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_348
timestamp 1698175906
transform 1 0 40320 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_28
timestamp 1698175906
transform 1 0 4480 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_32
timestamp 1698175906
transform 1 0 4928 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698175906
transform 1 0 5152 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_37
timestamp 1698175906
transform 1 0 5488 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_101
timestamp 1698175906
transform 1 0 12656 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_107
timestamp 1698175906
transform 1 0 13328 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_111
timestamp 1698175906
transform 1 0 13776 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_113
timestamp 1698175906
transform 1 0 14000 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_119
timestamp 1698175906
transform 1 0 14672 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_133
timestamp 1698175906
transform 1 0 16240 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_165
timestamp 1698175906
transform 1 0 19824 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_199
timestamp 1698175906
transform 1 0 23632 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_207
timestamp 1698175906
transform 1 0 24528 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_243
timestamp 1698175906
transform 1 0 28560 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_276
timestamp 1698175906
transform 1 0 32256 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_308
timestamp 1698175906
transform 1 0 35840 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_312
timestamp 1698175906
transform 1 0 36288 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_314
timestamp 1698175906
transform 1 0 36512 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_317
timestamp 1698175906
transform 1 0 36848 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_321
timestamp 1698175906
transform 1 0 37296 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_28
timestamp 1698175906
transform 1 0 4480 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_60
timestamp 1698175906
transform 1 0 8064 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_68
timestamp 1698175906
transform 1 0 8960 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_72
timestamp 1698175906
transform 1 0 9408 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_88
timestamp 1698175906
transform 1 0 11200 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_96
timestamp 1698175906
transform 1 0 12096 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_100
timestamp 1698175906
transform 1 0 12544 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_130
timestamp 1698175906
transform 1 0 15904 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_134
timestamp 1698175906
transform 1 0 16352 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_138
timestamp 1698175906
transform 1 0 16800 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_147
timestamp 1698175906
transform 1 0 17808 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_151
timestamp 1698175906
transform 1 0 18256 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_157
timestamp 1698175906
transform 1 0 18928 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_161
timestamp 1698175906
transform 1 0 19376 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_165
timestamp 1698175906
transform 1 0 19824 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_198
timestamp 1698175906
transform 1 0 23520 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_206
timestamp 1698175906
transform 1 0 24416 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_212
timestamp 1698175906
transform 1 0 25088 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_214
timestamp 1698175906
transform 1 0 25312 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_244
timestamp 1698175906
transform 1 0 28672 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_249
timestamp 1698175906
transform 1 0 29232 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_253
timestamp 1698175906
transform 1 0 29680 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_257
timestamp 1698175906
transform 1 0 30128 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_273
timestamp 1698175906
transform 1 0 31920 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_277
timestamp 1698175906
transform 1 0 32368 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_279
timestamp 1698175906
transform 1 0 32592 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_282
timestamp 1698175906
transform 1 0 32928 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_314
timestamp 1698175906
transform 1 0 36512 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_322
timestamp 1698175906
transform 1 0 37408 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_2
timestamp 1698175906
transform 1 0 1568 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698175906
transform 1 0 5152 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_37
timestamp 1698175906
transform 1 0 5488 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_101
timestamp 1698175906
transform 1 0 12656 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_107
timestamp 1698175906
transform 1 0 13328 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_123
timestamp 1698175906
transform 1 0 15120 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_127
timestamp 1698175906
transform 1 0 15568 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_158
timestamp 1698175906
transform 1 0 19040 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_170
timestamp 1698175906
transform 1 0 20384 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_174
timestamp 1698175906
transform 1 0 20832 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_177
timestamp 1698175906
transform 1 0 21168 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_184
timestamp 1698175906
transform 1 0 21952 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_186
timestamp 1698175906
transform 1 0 22176 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_192
timestamp 1698175906
transform 1 0 22848 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_194
timestamp 1698175906
transform 1 0 23072 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_201
timestamp 1698175906
transform 1 0 23856 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_233
timestamp 1698175906
transform 1 0 27440 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_241
timestamp 1698175906
transform 1 0 28336 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_247
timestamp 1698175906
transform 1 0 29008 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_311
timestamp 1698175906
transform 1 0 36176 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_317
timestamp 1698175906
transform 1 0 36848 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_321
timestamp 1698175906
transform 1 0 37296 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_2
timestamp 1698175906
transform 1 0 1568 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_66
timestamp 1698175906
transform 1 0 8736 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_72
timestamp 1698175906
transform 1 0 9408 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_136
timestamp 1698175906
transform 1 0 16576 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_171
timestamp 1698175906
transform 1 0 20496 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_175
timestamp 1698175906
transform 1 0 20944 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_207
timestamp 1698175906
transform 1 0 24528 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_209
timestamp 1698175906
transform 1 0 24752 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_212
timestamp 1698175906
transform 1 0 25088 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_216
timestamp 1698175906
transform 1 0 25536 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_282
timestamp 1698175906
transform 1 0 32928 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_346
timestamp 1698175906
transform 1 0 40096 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_348
timestamp 1698175906
transform 1 0 40320 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_2
timestamp 1698175906
transform 1 0 1568 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698175906
transform 1 0 5152 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_37
timestamp 1698175906
transform 1 0 5488 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_101
timestamp 1698175906
transform 1 0 12656 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_107
timestamp 1698175906
transform 1 0 13328 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_171
timestamp 1698175906
transform 1 0 20496 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_177
timestamp 1698175906
transform 1 0 21168 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_193
timestamp 1698175906
transform 1 0 22960 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_201
timestamp 1698175906
transform 1 0 23856 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_233
timestamp 1698175906
transform 1 0 27440 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_241
timestamp 1698175906
transform 1 0 28336 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_247
timestamp 1698175906
transform 1 0 29008 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_311
timestamp 1698175906
transform 1 0 36176 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_317
timestamp 1698175906
transform 1 0 36848 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_2
timestamp 1698175906
transform 1 0 1568 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_66
timestamp 1698175906
transform 1 0 8736 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_72
timestamp 1698175906
transform 1 0 9408 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_136
timestamp 1698175906
transform 1 0 16576 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_142
timestamp 1698175906
transform 1 0 17248 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_206
timestamp 1698175906
transform 1 0 24416 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_212
timestamp 1698175906
transform 1 0 25088 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_276
timestamp 1698175906
transform 1 0 32256 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_282
timestamp 1698175906
transform 1 0 32928 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_346
timestamp 1698175906
transform 1 0 40096 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_348
timestamp 1698175906
transform 1 0 40320 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698175906
transform 1 0 1568 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698175906
transform 1 0 5152 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_37
timestamp 1698175906
transform 1 0 5488 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_101
timestamp 1698175906
transform 1 0 12656 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_107
timestamp 1698175906
transform 1 0 13328 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_171
timestamp 1698175906
transform 1 0 20496 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_177
timestamp 1698175906
transform 1 0 21168 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_241
timestamp 1698175906
transform 1 0 28336 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_247
timestamp 1698175906
transform 1 0 29008 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_311
timestamp 1698175906
transform 1 0 36176 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_317
timestamp 1698175906
transform 1 0 36848 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2
timestamp 1698175906
transform 1 0 1568 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_66
timestamp 1698175906
transform 1 0 8736 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_72
timestamp 1698175906
transform 1 0 9408 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_136
timestamp 1698175906
transform 1 0 16576 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_142
timestamp 1698175906
transform 1 0 17248 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_206
timestamp 1698175906
transform 1 0 24416 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_212
timestamp 1698175906
transform 1 0 25088 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_276
timestamp 1698175906
transform 1 0 32256 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_282
timestamp 1698175906
transform 1 0 32928 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_346
timestamp 1698175906
transform 1 0 40096 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_348
timestamp 1698175906
transform 1 0 40320 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_2
timestamp 1698175906
transform 1 0 1568 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698175906
transform 1 0 5152 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_37
timestamp 1698175906
transform 1 0 5488 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_101
timestamp 1698175906
transform 1 0 12656 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_107
timestamp 1698175906
transform 1 0 13328 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_171
timestamp 1698175906
transform 1 0 20496 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_177
timestamp 1698175906
transform 1 0 21168 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_241
timestamp 1698175906
transform 1 0 28336 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_247
timestamp 1698175906
transform 1 0 29008 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_311
timestamp 1698175906
transform 1 0 36176 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_317
timestamp 1698175906
transform 1 0 36848 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2
timestamp 1698175906
transform 1 0 1568 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_66
timestamp 1698175906
transform 1 0 8736 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_72
timestamp 1698175906
transform 1 0 9408 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_136
timestamp 1698175906
transform 1 0 16576 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_142
timestamp 1698175906
transform 1 0 17248 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_206
timestamp 1698175906
transform 1 0 24416 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_212
timestamp 1698175906
transform 1 0 25088 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_276
timestamp 1698175906
transform 1 0 32256 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_282
timestamp 1698175906
transform 1 0 32928 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_346
timestamp 1698175906
transform 1 0 40096 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_348
timestamp 1698175906
transform 1 0 40320 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698175906
transform 1 0 1568 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698175906
transform 1 0 5152 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_37
timestamp 1698175906
transform 1 0 5488 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_101
timestamp 1698175906
transform 1 0 12656 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_107
timestamp 1698175906
transform 1 0 13328 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_171
timestamp 1698175906
transform 1 0 20496 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_177
timestamp 1698175906
transform 1 0 21168 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_241
timestamp 1698175906
transform 1 0 28336 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_247
timestamp 1698175906
transform 1 0 29008 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_311
timestamp 1698175906
transform 1 0 36176 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_317
timestamp 1698175906
transform 1 0 36848 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_2
timestamp 1698175906
transform 1 0 1568 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_66
timestamp 1698175906
transform 1 0 8736 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_72
timestamp 1698175906
transform 1 0 9408 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_136
timestamp 1698175906
transform 1 0 16576 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_142
timestamp 1698175906
transform 1 0 17248 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_206
timestamp 1698175906
transform 1 0 24416 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_212
timestamp 1698175906
transform 1 0 25088 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_276
timestamp 1698175906
transform 1 0 32256 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_282
timestamp 1698175906
transform 1 0 32928 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_346
timestamp 1698175906
transform 1 0 40096 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_348
timestamp 1698175906
transform 1 0 40320 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698175906
transform 1 0 1568 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698175906
transform 1 0 5152 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_37
timestamp 1698175906
transform 1 0 5488 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_101
timestamp 1698175906
transform 1 0 12656 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_107
timestamp 1698175906
transform 1 0 13328 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_171
timestamp 1698175906
transform 1 0 20496 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_177
timestamp 1698175906
transform 1 0 21168 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_241
timestamp 1698175906
transform 1 0 28336 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_247
timestamp 1698175906
transform 1 0 29008 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_311
timestamp 1698175906
transform 1 0 36176 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_317
timestamp 1698175906
transform 1 0 36848 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2
timestamp 1698175906
transform 1 0 1568 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1698175906
transform 1 0 8736 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_72
timestamp 1698175906
transform 1 0 9408 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_136
timestamp 1698175906
transform 1 0 16576 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_142
timestamp 1698175906
transform 1 0 17248 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_206
timestamp 1698175906
transform 1 0 24416 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_212
timestamp 1698175906
transform 1 0 25088 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_276
timestamp 1698175906
transform 1 0 32256 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_282
timestamp 1698175906
transform 1 0 32928 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_346
timestamp 1698175906
transform 1 0 40096 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_348
timestamp 1698175906
transform 1 0 40320 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_2
timestamp 1698175906
transform 1 0 1568 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698175906
transform 1 0 5152 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_37
timestamp 1698175906
transform 1 0 5488 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_101
timestamp 1698175906
transform 1 0 12656 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_107
timestamp 1698175906
transform 1 0 13328 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_171
timestamp 1698175906
transform 1 0 20496 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_177
timestamp 1698175906
transform 1 0 21168 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_193
timestamp 1698175906
transform 1 0 22960 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_197
timestamp 1698175906
transform 1 0 23408 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_225
timestamp 1698175906
transform 1 0 26544 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_241
timestamp 1698175906
transform 1 0 28336 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_247
timestamp 1698175906
transform 1 0 29008 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_311
timestamp 1698175906
transform 1 0 36176 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_317
timestamp 1698175906
transform 1 0 36848 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_2
timestamp 1698175906
transform 1 0 1568 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_66
timestamp 1698175906
transform 1 0 8736 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_72
timestamp 1698175906
transform 1 0 9408 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_136
timestamp 1698175906
transform 1 0 16576 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_142
timestamp 1698175906
transform 1 0 17248 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_158
timestamp 1698175906
transform 1 0 19040 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_166
timestamp 1698175906
transform 1 0 19936 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_168
timestamp 1698175906
transform 1 0 20160 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_195
timestamp 1698175906
transform 1 0 23184 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_203
timestamp 1698175906
transform 1 0 24080 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_207
timestamp 1698175906
transform 1 0 24528 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_209
timestamp 1698175906
transform 1 0 24752 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_238
timestamp 1698175906
transform 1 0 28000 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_270
timestamp 1698175906
transform 1 0 31584 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_278
timestamp 1698175906
transform 1 0 32480 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_282
timestamp 1698175906
transform 1 0 32928 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_346
timestamp 1698175906
transform 1 0 40096 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_348
timestamp 1698175906
transform 1 0 40320 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_2
timestamp 1698175906
transform 1 0 1568 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_36
timestamp 1698175906
transform 1 0 5376 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_70
timestamp 1698175906
transform 1 0 9184 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_104
timestamp 1698175906
transform 1 0 12992 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_138
timestamp 1698175906
transform 1 0 16800 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_142
timestamp 1698175906
transform 1 0 17248 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_172
timestamp 1698175906
transform 1 0 20608 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_176
timestamp 1698175906
transform 1 0 21056 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_232
timestamp 1698175906
transform 1 0 27328 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_236
timestamp 1698175906
transform 1 0 27776 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_240
timestamp 1698175906
transform 1 0 28224 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_274
timestamp 1698175906
transform 1 0 32032 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_308
timestamp 1698175906
transform 1 0 35840 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_342
timestamp 1698175906
transform 1 0 39648 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_346
timestamp 1698175906
transform 1 0 40096 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_348
timestamp 1698175906
transform 1 0 40320 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 25088 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output2
timestamp 1698175906
transform 1 0 24416 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output3
timestamp 1698175906
transform 1 0 24416 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output4
timestamp 1698175906
transform 1 0 37520 0 1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output5
timestamp 1698175906
transform 1 0 37520 0 -1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output6
timestamp 1698175906
transform 1 0 28560 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output7
timestamp 1698175906
transform -1 0 4480 0 1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output8
timestamp 1698175906
transform -1 0 24192 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output9
timestamp 1698175906
transform 1 0 25648 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output10
timestamp 1698175906
transform -1 0 4480 0 -1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output11
timestamp 1698175906
transform 1 0 37520 0 -1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output12
timestamp 1698175906
transform 1 0 37520 0 1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output13
timestamp 1698175906
transform 1 0 37520 0 1 14112
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output14
timestamp 1698175906
transform 1 0 37520 0 1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output15
timestamp 1698175906
transform -1 0 4480 0 -1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output16
timestamp 1698175906
transform 1 0 37520 0 1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output17
timestamp 1698175906
transform 1 0 37520 0 -1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output18
timestamp 1698175906
transform -1 0 4480 0 -1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output19
timestamp 1698175906
transform 1 0 17472 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output20
timestamp 1698175906
transform 1 0 21280 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output21
timestamp 1698175906
transform 1 0 37520 0 -1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output22
timestamp 1698175906
transform -1 0 4480 0 1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output23
timestamp 1698175906
transform 1 0 28224 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output24
timestamp 1698175906
transform 1 0 20272 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output25
timestamp 1698175906
transform 1 0 23632 0 1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output26
timestamp 1698175906
transform 1 0 37520 0 1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_45 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698175906
transform -1 0 40656 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_46
timestamp 1698175906
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698175906
transform -1 0 40656 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_47
timestamp 1698175906
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698175906
transform -1 0 40656 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_48
timestamp 1698175906
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698175906
transform -1 0 40656 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_49
timestamp 1698175906
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698175906
transform -1 0 40656 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_50
timestamp 1698175906
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698175906
transform -1 0 40656 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_51
timestamp 1698175906
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698175906
transform -1 0 40656 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_52
timestamp 1698175906
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698175906
transform -1 0 40656 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_53
timestamp 1698175906
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698175906
transform -1 0 40656 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_54
timestamp 1698175906
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698175906
transform -1 0 40656 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_55
timestamp 1698175906
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698175906
transform -1 0 40656 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_56
timestamp 1698175906
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698175906
transform -1 0 40656 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_57
timestamp 1698175906
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698175906
transform -1 0 40656 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_58
timestamp 1698175906
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698175906
transform -1 0 40656 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_59
timestamp 1698175906
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698175906
transform -1 0 40656 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_60
timestamp 1698175906
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698175906
transform -1 0 40656 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_61
timestamp 1698175906
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698175906
transform -1 0 40656 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_62
timestamp 1698175906
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698175906
transform -1 0 40656 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_63
timestamp 1698175906
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698175906
transform -1 0 40656 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_64
timestamp 1698175906
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698175906
transform -1 0 40656 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_65
timestamp 1698175906
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698175906
transform -1 0 40656 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_66
timestamp 1698175906
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698175906
transform -1 0 40656 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_67
timestamp 1698175906
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698175906
transform -1 0 40656 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_68
timestamp 1698175906
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698175906
transform -1 0 40656 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_69
timestamp 1698175906
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698175906
transform -1 0 40656 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_70
timestamp 1698175906
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698175906
transform -1 0 40656 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_71
timestamp 1698175906
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698175906
transform -1 0 40656 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_72
timestamp 1698175906
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698175906
transform -1 0 40656 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_73
timestamp 1698175906
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698175906
transform -1 0 40656 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_74
timestamp 1698175906
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698175906
transform -1 0 40656 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_75
timestamp 1698175906
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698175906
transform -1 0 40656 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_76
timestamp 1698175906
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698175906
transform -1 0 40656 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_77
timestamp 1698175906
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698175906
transform -1 0 40656 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_78
timestamp 1698175906
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698175906
transform -1 0 40656 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_79
timestamp 1698175906
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698175906
transform -1 0 40656 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_80
timestamp 1698175906
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698175906
transform -1 0 40656 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_81
timestamp 1698175906
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698175906
transform -1 0 40656 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_82
timestamp 1698175906
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698175906
transform -1 0 40656 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_83
timestamp 1698175906
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698175906
transform -1 0 40656 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_84
timestamp 1698175906
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698175906
transform -1 0 40656 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_85
timestamp 1698175906
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698175906
transform -1 0 40656 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_86
timestamp 1698175906
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698175906
transform -1 0 40656 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_87
timestamp 1698175906
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698175906
transform -1 0 40656 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_88
timestamp 1698175906
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698175906
transform -1 0 40656 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_89
timestamp 1698175906
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698175906
transform -1 0 40656 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_90 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_91
timestamp 1698175906
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_92
timestamp 1698175906
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_93
timestamp 1698175906
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_94
timestamp 1698175906
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_95
timestamp 1698175906
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_96
timestamp 1698175906
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_97
timestamp 1698175906
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_98
timestamp 1698175906
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_99
timestamp 1698175906
transform 1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_100
timestamp 1698175906
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_101
timestamp 1698175906
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_102
timestamp 1698175906
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_103
timestamp 1698175906
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_104
timestamp 1698175906
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_105
timestamp 1698175906
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_106
timestamp 1698175906
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_107
timestamp 1698175906
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_108
timestamp 1698175906
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_109
timestamp 1698175906
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_110
timestamp 1698175906
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_111
timestamp 1698175906
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_112
timestamp 1698175906
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_113
timestamp 1698175906
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_114
timestamp 1698175906
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_115
timestamp 1698175906
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_116
timestamp 1698175906
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_117
timestamp 1698175906
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_118
timestamp 1698175906
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_119
timestamp 1698175906
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_120
timestamp 1698175906
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_121
timestamp 1698175906
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_122
timestamp 1698175906
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_123
timestamp 1698175906
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_124
timestamp 1698175906
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_125
timestamp 1698175906
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_126
timestamp 1698175906
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_127
timestamp 1698175906
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_128
timestamp 1698175906
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_129
timestamp 1698175906
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_130
timestamp 1698175906
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_131
timestamp 1698175906
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_132
timestamp 1698175906
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_133
timestamp 1698175906
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_134
timestamp 1698175906
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_135
timestamp 1698175906
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_136
timestamp 1698175906
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_137
timestamp 1698175906
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_138
timestamp 1698175906
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_139
timestamp 1698175906
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_140
timestamp 1698175906
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_141
timestamp 1698175906
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_142
timestamp 1698175906
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_143
timestamp 1698175906
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_144
timestamp 1698175906
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_145
timestamp 1698175906
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_146
timestamp 1698175906
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_147
timestamp 1698175906
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_148
timestamp 1698175906
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_149
timestamp 1698175906
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_150
timestamp 1698175906
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_151
timestamp 1698175906
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_152
timestamp 1698175906
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_153
timestamp 1698175906
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_154
timestamp 1698175906
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_155
timestamp 1698175906
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_156
timestamp 1698175906
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_157
timestamp 1698175906
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_158
timestamp 1698175906
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_159
timestamp 1698175906
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_160
timestamp 1698175906
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_161
timestamp 1698175906
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_162
timestamp 1698175906
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_163
timestamp 1698175906
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_164
timestamp 1698175906
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_165
timestamp 1698175906
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_166
timestamp 1698175906
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_167
timestamp 1698175906
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_168
timestamp 1698175906
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_169
timestamp 1698175906
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_170
timestamp 1698175906
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_171
timestamp 1698175906
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_172
timestamp 1698175906
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_173
timestamp 1698175906
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_174
timestamp 1698175906
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_175
timestamp 1698175906
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_176
timestamp 1698175906
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_177
timestamp 1698175906
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_178
timestamp 1698175906
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_179
timestamp 1698175906
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_180
timestamp 1698175906
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_181
timestamp 1698175906
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_182
timestamp 1698175906
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_183
timestamp 1698175906
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_184
timestamp 1698175906
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_185
timestamp 1698175906
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_186
timestamp 1698175906
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_187
timestamp 1698175906
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_188
timestamp 1698175906
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_189
timestamp 1698175906
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_190
timestamp 1698175906
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_191
timestamp 1698175906
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_192
timestamp 1698175906
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_193
timestamp 1698175906
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_194
timestamp 1698175906
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_195
timestamp 1698175906
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_196
timestamp 1698175906
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_197
timestamp 1698175906
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_198
timestamp 1698175906
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_199
timestamp 1698175906
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_200
timestamp 1698175906
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_201
timestamp 1698175906
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_202
timestamp 1698175906
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_203
timestamp 1698175906
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_204
timestamp 1698175906
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_205
timestamp 1698175906
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_206
timestamp 1698175906
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_207
timestamp 1698175906
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_208
timestamp 1698175906
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_209
timestamp 1698175906
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_210
timestamp 1698175906
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_211
timestamp 1698175906
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_212
timestamp 1698175906
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_213
timestamp 1698175906
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_214
timestamp 1698175906
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_215
timestamp 1698175906
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_216
timestamp 1698175906
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_217
timestamp 1698175906
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_218
timestamp 1698175906
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_219
timestamp 1698175906
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_220
timestamp 1698175906
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_221
timestamp 1698175906
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_222
timestamp 1698175906
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_223
timestamp 1698175906
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_224
timestamp 1698175906
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_225
timestamp 1698175906
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_226
timestamp 1698175906
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_227
timestamp 1698175906
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_228
timestamp 1698175906
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_229
timestamp 1698175906
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_230
timestamp 1698175906
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_231
timestamp 1698175906
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_232
timestamp 1698175906
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_233
timestamp 1698175906
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_234
timestamp 1698175906
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_235
timestamp 1698175906
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_236
timestamp 1698175906
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_237
timestamp 1698175906
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_238
timestamp 1698175906
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_239
timestamp 1698175906
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_240
timestamp 1698175906
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_241
timestamp 1698175906
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_242
timestamp 1698175906
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_243
timestamp 1698175906
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_244
timestamp 1698175906
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_245
timestamp 1698175906
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_246
timestamp 1698175906
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_247
timestamp 1698175906
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_248
timestamp 1698175906
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_249
timestamp 1698175906
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_250
timestamp 1698175906
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_251
timestamp 1698175906
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_252
timestamp 1698175906
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_253
timestamp 1698175906
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_254
timestamp 1698175906
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_255
timestamp 1698175906
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_256
timestamp 1698175906
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_257
timestamp 1698175906
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_258
timestamp 1698175906
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_259
timestamp 1698175906
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_260
timestamp 1698175906
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_261
timestamp 1698175906
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_262
timestamp 1698175906
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_263
timestamp 1698175906
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_264
timestamp 1698175906
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_265
timestamp 1698175906
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_266
timestamp 1698175906
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_267
timestamp 1698175906
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_268
timestamp 1698175906
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_269
timestamp 1698175906
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_270
timestamp 1698175906
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_271
timestamp 1698175906
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_272
timestamp 1698175906
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_273
timestamp 1698175906
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_274
timestamp 1698175906
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_275
timestamp 1698175906
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_276
timestamp 1698175906
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_277
timestamp 1698175906
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_278
timestamp 1698175906
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_279
timestamp 1698175906
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_280
timestamp 1698175906
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_281
timestamp 1698175906
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_282
timestamp 1698175906
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_283
timestamp 1698175906
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_284
timestamp 1698175906
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_285
timestamp 1698175906
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_286
timestamp 1698175906
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_287
timestamp 1698175906
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_288
timestamp 1698175906
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_289
timestamp 1698175906
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_290
timestamp 1698175906
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_291
timestamp 1698175906
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_292
timestamp 1698175906
transform 1 0 32704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_293
timestamp 1698175906
transform 1 0 5152 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_294
timestamp 1698175906
transform 1 0 8960 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_295
timestamp 1698175906
transform 1 0 12768 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_296
timestamp 1698175906
transform 1 0 16576 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_297
timestamp 1698175906
transform 1 0 20384 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_298
timestamp 1698175906
transform 1 0 24192 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_299
timestamp 1698175906
transform 1 0 28000 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_300
timestamp 1698175906
transform 1 0 31808 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_301
timestamp 1698175906
transform 1 0 35616 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_302
timestamp 1698175906
transform 1 0 39424 0 1 37632
box -86 -86 310 870
<< labels >>
flabel metal3 s 0 27552 800 27664 0 FreeSans 448 0 0 0 clk
port 0 nsew signal input
flabel metal2 s 24192 41200 24304 42000 0 FreeSans 448 90 0 0 segm[0]
port 1 nsew signal tristate
flabel metal2 s 24192 0 24304 800 0 FreeSans 448 90 0 0 segm[10]
port 2 nsew signal tristate
flabel metal2 s 22848 41200 22960 42000 0 FreeSans 448 90 0 0 segm[11]
port 3 nsew signal tristate
flabel metal3 s 41200 17472 42000 17584 0 FreeSans 448 0 0 0 segm[12]
port 4 nsew signal tristate
flabel metal3 s 41200 16800 42000 16912 0 FreeSans 448 0 0 0 segm[13]
port 5 nsew signal tristate
flabel metal2 s 26880 0 26992 800 0 FreeSans 448 90 0 0 segm[1]
port 6 nsew signal tristate
flabel metal3 s 0 24864 800 24976 0 FreeSans 448 0 0 0 segm[2]
port 7 nsew signal tristate
flabel metal2 s 22176 41200 22288 42000 0 FreeSans 448 90 0 0 segm[3]
port 8 nsew signal tristate
flabel metal2 s 25536 0 25648 800 0 FreeSans 448 90 0 0 segm[4]
port 9 nsew signal tristate
flabel metal3 s 0 25536 800 25648 0 FreeSans 448 0 0 0 segm[5]
port 10 nsew signal tristate
flabel metal3 s 41200 21504 42000 21616 0 FreeSans 448 0 0 0 segm[6]
port 11 nsew signal tristate
flabel metal3 s 41200 26208 42000 26320 0 FreeSans 448 0 0 0 segm[7]
port 12 nsew signal tristate
flabel metal3 s 41200 14112 42000 14224 0 FreeSans 448 0 0 0 segm[8]
port 13 nsew signal tristate
flabel metal3 s 41200 24864 42000 24976 0 FreeSans 448 0 0 0 segm[9]
port 14 nsew signal tristate
flabel metal3 s 0 18144 800 18256 0 FreeSans 448 0 0 0 sel[0]
port 15 nsew signal tristate
flabel metal3 s 41200 22176 42000 22288 0 FreeSans 448 0 0 0 sel[10]
port 16 nsew signal tristate
flabel metal3 s 41200 25536 42000 25648 0 FreeSans 448 0 0 0 sel[11]
port 17 nsew signal tristate
flabel metal3 s 0 19488 800 19600 0 FreeSans 448 0 0 0 sel[1]
port 18 nsew signal tristate
flabel metal2 s 18816 41200 18928 42000 0 FreeSans 448 90 0 0 sel[2]
port 19 nsew signal tristate
flabel metal2 s 21504 0 21616 800 0 FreeSans 448 90 0 0 sel[3]
port 20 nsew signal tristate
flabel metal3 s 41200 19488 42000 19600 0 FreeSans 448 0 0 0 sel[4]
port 21 nsew signal tristate
flabel metal3 s 0 23520 800 23632 0 FreeSans 448 0 0 0 sel[5]
port 22 nsew signal tristate
flabel metal2 s 26208 0 26320 800 0 FreeSans 448 90 0 0 sel[6]
port 23 nsew signal tristate
flabel metal2 s 20160 41200 20272 42000 0 FreeSans 448 90 0 0 sel[7]
port 24 nsew signal tristate
flabel metal2 s 23520 41200 23632 42000 0 FreeSans 448 90 0 0 sel[8]
port 25 nsew signal tristate
flabel metal3 s 41200 20832 42000 20944 0 FreeSans 448 0 0 0 sel[9]
port 26 nsew signal tristate
flabel metal4 s 4448 3076 4768 38476 0 FreeSans 1280 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 35168 3076 35488 38476 0 FreeSans 1280 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 19808 3076 20128 38476 0 FreeSans 1280 90 0 0 vss
port 28 nsew ground bidirectional
rlabel metal1 21000 38416 21000 38416 0 vdd
rlabel metal1 21000 37632 21000 37632 0 vss
rlabel metal2 20104 27496 20104 27496 0 _000_
rlabel metal3 12880 24024 12880 24024 0 _001_
rlabel metal3 14336 24808 14336 24808 0 _002_
rlabel metal2 15232 25256 15232 25256 0 _003_
rlabel metal3 29064 19096 29064 19096 0 _004_
rlabel metal2 13272 21896 13272 21896 0 _005_
rlabel metal2 15512 17304 15512 17304 0 _006_
rlabel metal2 18424 15512 18424 15512 0 _007_
rlabel metal2 19656 24808 19656 24808 0 _008_
rlabel metal2 19096 15624 19096 15624 0 _009_
rlabel metal2 17528 26096 17528 26096 0 _010_
rlabel metal3 12880 19096 12880 19096 0 _011_
rlabel metal2 12152 18144 12152 18144 0 _012_
rlabel metal2 23408 22456 23408 22456 0 _013_
rlabel metal2 22344 15624 22344 15624 0 _014_
rlabel metal2 27776 16968 27776 16968 0 _015_
rlabel metal2 28616 15400 28616 15400 0 _016_
rlabel metal2 21672 27496 21672 27496 0 _017_
rlabel metal2 26488 14728 26488 14728 0 _018_
rlabel metal2 23800 13328 23800 13328 0 _019_
rlabel metal3 29064 22232 29064 22232 0 _020_
rlabel metal2 30016 25592 30016 25592 0 _021_
rlabel metal2 26376 25480 26376 25480 0 _022_
rlabel metal2 26320 24024 26320 24024 0 _023_
rlabel metal2 21280 26152 21280 26152 0 _024_
rlabel metal2 27048 20804 27048 20804 0 _025_
rlabel metal2 18200 16072 18200 16072 0 _026_
rlabel metal2 20272 19208 20272 19208 0 _027_
rlabel metal2 25648 20216 25648 20216 0 _028_
rlabel metal2 25312 18984 25312 18984 0 _029_
rlabel metal2 20664 16184 20664 16184 0 _030_
rlabel metal3 17976 26376 17976 26376 0 _031_
rlabel metal2 16744 23968 16744 23968 0 _032_
rlabel metal2 18088 20272 18088 20272 0 _033_
rlabel metal3 14476 19208 14476 19208 0 _034_
rlabel metal2 16632 19544 16632 19544 0 _035_
rlabel metal2 13832 19712 13832 19712 0 _036_
rlabel metal2 13496 19600 13496 19600 0 _037_
rlabel metal2 14336 21336 14336 21336 0 _038_
rlabel metal2 13720 18200 13720 18200 0 _039_
rlabel metal2 15064 18200 15064 18200 0 _040_
rlabel metal2 27608 17920 27608 17920 0 _041_
rlabel metal2 28056 22008 28056 22008 0 _042_
rlabel metal3 20664 21560 20664 21560 0 _043_
rlabel metal2 22568 21280 22568 21280 0 _044_
rlabel metal2 22120 20832 22120 20832 0 _045_
rlabel metal2 22456 21448 22456 21448 0 _046_
rlabel metal3 20776 17752 20776 17752 0 _047_
rlabel metal3 27412 17528 27412 17528 0 _048_
rlabel metal2 23016 18480 23016 18480 0 _049_
rlabel metal2 22792 18816 22792 18816 0 _050_
rlabel metal2 20888 20328 20888 20328 0 _051_
rlabel metal2 22456 18032 22456 18032 0 _052_
rlabel metal2 22792 16744 22792 16744 0 _053_
rlabel metal2 26936 15232 26936 15232 0 _054_
rlabel metal2 27160 15792 27160 15792 0 _055_
rlabel metal3 27328 17304 27328 17304 0 _056_
rlabel metal2 27272 16688 27272 16688 0 _057_
rlabel metal3 26908 21560 26908 21560 0 _058_
rlabel metal3 26824 18536 26824 18536 0 _059_
rlabel metal2 22064 26936 22064 26936 0 _060_
rlabel metal2 27272 14616 27272 14616 0 _061_
rlabel metal3 25256 15400 25256 15400 0 _062_
rlabel metal2 26544 15288 26544 15288 0 _063_
rlabel metal2 24808 14504 24808 14504 0 _064_
rlabel metal2 27720 23520 27720 23520 0 _065_
rlabel metal2 29736 22176 29736 22176 0 _066_
rlabel metal2 27832 24304 27832 24304 0 _067_
rlabel metal2 29008 24920 29008 24920 0 _068_
rlabel metal2 27496 24976 27496 24976 0 _069_
rlabel metal2 25928 22456 25928 22456 0 _070_
rlabel metal2 27272 24640 27272 24640 0 _071_
rlabel metal2 26824 24248 26824 24248 0 _072_
rlabel metal2 22680 25480 22680 25480 0 _073_
rlabel metal2 29064 20888 29064 20888 0 _074_
rlabel metal2 21448 20328 21448 20328 0 _075_
rlabel metal3 24192 20552 24192 20552 0 _076_
rlabel metal3 21560 22904 21560 22904 0 _077_
rlabel metal2 22568 23856 22568 23856 0 _078_
rlabel metal2 19432 26908 19432 26908 0 _079_
rlabel metal2 20104 26992 20104 26992 0 _080_
rlabel metal3 18536 22120 18536 22120 0 _081_
rlabel metal2 20664 22792 20664 22792 0 _082_
rlabel metal2 20104 19488 20104 19488 0 _083_
rlabel metal2 18312 18984 18312 18984 0 _084_
rlabel metal2 22008 20720 22008 20720 0 _085_
rlabel metal2 19264 20664 19264 20664 0 _086_
rlabel metal2 19600 23800 19600 23800 0 _087_
rlabel metal2 14504 22736 14504 22736 0 _088_
rlabel metal2 16296 21952 16296 21952 0 _089_
rlabel metal2 14672 22344 14672 22344 0 _090_
rlabel metal3 18144 19992 18144 19992 0 _091_
rlabel metal3 15736 17528 15736 17528 0 _092_
rlabel metal2 14280 22792 14280 22792 0 _093_
rlabel metal3 14000 23352 14000 23352 0 _094_
rlabel metal2 23800 17248 23800 17248 0 _095_
rlabel metal2 22456 18928 22456 18928 0 _096_
rlabel metal2 20664 19264 20664 19264 0 _097_
rlabel metal2 15064 23072 15064 23072 0 _098_
rlabel metal2 15064 24864 15064 24864 0 _099_
rlabel metal2 16800 20104 16800 20104 0 _100_
rlabel metal2 14728 21168 14728 21168 0 _101_
rlabel metal2 14840 23408 14840 23408 0 _102_
rlabel metal2 15288 25536 15288 25536 0 _103_
rlabel metal2 15904 21784 15904 21784 0 _104_
rlabel metal2 15512 25088 15512 25088 0 _105_
rlabel metal2 25592 18816 25592 18816 0 _106_
rlabel metal2 28056 18872 28056 18872 0 _107_
rlabel metal2 28168 24640 28168 24640 0 _108_
rlabel metal2 28504 24248 28504 24248 0 _109_
rlabel metal2 28728 19488 28728 19488 0 _110_
rlabel metal2 17808 18424 17808 18424 0 _111_
rlabel metal2 16408 17920 16408 17920 0 _112_
rlabel metal2 23352 21504 23352 21504 0 _113_
rlabel metal2 19880 16408 19880 16408 0 _114_
rlabel metal3 2478 27608 2478 27608 0 clk
rlabel metal2 23352 20440 23352 20440 0 clknet_0_clk
rlabel metal3 21168 14616 21168 14616 0 clknet_1_0__leaf_clk
rlabel metal2 28392 25088 28392 25088 0 clknet_1_1__leaf_clk
rlabel metal2 15736 20048 15736 20048 0 dut12.count\[0\]
rlabel metal2 16632 17584 16632 17584 0 dut12.count\[1\]
rlabel metal2 20440 14616 20440 14616 0 dut12.count\[2\]
rlabel metal2 21224 23296 21224 23296 0 dut12.count\[3\]
rlabel metal3 24528 26936 24528 26936 0 net1
rlabel metal2 12824 26208 12824 26208 0 net10
rlabel metal3 31920 21672 31920 21672 0 net11
rlabel metal3 28896 25368 28896 25368 0 net12
rlabel metal2 28616 14504 28616 14504 0 net13
rlabel metal2 27832 25536 27832 25536 0 net14
rlabel metal3 6356 18424 6356 18424 0 net15
rlabel metal2 30016 21784 30016 21784 0 net16
rlabel metal2 29176 24976 29176 24976 0 net17
rlabel metal3 6356 19992 6356 19992 0 net18
rlabel metal2 18760 27160 18760 27160 0 net19
rlabel metal2 24584 5964 24584 5964 0 net2
rlabel metal2 21448 5964 21448 5964 0 net20
rlabel metal3 31052 20104 31052 20104 0 net21
rlabel metal3 6356 23912 6356 23912 0 net22
rlabel metal3 27384 3528 27384 3528 0 net23
rlabel metal2 20328 27328 20328 27328 0 net24
rlabel metal2 23688 30212 23688 30212 0 net25
rlabel metal3 29512 20552 29512 20552 0 net26
rlabel metal3 23968 26152 23968 26152 0 net3
rlabel metal2 29960 17192 29960 17192 0 net4
rlabel metal2 30856 15624 30856 15624 0 net5
rlabel metal3 27776 13832 27776 13832 0 net6
rlabel metal2 4312 25368 4312 25368 0 net7
rlabel metal2 23464 28560 23464 28560 0 net8
rlabel metal2 25872 13048 25872 13048 0 net9
rlabel metal2 24248 39354 24248 39354 0 segm[0]
rlabel metal2 24248 2198 24248 2198 0 segm[10]
rlabel metal2 22904 39746 22904 39746 0 segm[11]
rlabel metal2 40040 17640 40040 17640 0 segm[12]
rlabel metal2 40040 16800 40040 16800 0 segm[13]
rlabel metal2 26936 2422 26936 2422 0 segm[1]
rlabel metal3 1414 24920 1414 24920 0 segm[2]
rlabel metal2 22232 39690 22232 39690 0 segm[3]
rlabel metal2 25592 2086 25592 2086 0 segm[4]
rlabel metal3 1358 25592 1358 25592 0 segm[5]
rlabel metal2 40040 21504 40040 21504 0 segm[6]
rlabel metal2 40040 26712 40040 26712 0 segm[7]
rlabel metal2 40040 14392 40040 14392 0 segm[8]
rlabel metal2 40040 25256 40040 25256 0 segm[9]
rlabel metal3 1358 18200 1358 18200 0 sel[0]
rlabel metal2 40040 22344 40040 22344 0 sel[10]
rlabel metal2 39928 25872 39928 25872 0 sel[11]
rlabel metal3 1358 19544 1358 19544 0 sel[1]
rlabel metal2 18872 39690 18872 39690 0 sel[2]
rlabel metal2 21560 2198 21560 2198 0 sel[3]
rlabel metal2 40040 19656 40040 19656 0 sel[4]
rlabel metal3 1358 23576 1358 23576 0 sel[5]
rlabel metal2 26264 2198 26264 2198 0 sel[6]
rlabel metal2 20216 39354 20216 39354 0 sel[7]
rlabel metal2 23576 38962 23576 38962 0 sel[8]
rlabel metal3 40642 20888 40642 20888 0 sel[9]
<< properties >>
string FIXED_BBOX 0 0 42000 42000
<< end >>
