magic
tech gf180mcuD
magscale 1 10
timestamp 1699642277
<< metal1 >>
rect 1344 38442 40656 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 40656 38442
rect 1344 38356 40656 38390
rect 19182 38274 19234 38286
rect 19182 38210 19234 38222
rect 22094 38274 22146 38286
rect 22094 38210 22146 38222
rect 25566 38274 25618 38286
rect 25566 38210 25618 38222
rect 19730 37998 19742 38050
rect 19794 37998 19806 38050
rect 21074 37998 21086 38050
rect 21138 37998 21150 38050
rect 24546 37998 24558 38050
rect 24610 37998 24622 38050
rect 1344 37658 40656 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 40656 37658
rect 1344 37572 40656 37606
rect 18398 37490 18450 37502
rect 18398 37426 18450 37438
rect 21422 37490 21474 37502
rect 21422 37426 21474 37438
rect 26238 37490 26290 37502
rect 26238 37426 26290 37438
rect 17714 37214 17726 37266
rect 17778 37214 17790 37266
rect 20514 37214 20526 37266
rect 20578 37214 20590 37266
rect 25218 37214 25230 37266
rect 25282 37214 25294 37266
rect 1344 36874 40656 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 40656 36874
rect 1344 36788 40656 36822
rect 17390 36706 17442 36718
rect 17390 36642 17442 36654
rect 16370 36430 16382 36482
rect 16434 36430 16446 36482
rect 1344 36090 40656 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 40656 36090
rect 1344 36004 40656 36038
rect 1344 35306 40656 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 40656 35306
rect 1344 35220 40656 35254
rect 1344 34522 40656 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 40656 34522
rect 1344 34436 40656 34470
rect 1344 33738 40656 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 40656 33738
rect 1344 33652 40656 33686
rect 1344 32954 40656 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 40656 32954
rect 1344 32868 40656 32902
rect 1344 32170 40656 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 40656 32170
rect 1344 32084 40656 32118
rect 1344 31386 40656 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 40656 31386
rect 1344 31300 40656 31334
rect 1344 30602 40656 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 40656 30602
rect 1344 30516 40656 30550
rect 1344 29818 40656 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 40656 29818
rect 1344 29732 40656 29766
rect 1344 29034 40656 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 40656 29034
rect 1344 28948 40656 28982
rect 1344 28250 40656 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 40656 28250
rect 1344 28164 40656 28198
rect 15934 28082 15986 28094
rect 15934 28018 15986 28030
rect 15710 27858 15762 27870
rect 15710 27794 15762 27806
rect 16046 27858 16098 27870
rect 17378 27806 17390 27858
rect 17442 27806 17454 27858
rect 21410 27806 21422 27858
rect 21474 27806 21486 27858
rect 37874 27806 37886 27858
rect 37938 27806 37950 27858
rect 16046 27794 16098 27806
rect 21198 27746 21250 27758
rect 18162 27694 18174 27746
rect 18226 27694 18238 27746
rect 20290 27694 20302 27746
rect 20354 27694 20366 27746
rect 22194 27694 22206 27746
rect 22258 27694 22270 27746
rect 24322 27694 24334 27746
rect 24386 27694 24398 27746
rect 21198 27682 21250 27694
rect 40014 27634 40066 27646
rect 40014 27570 40066 27582
rect 1344 27466 40656 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 40656 27466
rect 1344 27380 40656 27414
rect 23550 27298 23602 27310
rect 23550 27234 23602 27246
rect 40014 27186 40066 27198
rect 17266 27134 17278 27186
rect 17330 27134 17342 27186
rect 27570 27134 27582 27186
rect 27634 27134 27646 27186
rect 40014 27122 40066 27134
rect 17838 27074 17890 27086
rect 14466 27022 14478 27074
rect 14530 27022 14542 27074
rect 17838 27010 17890 27022
rect 18174 27074 18226 27086
rect 18174 27010 18226 27022
rect 19070 27074 19122 27086
rect 19070 27010 19122 27022
rect 22766 27074 22818 27086
rect 22766 27010 22818 27022
rect 23102 27074 23154 27086
rect 23102 27010 23154 27022
rect 23438 27074 23490 27086
rect 24546 27022 24558 27074
rect 24610 27022 24622 27074
rect 28130 27022 28142 27074
rect 28194 27022 28206 27074
rect 37650 27022 37662 27074
rect 37714 27022 37726 27074
rect 23438 27010 23490 27022
rect 17502 26962 17554 26974
rect 15138 26910 15150 26962
rect 15202 26910 15214 26962
rect 17502 26898 17554 26910
rect 17726 26962 17778 26974
rect 17726 26898 17778 26910
rect 18510 26962 18562 26974
rect 18510 26898 18562 26910
rect 18734 26962 18786 26974
rect 18734 26898 18786 26910
rect 18958 26962 19010 26974
rect 18958 26898 19010 26910
rect 23550 26962 23602 26974
rect 25330 26910 25342 26962
rect 25394 26910 25406 26962
rect 28354 26910 28366 26962
rect 28418 26910 28430 26962
rect 23550 26898 23602 26910
rect 18398 26850 18450 26862
rect 20526 26850 20578 26862
rect 20178 26798 20190 26850
rect 20242 26847 20254 26850
rect 20402 26847 20414 26850
rect 20242 26801 20414 26847
rect 20242 26798 20254 26801
rect 20402 26798 20414 26801
rect 20466 26798 20478 26850
rect 18398 26786 18450 26798
rect 20526 26786 20578 26798
rect 22990 26850 23042 26862
rect 22990 26786 23042 26798
rect 24222 26850 24274 26862
rect 24222 26786 24274 26798
rect 1344 26682 40656 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 40656 26682
rect 1344 26596 40656 26630
rect 16382 26514 16434 26526
rect 25902 26514 25954 26526
rect 20514 26462 20526 26514
rect 20578 26462 20590 26514
rect 23090 26462 23102 26514
rect 23154 26462 23166 26514
rect 16382 26450 16434 26462
rect 25902 26450 25954 26462
rect 16606 26402 16658 26414
rect 16606 26338 16658 26350
rect 16718 26402 16770 26414
rect 16718 26338 16770 26350
rect 25342 26402 25394 26414
rect 27122 26350 27134 26402
rect 27186 26350 27198 26402
rect 25342 26338 25394 26350
rect 25454 26290 25506 26302
rect 13346 26238 13358 26290
rect 13410 26238 13422 26290
rect 20290 26238 20302 26290
rect 20354 26238 20366 26290
rect 23314 26238 23326 26290
rect 23378 26238 23390 26290
rect 25454 26226 25506 26238
rect 25678 26290 25730 26302
rect 25678 26226 25730 26238
rect 26014 26290 26066 26302
rect 26898 26238 26910 26290
rect 26962 26238 26974 26290
rect 37650 26238 37662 26290
rect 37714 26238 37726 26290
rect 26014 26226 26066 26238
rect 17502 26178 17554 26190
rect 14018 26126 14030 26178
rect 14082 26126 14094 26178
rect 16146 26126 16158 26178
rect 16210 26126 16222 26178
rect 39890 26126 39902 26178
rect 39954 26126 39966 26178
rect 17502 26114 17554 26126
rect 25342 26066 25394 26078
rect 25342 26002 25394 26014
rect 1344 25898 40656 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 40656 25898
rect 1344 25812 40656 25846
rect 22878 25730 22930 25742
rect 22878 25666 22930 25678
rect 20738 25566 20750 25618
rect 20802 25566 20814 25618
rect 14926 25506 14978 25518
rect 14926 25442 14978 25454
rect 15262 25506 15314 25518
rect 17826 25454 17838 25506
rect 17890 25454 17902 25506
rect 15262 25442 15314 25454
rect 22766 25394 22818 25406
rect 18610 25342 18622 25394
rect 18674 25342 18686 25394
rect 22766 25330 22818 25342
rect 15150 25282 15202 25294
rect 15150 25218 15202 25230
rect 16382 25282 16434 25294
rect 16382 25218 16434 25230
rect 21422 25282 21474 25294
rect 21422 25218 21474 25230
rect 22878 25282 22930 25294
rect 22878 25218 22930 25230
rect 23886 25282 23938 25294
rect 23886 25218 23938 25230
rect 1344 25114 40656 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 40656 25114
rect 1344 25028 40656 25062
rect 19070 24946 19122 24958
rect 19070 24882 19122 24894
rect 19294 24946 19346 24958
rect 19294 24882 19346 24894
rect 19630 24946 19682 24958
rect 19630 24882 19682 24894
rect 19854 24946 19906 24958
rect 19854 24882 19906 24894
rect 24558 24946 24610 24958
rect 24558 24882 24610 24894
rect 24334 24834 24386 24846
rect 24334 24770 24386 24782
rect 19406 24722 19458 24734
rect 19406 24658 19458 24670
rect 19966 24722 20018 24734
rect 24222 24722 24274 24734
rect 20738 24670 20750 24722
rect 20802 24670 20814 24722
rect 19966 24658 20018 24670
rect 24222 24658 24274 24670
rect 21522 24558 21534 24610
rect 21586 24558 21598 24610
rect 23650 24558 23662 24610
rect 23714 24558 23726 24610
rect 1344 24330 40656 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 40656 24330
rect 1344 24244 40656 24278
rect 18286 24162 18338 24174
rect 18286 24098 18338 24110
rect 1934 24050 1986 24062
rect 19854 24050 19906 24062
rect 14578 23998 14590 24050
rect 14642 23998 14654 24050
rect 1934 23986 1986 23998
rect 19854 23986 19906 23998
rect 21870 24050 21922 24062
rect 21870 23986 21922 23998
rect 22990 24050 23042 24062
rect 22990 23986 23042 23998
rect 25230 24050 25282 24062
rect 40014 24050 40066 24062
rect 28466 23998 28478 24050
rect 28530 23998 28542 24050
rect 25230 23986 25282 23998
rect 40014 23986 40066 23998
rect 15262 23938 15314 23950
rect 4274 23886 4286 23938
rect 4338 23886 4350 23938
rect 15262 23874 15314 23886
rect 19630 23938 19682 23950
rect 19630 23874 19682 23886
rect 21646 23938 21698 23950
rect 21646 23874 21698 23886
rect 22094 23938 22146 23950
rect 22094 23874 22146 23886
rect 22654 23938 22706 23950
rect 22654 23874 22706 23886
rect 22878 23938 22930 23950
rect 22878 23874 22930 23886
rect 23438 23938 23490 23950
rect 23438 23874 23490 23886
rect 23662 23938 23714 23950
rect 23662 23874 23714 23886
rect 24110 23938 24162 23950
rect 24110 23874 24162 23886
rect 24446 23938 24498 23950
rect 25554 23886 25566 23938
rect 25618 23886 25630 23938
rect 37650 23886 37662 23938
rect 37714 23886 37726 23938
rect 24446 23874 24498 23886
rect 14702 23826 14754 23838
rect 14702 23762 14754 23774
rect 14926 23826 14978 23838
rect 14926 23762 14978 23774
rect 18174 23826 18226 23838
rect 18174 23762 18226 23774
rect 20078 23826 20130 23838
rect 20078 23762 20130 23774
rect 20302 23826 20354 23838
rect 23998 23826 24050 23838
rect 22306 23774 22318 23826
rect 22370 23774 22382 23826
rect 26338 23774 26350 23826
rect 26402 23774 26414 23826
rect 20302 23762 20354 23774
rect 23998 23762 24050 23774
rect 15374 23714 15426 23726
rect 15374 23650 15426 23662
rect 15822 23714 15874 23726
rect 15822 23650 15874 23662
rect 18286 23714 18338 23726
rect 18286 23650 18338 23662
rect 21534 23714 21586 23726
rect 21534 23650 21586 23662
rect 23886 23714 23938 23726
rect 23886 23650 23938 23662
rect 24558 23714 24610 23726
rect 24558 23650 24610 23662
rect 1344 23546 40656 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 40656 23546
rect 1344 23460 40656 23494
rect 15598 23378 15650 23390
rect 15598 23314 15650 23326
rect 25678 23378 25730 23390
rect 25678 23314 25730 23326
rect 16270 23266 16322 23278
rect 16270 23202 16322 23214
rect 16830 23266 16882 23278
rect 20178 23214 20190 23266
rect 20242 23214 20254 23266
rect 16830 23202 16882 23214
rect 15486 23154 15538 23166
rect 4274 23102 4286 23154
rect 4338 23102 4350 23154
rect 14914 23102 14926 23154
rect 14978 23102 14990 23154
rect 15250 23102 15262 23154
rect 15314 23102 15326 23154
rect 15486 23090 15538 23102
rect 15710 23154 15762 23166
rect 16494 23154 16546 23166
rect 15922 23102 15934 23154
rect 15986 23102 15998 23154
rect 24658 23102 24670 23154
rect 24722 23102 24734 23154
rect 26002 23102 26014 23154
rect 26066 23102 26078 23154
rect 37650 23102 37662 23154
rect 37714 23102 37726 23154
rect 15710 23090 15762 23102
rect 16494 23090 16546 23102
rect 16382 23042 16434 23054
rect 12002 22990 12014 23042
rect 12066 22990 12078 23042
rect 14130 22990 14142 23042
rect 14194 22990 14206 23042
rect 26786 22990 26798 23042
rect 26850 22990 26862 23042
rect 28914 22990 28926 23042
rect 28978 22990 28990 23042
rect 16382 22978 16434 22990
rect 1934 22930 1986 22942
rect 1934 22866 1986 22878
rect 40014 22930 40066 22942
rect 40014 22866 40066 22878
rect 1344 22762 40656 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 40656 22762
rect 1344 22676 40656 22710
rect 20638 22482 20690 22494
rect 20178 22430 20190 22482
rect 20242 22430 20254 22482
rect 20638 22418 20690 22430
rect 21422 22482 21474 22494
rect 40014 22482 40066 22494
rect 25330 22430 25342 22482
rect 25394 22430 25406 22482
rect 26226 22430 26238 22482
rect 26290 22430 26302 22482
rect 21422 22418 21474 22430
rect 40014 22418 40066 22430
rect 15486 22370 15538 22382
rect 13682 22318 13694 22370
rect 13746 22318 13758 22370
rect 15138 22318 15150 22370
rect 15202 22318 15214 22370
rect 15486 22306 15538 22318
rect 15598 22370 15650 22382
rect 25790 22370 25842 22382
rect 26910 22370 26962 22382
rect 17266 22318 17278 22370
rect 17330 22318 17342 22370
rect 21858 22318 21870 22370
rect 21922 22318 21934 22370
rect 22418 22318 22430 22370
rect 22482 22318 22494 22370
rect 26338 22318 26350 22370
rect 26402 22318 26414 22370
rect 15598 22306 15650 22318
rect 25790 22306 25842 22318
rect 26910 22306 26962 22318
rect 27470 22370 27522 22382
rect 27470 22306 27522 22318
rect 27806 22370 27858 22382
rect 37650 22318 37662 22370
rect 37714 22318 37726 22370
rect 27806 22306 27858 22318
rect 13918 22258 13970 22270
rect 13918 22194 13970 22206
rect 15374 22258 15426 22270
rect 27134 22258 27186 22270
rect 18050 22206 18062 22258
rect 18114 22206 18126 22258
rect 23202 22206 23214 22258
rect 23266 22206 23278 22258
rect 15374 22194 15426 22206
rect 27134 22194 27186 22206
rect 27246 22258 27298 22270
rect 27246 22194 27298 22206
rect 14702 22146 14754 22158
rect 25902 22146 25954 22158
rect 22082 22094 22094 22146
rect 22146 22094 22158 22146
rect 14702 22082 14754 22094
rect 25902 22082 25954 22094
rect 26126 22146 26178 22158
rect 26126 22082 26178 22094
rect 27694 22146 27746 22158
rect 27694 22082 27746 22094
rect 1344 21978 40656 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 40656 21978
rect 1344 21892 40656 21926
rect 14702 21810 14754 21822
rect 14702 21746 14754 21758
rect 15262 21810 15314 21822
rect 15262 21746 15314 21758
rect 15822 21810 15874 21822
rect 17614 21810 17666 21822
rect 16818 21758 16830 21810
rect 16882 21758 16894 21810
rect 15822 21746 15874 21758
rect 17614 21746 17666 21758
rect 18062 21810 18114 21822
rect 23326 21810 23378 21822
rect 20178 21758 20190 21810
rect 20242 21758 20254 21810
rect 18062 21746 18114 21758
rect 23326 21746 23378 21758
rect 25566 21810 25618 21822
rect 25566 21746 25618 21758
rect 15486 21698 15538 21710
rect 13458 21646 13470 21698
rect 13522 21646 13534 21698
rect 15486 21634 15538 21646
rect 16046 21698 16098 21710
rect 16046 21634 16098 21646
rect 17838 21698 17890 21710
rect 17838 21634 17890 21646
rect 18286 21698 18338 21710
rect 25230 21698 25282 21710
rect 21410 21646 21422 21698
rect 21474 21646 21486 21698
rect 18286 21634 18338 21646
rect 25230 21634 25282 21646
rect 25342 21698 25394 21710
rect 25342 21634 25394 21646
rect 15598 21586 15650 21598
rect 14242 21534 14254 21586
rect 14306 21534 14318 21586
rect 15598 21522 15650 21534
rect 16158 21586 16210 21598
rect 16158 21522 16210 21534
rect 16494 21586 16546 21598
rect 16494 21522 16546 21534
rect 17278 21586 17330 21598
rect 17278 21522 17330 21534
rect 18398 21586 18450 21598
rect 23438 21586 23490 21598
rect 20402 21534 20414 21586
rect 20466 21534 20478 21586
rect 21186 21534 21198 21586
rect 21250 21534 21262 21586
rect 18398 21522 18450 21534
rect 23438 21522 23490 21534
rect 23662 21586 23714 21598
rect 23662 21522 23714 21534
rect 23886 21586 23938 21598
rect 23886 21522 23938 21534
rect 23998 21586 24050 21598
rect 24322 21534 24334 21586
rect 24386 21534 24398 21586
rect 37874 21534 37886 21586
rect 37938 21534 37950 21586
rect 23998 21522 24050 21534
rect 17502 21474 17554 21486
rect 11330 21422 11342 21474
rect 11394 21422 11406 21474
rect 39890 21422 39902 21474
rect 39954 21422 39966 21474
rect 17502 21410 17554 21422
rect 1344 21194 40656 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 40656 21194
rect 1344 21108 40656 21142
rect 20414 21026 20466 21038
rect 20414 20962 20466 20974
rect 1934 20914 1986 20926
rect 13694 20914 13746 20926
rect 20526 20914 20578 20926
rect 9986 20862 9998 20914
rect 10050 20862 10062 20914
rect 14242 20862 14254 20914
rect 14306 20862 14318 20914
rect 1934 20850 1986 20862
rect 13694 20850 13746 20862
rect 20526 20850 20578 20862
rect 40014 20914 40066 20926
rect 40014 20850 40066 20862
rect 4274 20750 4286 20802
rect 4338 20750 4350 20802
rect 12114 20750 12126 20802
rect 12178 20750 12190 20802
rect 12898 20750 12910 20802
rect 12962 20750 12974 20802
rect 14802 20750 14814 20802
rect 14866 20750 14878 20802
rect 21298 20750 21310 20802
rect 21362 20750 21374 20802
rect 37650 20750 37662 20802
rect 37714 20750 37726 20802
rect 25106 20638 25118 20690
rect 25170 20638 25182 20690
rect 14254 20578 14306 20590
rect 14254 20514 14306 20526
rect 14366 20578 14418 20590
rect 14366 20514 14418 20526
rect 14590 20578 14642 20590
rect 14590 20514 14642 20526
rect 20190 20578 20242 20590
rect 20190 20514 20242 20526
rect 20638 20578 20690 20590
rect 20638 20514 20690 20526
rect 27022 20578 27074 20590
rect 27022 20514 27074 20526
rect 1344 20410 40656 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 40656 20410
rect 1344 20324 40656 20358
rect 14590 20242 14642 20254
rect 14590 20178 14642 20190
rect 15710 20242 15762 20254
rect 15710 20178 15762 20190
rect 15822 20242 15874 20254
rect 15822 20178 15874 20190
rect 18622 20242 18674 20254
rect 18622 20178 18674 20190
rect 21198 20242 21250 20254
rect 21198 20178 21250 20190
rect 13358 20130 13410 20142
rect 13358 20066 13410 20078
rect 13694 20130 13746 20142
rect 13694 20066 13746 20078
rect 14254 20130 14306 20142
rect 14254 20066 14306 20078
rect 14814 20130 14866 20142
rect 18510 20130 18562 20142
rect 16482 20078 16494 20130
rect 16546 20078 16558 20130
rect 14814 20066 14866 20078
rect 18510 20066 18562 20078
rect 19182 20130 19234 20142
rect 19182 20066 19234 20078
rect 19742 20130 19794 20142
rect 19742 20066 19794 20078
rect 21758 20130 21810 20142
rect 21758 20066 21810 20078
rect 23102 20130 23154 20142
rect 23102 20066 23154 20078
rect 23550 20130 23602 20142
rect 23874 20078 23886 20130
rect 23938 20078 23950 20130
rect 24658 20078 24670 20130
rect 24722 20078 24734 20130
rect 30146 20078 30158 20130
rect 30210 20078 30222 20130
rect 23550 20066 23602 20078
rect 13918 20018 13970 20030
rect 4274 19966 4286 20018
rect 4338 19966 4350 20018
rect 13918 19954 13970 19966
rect 14478 20018 14530 20030
rect 14478 19954 14530 19966
rect 14702 20018 14754 20030
rect 15486 20018 15538 20030
rect 19070 20018 19122 20030
rect 15250 19966 15262 20018
rect 15314 19966 15326 20018
rect 16706 19966 16718 20018
rect 16770 19966 16782 20018
rect 14702 19954 14754 19966
rect 15486 19954 15538 19966
rect 19070 19954 19122 19966
rect 19406 20018 19458 20030
rect 19406 19954 19458 19966
rect 20862 20018 20914 20030
rect 20862 19954 20914 19966
rect 24334 20018 24386 20030
rect 24334 19954 24386 19966
rect 25454 20018 25506 20030
rect 25454 19954 25506 19966
rect 26126 20018 26178 20030
rect 29822 20018 29874 20030
rect 26674 19966 26686 20018
rect 26738 19966 26750 20018
rect 26126 19954 26178 19966
rect 29822 19954 29874 19966
rect 13470 19906 13522 19918
rect 13470 19842 13522 19854
rect 15598 19906 15650 19918
rect 21870 19906 21922 19918
rect 21074 19854 21086 19906
rect 21138 19854 21150 19906
rect 15598 19842 15650 19854
rect 21870 19842 21922 19854
rect 25678 19906 25730 19918
rect 27346 19854 27358 19906
rect 27410 19854 27422 19906
rect 29474 19854 29486 19906
rect 29538 19854 29550 19906
rect 25678 19842 25730 19854
rect 1934 19794 1986 19806
rect 1934 19730 1986 19742
rect 18734 19794 18786 19806
rect 18734 19730 18786 19742
rect 19630 19794 19682 19806
rect 19630 19730 19682 19742
rect 22878 19794 22930 19806
rect 22878 19730 22930 19742
rect 23214 19794 23266 19806
rect 23214 19730 23266 19742
rect 26126 19794 26178 19806
rect 26126 19730 26178 19742
rect 26238 19794 26290 19806
rect 26238 19730 26290 19742
rect 1344 19626 40656 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 40656 19626
rect 1344 19540 40656 19574
rect 18174 19458 18226 19470
rect 18174 19394 18226 19406
rect 24222 19458 24274 19470
rect 24222 19394 24274 19406
rect 26574 19458 26626 19470
rect 26574 19394 26626 19406
rect 19742 19346 19794 19358
rect 9986 19294 9998 19346
rect 10050 19294 10062 19346
rect 12114 19294 12126 19346
rect 12178 19294 12190 19346
rect 19742 19282 19794 19294
rect 13582 19234 13634 19246
rect 12898 19182 12910 19234
rect 12962 19182 12974 19234
rect 13582 19170 13634 19182
rect 15150 19234 15202 19246
rect 15150 19170 15202 19182
rect 15486 19234 15538 19246
rect 15486 19170 15538 19182
rect 16158 19234 16210 19246
rect 16158 19170 16210 19182
rect 17950 19234 18002 19246
rect 19182 19234 19234 19246
rect 20526 19234 20578 19246
rect 24334 19234 24386 19246
rect 18498 19182 18510 19234
rect 18562 19182 18574 19234
rect 20290 19182 20302 19234
rect 20354 19182 20366 19234
rect 22530 19182 22542 19234
rect 22594 19182 22606 19234
rect 17950 19170 18002 19182
rect 19182 19170 19234 19182
rect 20526 19170 20578 19182
rect 24334 19170 24386 19182
rect 26462 19234 26514 19246
rect 26462 19170 26514 19182
rect 17614 19122 17666 19134
rect 15810 19070 15822 19122
rect 15874 19070 15886 19122
rect 16482 19070 16494 19122
rect 16546 19070 16558 19122
rect 17614 19058 17666 19070
rect 19406 19122 19458 19134
rect 24222 19122 24274 19134
rect 21970 19070 21982 19122
rect 22034 19070 22046 19122
rect 22306 19070 22318 19122
rect 22370 19070 22382 19122
rect 19406 19058 19458 19070
rect 24222 19058 24274 19070
rect 26574 19122 26626 19134
rect 26574 19058 26626 19070
rect 15374 19010 15426 19022
rect 15374 18946 15426 18958
rect 16830 19010 16882 19022
rect 16830 18946 16882 18958
rect 17726 19010 17778 19022
rect 17726 18946 17778 18958
rect 18286 19010 18338 19022
rect 18286 18946 18338 18958
rect 18958 19010 19010 19022
rect 18958 18946 19010 18958
rect 19294 19010 19346 19022
rect 19294 18946 19346 18958
rect 21646 19010 21698 19022
rect 21646 18946 21698 18958
rect 1344 18842 40656 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 40656 18842
rect 1344 18756 40656 18790
rect 18398 18674 18450 18686
rect 18398 18610 18450 18622
rect 19070 18674 19122 18686
rect 19070 18610 19122 18622
rect 26574 18674 26626 18686
rect 26574 18610 26626 18622
rect 18174 18562 18226 18574
rect 23886 18562 23938 18574
rect 15474 18510 15486 18562
rect 15538 18510 15550 18562
rect 22306 18510 22318 18562
rect 22370 18510 22382 18562
rect 23426 18510 23438 18562
rect 23490 18510 23502 18562
rect 18174 18498 18226 18510
rect 23886 18498 23938 18510
rect 25790 18562 25842 18574
rect 25790 18498 25842 18510
rect 14814 18450 14866 18462
rect 14130 18398 14142 18450
rect 14194 18398 14206 18450
rect 14814 18386 14866 18398
rect 15038 18450 15090 18462
rect 15038 18386 15090 18398
rect 15822 18450 15874 18462
rect 15822 18386 15874 18398
rect 18846 18450 18898 18462
rect 18846 18386 18898 18398
rect 20638 18450 20690 18462
rect 21982 18450 22034 18462
rect 20962 18398 20974 18450
rect 21026 18398 21038 18450
rect 20638 18386 20690 18398
rect 21982 18386 22034 18398
rect 23102 18450 23154 18462
rect 23102 18386 23154 18398
rect 23774 18450 23826 18462
rect 23774 18386 23826 18398
rect 26126 18450 26178 18462
rect 26338 18398 26350 18450
rect 26402 18398 26414 18450
rect 26898 18398 26910 18450
rect 26962 18398 26974 18450
rect 37650 18398 37662 18450
rect 37714 18398 37726 18450
rect 26126 18386 26178 18398
rect 14478 18338 14530 18350
rect 14242 18286 14254 18338
rect 14306 18286 14318 18338
rect 14478 18274 14530 18286
rect 14926 18338 14978 18350
rect 14926 18274 14978 18286
rect 18286 18338 18338 18350
rect 18286 18274 18338 18286
rect 19630 18338 19682 18350
rect 19630 18274 19682 18286
rect 20526 18338 20578 18350
rect 20526 18274 20578 18286
rect 25454 18338 25506 18350
rect 27682 18286 27694 18338
rect 27746 18286 27758 18338
rect 29810 18286 29822 18338
rect 29874 18286 29886 18338
rect 25454 18274 25506 18286
rect 15262 18226 15314 18238
rect 15262 18162 15314 18174
rect 23886 18226 23938 18238
rect 40014 18226 40066 18238
rect 26338 18174 26350 18226
rect 26402 18174 26414 18226
rect 23886 18162 23938 18174
rect 40014 18162 40066 18174
rect 1344 18058 40656 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 40656 18058
rect 1344 17972 40656 18006
rect 14926 17890 14978 17902
rect 28142 17890 28194 17902
rect 27234 17838 27246 17890
rect 27298 17838 27310 17890
rect 14926 17826 14978 17838
rect 28142 17826 28194 17838
rect 1934 17778 1986 17790
rect 1934 17714 1986 17726
rect 20750 17778 20802 17790
rect 20750 17714 20802 17726
rect 27694 17778 27746 17790
rect 27694 17714 27746 17726
rect 28254 17778 28306 17790
rect 28254 17714 28306 17726
rect 29262 17778 29314 17790
rect 29262 17714 29314 17726
rect 40014 17778 40066 17790
rect 40014 17714 40066 17726
rect 15150 17666 15202 17678
rect 4274 17614 4286 17666
rect 4338 17614 4350 17666
rect 15150 17602 15202 17614
rect 15710 17666 15762 17678
rect 15710 17602 15762 17614
rect 16046 17666 16098 17678
rect 16046 17602 16098 17614
rect 18846 17666 18898 17678
rect 18846 17602 18898 17614
rect 19854 17666 19906 17678
rect 19854 17602 19906 17614
rect 20526 17666 20578 17678
rect 27806 17666 27858 17678
rect 25218 17614 25230 17666
rect 25282 17614 25294 17666
rect 27122 17614 27134 17666
rect 27186 17614 27198 17666
rect 28466 17614 28478 17666
rect 28530 17614 28542 17666
rect 37650 17614 37662 17666
rect 37714 17614 37726 17666
rect 20526 17602 20578 17614
rect 27806 17602 27858 17614
rect 15934 17554 15986 17566
rect 29150 17554 29202 17566
rect 18050 17502 18062 17554
rect 18114 17502 18126 17554
rect 22978 17502 22990 17554
rect 23042 17502 23054 17554
rect 27570 17502 27582 17554
rect 27634 17502 27646 17554
rect 15934 17490 15986 17502
rect 29150 17490 29202 17502
rect 18398 17442 18450 17454
rect 14578 17390 14590 17442
rect 14642 17390 14654 17442
rect 18398 17378 18450 17390
rect 18734 17442 18786 17454
rect 19506 17390 19518 17442
rect 19570 17390 19582 17442
rect 20178 17390 20190 17442
rect 20242 17390 20254 17442
rect 18734 17378 18786 17390
rect 1344 17274 40656 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 40656 17274
rect 1344 17188 40656 17222
rect 14814 17106 14866 17118
rect 23550 17106 23602 17118
rect 19506 17054 19518 17106
rect 19570 17054 19582 17106
rect 14814 17042 14866 17054
rect 23550 17042 23602 17054
rect 23774 17106 23826 17118
rect 23774 17042 23826 17054
rect 25566 17106 25618 17118
rect 25566 17042 25618 17054
rect 16046 16994 16098 17006
rect 16046 16930 16098 16942
rect 17502 16994 17554 17006
rect 17502 16930 17554 16942
rect 17614 16994 17666 17006
rect 17614 16930 17666 16942
rect 18622 16994 18674 17006
rect 18622 16930 18674 16942
rect 20638 16994 20690 17006
rect 20638 16930 20690 16942
rect 23438 16994 23490 17006
rect 23438 16930 23490 16942
rect 25790 16994 25842 17006
rect 27010 16942 27022 16994
rect 27074 16942 27086 16994
rect 25790 16930 25842 16942
rect 17278 16882 17330 16894
rect 20190 16882 20242 16894
rect 14354 16830 14366 16882
rect 14418 16830 14430 16882
rect 16594 16830 16606 16882
rect 16658 16830 16670 16882
rect 18050 16830 18062 16882
rect 18114 16830 18126 16882
rect 25218 16830 25230 16882
rect 25282 16830 25294 16882
rect 26338 16830 26350 16882
rect 26402 16830 26414 16882
rect 37650 16830 37662 16882
rect 37714 16830 37726 16882
rect 17278 16818 17330 16830
rect 20190 16818 20242 16830
rect 16270 16770 16322 16782
rect 11442 16718 11454 16770
rect 11506 16718 11518 16770
rect 13570 16718 13582 16770
rect 13634 16718 13646 16770
rect 16270 16706 16322 16718
rect 25678 16770 25730 16782
rect 40014 16770 40066 16782
rect 29138 16718 29150 16770
rect 29202 16718 29214 16770
rect 25678 16706 25730 16718
rect 40014 16706 40066 16718
rect 1344 16490 40656 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 40656 16490
rect 1344 16404 40656 16438
rect 21310 16210 21362 16222
rect 17266 16158 17278 16210
rect 17330 16158 17342 16210
rect 23762 16158 23774 16210
rect 23826 16158 23838 16210
rect 25890 16158 25902 16210
rect 25954 16158 25966 16210
rect 21310 16146 21362 16158
rect 13806 16098 13858 16110
rect 13806 16034 13858 16046
rect 15822 16098 15874 16110
rect 16718 16098 16770 16110
rect 16258 16046 16270 16098
rect 16322 16046 16334 16098
rect 17602 16046 17614 16098
rect 17666 16046 17678 16098
rect 18834 16046 18846 16098
rect 18898 16046 18910 16098
rect 19842 16046 19854 16098
rect 19906 16046 19918 16098
rect 20738 16046 20750 16098
rect 20802 16046 20814 16098
rect 21746 16046 21758 16098
rect 21810 16046 21822 16098
rect 22978 16046 22990 16098
rect 23042 16046 23054 16098
rect 15822 16034 15874 16046
rect 16718 16034 16770 16046
rect 13470 15986 13522 15998
rect 17154 15934 17166 15986
rect 17218 15934 17230 15986
rect 20402 15934 20414 15986
rect 20466 15934 20478 15986
rect 13470 15922 13522 15934
rect 15486 15874 15538 15886
rect 15486 15810 15538 15822
rect 15710 15874 15762 15886
rect 15710 15810 15762 15822
rect 26350 15874 26402 15886
rect 26350 15810 26402 15822
rect 26798 15874 26850 15886
rect 26798 15810 26850 15822
rect 1344 15706 40656 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 40656 15706
rect 1344 15620 40656 15654
rect 17390 15538 17442 15550
rect 17390 15474 17442 15486
rect 19070 15538 19122 15550
rect 19070 15474 19122 15486
rect 20638 15538 20690 15550
rect 25666 15486 25678 15538
rect 25730 15486 25742 15538
rect 20638 15474 20690 15486
rect 22878 15426 22930 15438
rect 14354 15374 14366 15426
rect 14418 15374 14430 15426
rect 22878 15362 22930 15374
rect 26014 15426 26066 15438
rect 26014 15362 26066 15374
rect 17950 15314 18002 15326
rect 19742 15314 19794 15326
rect 13682 15262 13694 15314
rect 13746 15262 13758 15314
rect 18498 15262 18510 15314
rect 18562 15262 18574 15314
rect 18834 15262 18846 15314
rect 18898 15262 18910 15314
rect 17950 15250 18002 15262
rect 19742 15250 19794 15262
rect 20190 15314 20242 15326
rect 22094 15314 22146 15326
rect 21634 15262 21646 15314
rect 21698 15262 21710 15314
rect 20190 15250 20242 15262
rect 22094 15250 22146 15262
rect 22766 15314 22818 15326
rect 22766 15250 22818 15262
rect 23326 15314 23378 15326
rect 25218 15262 25230 15314
rect 25282 15262 25294 15314
rect 25778 15262 25790 15314
rect 25842 15262 25854 15314
rect 23326 15250 23378 15262
rect 23102 15202 23154 15214
rect 16482 15150 16494 15202
rect 16546 15150 16558 15202
rect 23102 15138 23154 15150
rect 19966 15090 20018 15102
rect 19966 15026 20018 15038
rect 25566 15090 25618 15102
rect 25566 15026 25618 15038
rect 1344 14922 40656 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 40656 14922
rect 1344 14836 40656 14870
rect 19854 14754 19906 14766
rect 19854 14690 19906 14702
rect 16718 14642 16770 14654
rect 16718 14578 16770 14590
rect 18846 14642 18898 14654
rect 24658 14590 24670 14642
rect 24722 14590 24734 14642
rect 25778 14590 25790 14642
rect 25842 14590 25854 14642
rect 27906 14590 27918 14642
rect 27970 14590 27982 14642
rect 18846 14578 18898 14590
rect 19394 14478 19406 14530
rect 19458 14478 19470 14530
rect 20178 14478 20190 14530
rect 20242 14478 20254 14530
rect 21858 14478 21870 14530
rect 21922 14478 21934 14530
rect 24994 14478 25006 14530
rect 25058 14478 25070 14530
rect 17950 14418 18002 14430
rect 17602 14366 17614 14418
rect 17666 14366 17678 14418
rect 19170 14366 19182 14418
rect 19234 14366 19246 14418
rect 22530 14366 22542 14418
rect 22594 14366 22606 14418
rect 17950 14354 18002 14366
rect 18286 14306 18338 14318
rect 18286 14242 18338 14254
rect 19966 14306 20018 14318
rect 19966 14242 20018 14254
rect 1344 14138 40656 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 40656 14138
rect 1344 14052 40656 14086
rect 22094 13970 22146 13982
rect 22094 13906 22146 13918
rect 23438 13970 23490 13982
rect 23438 13906 23490 13918
rect 24670 13970 24722 13982
rect 24670 13906 24722 13918
rect 25342 13970 25394 13982
rect 25342 13906 25394 13918
rect 26350 13970 26402 13982
rect 26350 13906 26402 13918
rect 23662 13858 23714 13870
rect 19506 13806 19518 13858
rect 19570 13806 19582 13858
rect 23662 13794 23714 13806
rect 23774 13858 23826 13870
rect 23774 13794 23826 13806
rect 18722 13694 18734 13746
rect 18786 13694 18798 13746
rect 26462 13634 26514 13646
rect 21634 13582 21646 13634
rect 21698 13582 21710 13634
rect 26462 13570 26514 13582
rect 1344 13354 40656 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 40656 13354
rect 1344 13268 40656 13302
rect 18734 13074 18786 13086
rect 16034 13022 16046 13074
rect 16098 13022 16110 13074
rect 18162 13022 18174 13074
rect 18226 13022 18238 13074
rect 18734 13010 18786 13022
rect 15362 12910 15374 12962
rect 15426 12910 15438 12962
rect 1344 12570 40656 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 40656 12570
rect 1344 12484 40656 12518
rect 1344 11786 40656 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 40656 11786
rect 1344 11700 40656 11734
rect 1344 11002 40656 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 40656 11002
rect 1344 10916 40656 10950
rect 1344 10218 40656 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 40656 10218
rect 1344 10132 40656 10166
rect 1344 9434 40656 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 40656 9434
rect 1344 9348 40656 9382
rect 1344 8650 40656 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 40656 8650
rect 1344 8564 40656 8598
rect 1344 7866 40656 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 40656 7866
rect 1344 7780 40656 7814
rect 1344 7082 40656 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 40656 7082
rect 1344 6996 40656 7030
rect 1344 6298 40656 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 40656 6298
rect 1344 6212 40656 6246
rect 1344 5514 40656 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 40656 5514
rect 1344 5428 40656 5462
rect 1344 4730 40656 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 40656 4730
rect 1344 4644 40656 4678
rect 27122 4286 27134 4338
rect 27186 4286 27198 4338
rect 28142 4114 28194 4126
rect 28142 4050 28194 4062
rect 1344 3946 40656 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 40656 3946
rect 1344 3860 40656 3894
rect 25566 3666 25618 3678
rect 25566 3602 25618 3614
rect 24546 3502 24558 3554
rect 24610 3502 24622 3554
rect 12350 3330 12402 3342
rect 12350 3266 12402 3278
rect 1344 3162 40656 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 40656 3162
rect 1344 3076 40656 3110
<< via1 >>
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 19182 38222 19234 38274
rect 22094 38222 22146 38274
rect 25566 38222 25618 38274
rect 19742 37998 19794 38050
rect 21086 37998 21138 38050
rect 24558 37998 24610 38050
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 18398 37438 18450 37490
rect 21422 37438 21474 37490
rect 26238 37438 26290 37490
rect 17726 37214 17778 37266
rect 20526 37214 20578 37266
rect 25230 37214 25282 37266
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 17390 36654 17442 36706
rect 16382 36430 16434 36482
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 15934 28030 15986 28082
rect 15710 27806 15762 27858
rect 16046 27806 16098 27858
rect 17390 27806 17442 27858
rect 21422 27806 21474 27858
rect 37886 27806 37938 27858
rect 18174 27694 18226 27746
rect 20302 27694 20354 27746
rect 21198 27694 21250 27746
rect 22206 27694 22258 27746
rect 24334 27694 24386 27746
rect 40014 27582 40066 27634
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 23550 27246 23602 27298
rect 17278 27134 17330 27186
rect 27582 27134 27634 27186
rect 40014 27134 40066 27186
rect 14478 27022 14530 27074
rect 17838 27022 17890 27074
rect 18174 27022 18226 27074
rect 19070 27022 19122 27074
rect 22766 27022 22818 27074
rect 23102 27022 23154 27074
rect 23438 27022 23490 27074
rect 24558 27022 24610 27074
rect 28142 27022 28194 27074
rect 37662 27022 37714 27074
rect 15150 26910 15202 26962
rect 17502 26910 17554 26962
rect 17726 26910 17778 26962
rect 18510 26910 18562 26962
rect 18734 26910 18786 26962
rect 18958 26910 19010 26962
rect 23550 26910 23602 26962
rect 25342 26910 25394 26962
rect 28366 26910 28418 26962
rect 18398 26798 18450 26850
rect 20190 26798 20242 26850
rect 20414 26798 20466 26850
rect 20526 26798 20578 26850
rect 22990 26798 23042 26850
rect 24222 26798 24274 26850
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 16382 26462 16434 26514
rect 20526 26462 20578 26514
rect 23102 26462 23154 26514
rect 25902 26462 25954 26514
rect 16606 26350 16658 26402
rect 16718 26350 16770 26402
rect 25342 26350 25394 26402
rect 27134 26350 27186 26402
rect 13358 26238 13410 26290
rect 20302 26238 20354 26290
rect 23326 26238 23378 26290
rect 25454 26238 25506 26290
rect 25678 26238 25730 26290
rect 26014 26238 26066 26290
rect 26910 26238 26962 26290
rect 37662 26238 37714 26290
rect 14030 26126 14082 26178
rect 16158 26126 16210 26178
rect 17502 26126 17554 26178
rect 39902 26126 39954 26178
rect 25342 26014 25394 26066
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 22878 25678 22930 25730
rect 20750 25566 20802 25618
rect 14926 25454 14978 25506
rect 15262 25454 15314 25506
rect 17838 25454 17890 25506
rect 18622 25342 18674 25394
rect 22766 25342 22818 25394
rect 15150 25230 15202 25282
rect 16382 25230 16434 25282
rect 21422 25230 21474 25282
rect 22878 25230 22930 25282
rect 23886 25230 23938 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 19070 24894 19122 24946
rect 19294 24894 19346 24946
rect 19630 24894 19682 24946
rect 19854 24894 19906 24946
rect 24558 24894 24610 24946
rect 24334 24782 24386 24834
rect 19406 24670 19458 24722
rect 19966 24670 20018 24722
rect 20750 24670 20802 24722
rect 24222 24670 24274 24722
rect 21534 24558 21586 24610
rect 23662 24558 23714 24610
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 18286 24110 18338 24162
rect 1934 23998 1986 24050
rect 14590 23998 14642 24050
rect 19854 23998 19906 24050
rect 21870 23998 21922 24050
rect 22990 23998 23042 24050
rect 25230 23998 25282 24050
rect 28478 23998 28530 24050
rect 40014 23998 40066 24050
rect 4286 23886 4338 23938
rect 15262 23886 15314 23938
rect 19630 23886 19682 23938
rect 21646 23886 21698 23938
rect 22094 23886 22146 23938
rect 22654 23886 22706 23938
rect 22878 23886 22930 23938
rect 23438 23886 23490 23938
rect 23662 23886 23714 23938
rect 24110 23886 24162 23938
rect 24446 23886 24498 23938
rect 25566 23886 25618 23938
rect 37662 23886 37714 23938
rect 14702 23774 14754 23826
rect 14926 23774 14978 23826
rect 18174 23774 18226 23826
rect 20078 23774 20130 23826
rect 20302 23774 20354 23826
rect 22318 23774 22370 23826
rect 23998 23774 24050 23826
rect 26350 23774 26402 23826
rect 15374 23662 15426 23714
rect 15822 23662 15874 23714
rect 18286 23662 18338 23714
rect 21534 23662 21586 23714
rect 23886 23662 23938 23714
rect 24558 23662 24610 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 15598 23326 15650 23378
rect 25678 23326 25730 23378
rect 16270 23214 16322 23266
rect 16830 23214 16882 23266
rect 20190 23214 20242 23266
rect 4286 23102 4338 23154
rect 14926 23102 14978 23154
rect 15262 23102 15314 23154
rect 15486 23102 15538 23154
rect 15710 23102 15762 23154
rect 15934 23102 15986 23154
rect 16494 23102 16546 23154
rect 24670 23102 24722 23154
rect 26014 23102 26066 23154
rect 37662 23102 37714 23154
rect 12014 22990 12066 23042
rect 14142 22990 14194 23042
rect 16382 22990 16434 23042
rect 26798 22990 26850 23042
rect 28926 22990 28978 23042
rect 1934 22878 1986 22930
rect 40014 22878 40066 22930
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 20190 22430 20242 22482
rect 20638 22430 20690 22482
rect 21422 22430 21474 22482
rect 25342 22430 25394 22482
rect 26238 22430 26290 22482
rect 40014 22430 40066 22482
rect 13694 22318 13746 22370
rect 15150 22318 15202 22370
rect 15486 22318 15538 22370
rect 15598 22318 15650 22370
rect 17278 22318 17330 22370
rect 21870 22318 21922 22370
rect 22430 22318 22482 22370
rect 25790 22318 25842 22370
rect 26350 22318 26402 22370
rect 26910 22318 26962 22370
rect 27470 22318 27522 22370
rect 27806 22318 27858 22370
rect 37662 22318 37714 22370
rect 13918 22206 13970 22258
rect 15374 22206 15426 22258
rect 18062 22206 18114 22258
rect 23214 22206 23266 22258
rect 27134 22206 27186 22258
rect 27246 22206 27298 22258
rect 14702 22094 14754 22146
rect 22094 22094 22146 22146
rect 25902 22094 25954 22146
rect 26126 22094 26178 22146
rect 27694 22094 27746 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 14702 21758 14754 21810
rect 15262 21758 15314 21810
rect 15822 21758 15874 21810
rect 16830 21758 16882 21810
rect 17614 21758 17666 21810
rect 18062 21758 18114 21810
rect 20190 21758 20242 21810
rect 23326 21758 23378 21810
rect 25566 21758 25618 21810
rect 13470 21646 13522 21698
rect 15486 21646 15538 21698
rect 16046 21646 16098 21698
rect 17838 21646 17890 21698
rect 18286 21646 18338 21698
rect 21422 21646 21474 21698
rect 25230 21646 25282 21698
rect 25342 21646 25394 21698
rect 14254 21534 14306 21586
rect 15598 21534 15650 21586
rect 16158 21534 16210 21586
rect 16494 21534 16546 21586
rect 17278 21534 17330 21586
rect 18398 21534 18450 21586
rect 20414 21534 20466 21586
rect 21198 21534 21250 21586
rect 23438 21534 23490 21586
rect 23662 21534 23714 21586
rect 23886 21534 23938 21586
rect 23998 21534 24050 21586
rect 24334 21534 24386 21586
rect 37886 21534 37938 21586
rect 11342 21422 11394 21474
rect 17502 21422 17554 21474
rect 39902 21422 39954 21474
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 20414 20974 20466 21026
rect 1934 20862 1986 20914
rect 9998 20862 10050 20914
rect 13694 20862 13746 20914
rect 14254 20862 14306 20914
rect 20526 20862 20578 20914
rect 40014 20862 40066 20914
rect 4286 20750 4338 20802
rect 12126 20750 12178 20802
rect 12910 20750 12962 20802
rect 14814 20750 14866 20802
rect 21310 20750 21362 20802
rect 37662 20750 37714 20802
rect 25118 20638 25170 20690
rect 14254 20526 14306 20578
rect 14366 20526 14418 20578
rect 14590 20526 14642 20578
rect 20190 20526 20242 20578
rect 20638 20526 20690 20578
rect 27022 20526 27074 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 14590 20190 14642 20242
rect 15710 20190 15762 20242
rect 15822 20190 15874 20242
rect 18622 20190 18674 20242
rect 21198 20190 21250 20242
rect 13358 20078 13410 20130
rect 13694 20078 13746 20130
rect 14254 20078 14306 20130
rect 14814 20078 14866 20130
rect 16494 20078 16546 20130
rect 18510 20078 18562 20130
rect 19182 20078 19234 20130
rect 19742 20078 19794 20130
rect 21758 20078 21810 20130
rect 23102 20078 23154 20130
rect 23550 20078 23602 20130
rect 23886 20078 23938 20130
rect 24670 20078 24722 20130
rect 30158 20078 30210 20130
rect 4286 19966 4338 20018
rect 13918 19966 13970 20018
rect 14478 19966 14530 20018
rect 14702 19966 14754 20018
rect 15262 19966 15314 20018
rect 15486 19966 15538 20018
rect 16718 19966 16770 20018
rect 19070 19966 19122 20018
rect 19406 19966 19458 20018
rect 20862 19966 20914 20018
rect 24334 19966 24386 20018
rect 25454 19966 25506 20018
rect 26126 19966 26178 20018
rect 26686 19966 26738 20018
rect 29822 19966 29874 20018
rect 13470 19854 13522 19906
rect 15598 19854 15650 19906
rect 21086 19854 21138 19906
rect 21870 19854 21922 19906
rect 25678 19854 25730 19906
rect 27358 19854 27410 19906
rect 29486 19854 29538 19906
rect 1934 19742 1986 19794
rect 18734 19742 18786 19794
rect 19630 19742 19682 19794
rect 22878 19742 22930 19794
rect 23214 19742 23266 19794
rect 26126 19742 26178 19794
rect 26238 19742 26290 19794
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 18174 19406 18226 19458
rect 24222 19406 24274 19458
rect 26574 19406 26626 19458
rect 9998 19294 10050 19346
rect 12126 19294 12178 19346
rect 19742 19294 19794 19346
rect 12910 19182 12962 19234
rect 13582 19182 13634 19234
rect 15150 19182 15202 19234
rect 15486 19182 15538 19234
rect 16158 19182 16210 19234
rect 17950 19182 18002 19234
rect 18510 19182 18562 19234
rect 19182 19182 19234 19234
rect 20302 19182 20354 19234
rect 20526 19182 20578 19234
rect 22542 19182 22594 19234
rect 24334 19182 24386 19234
rect 26462 19182 26514 19234
rect 15822 19070 15874 19122
rect 16494 19070 16546 19122
rect 17614 19070 17666 19122
rect 19406 19070 19458 19122
rect 21982 19070 22034 19122
rect 22318 19070 22370 19122
rect 24222 19070 24274 19122
rect 26574 19070 26626 19122
rect 15374 18958 15426 19010
rect 16830 18958 16882 19010
rect 17726 18958 17778 19010
rect 18286 18958 18338 19010
rect 18958 18958 19010 19010
rect 19294 18958 19346 19010
rect 21646 18958 21698 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 18398 18622 18450 18674
rect 19070 18622 19122 18674
rect 26574 18622 26626 18674
rect 15486 18510 15538 18562
rect 18174 18510 18226 18562
rect 22318 18510 22370 18562
rect 23438 18510 23490 18562
rect 23886 18510 23938 18562
rect 25790 18510 25842 18562
rect 14142 18398 14194 18450
rect 14814 18398 14866 18450
rect 15038 18398 15090 18450
rect 15822 18398 15874 18450
rect 18846 18398 18898 18450
rect 20638 18398 20690 18450
rect 20974 18398 21026 18450
rect 21982 18398 22034 18450
rect 23102 18398 23154 18450
rect 23774 18398 23826 18450
rect 26126 18398 26178 18450
rect 26350 18398 26402 18450
rect 26910 18398 26962 18450
rect 37662 18398 37714 18450
rect 14254 18286 14306 18338
rect 14478 18286 14530 18338
rect 14926 18286 14978 18338
rect 18286 18286 18338 18338
rect 19630 18286 19682 18338
rect 20526 18286 20578 18338
rect 25454 18286 25506 18338
rect 27694 18286 27746 18338
rect 29822 18286 29874 18338
rect 15262 18174 15314 18226
rect 23886 18174 23938 18226
rect 26350 18174 26402 18226
rect 40014 18174 40066 18226
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 14926 17838 14978 17890
rect 27246 17838 27298 17890
rect 28142 17838 28194 17890
rect 1934 17726 1986 17778
rect 20750 17726 20802 17778
rect 27694 17726 27746 17778
rect 28254 17726 28306 17778
rect 29262 17726 29314 17778
rect 40014 17726 40066 17778
rect 4286 17614 4338 17666
rect 15150 17614 15202 17666
rect 15710 17614 15762 17666
rect 16046 17614 16098 17666
rect 18846 17614 18898 17666
rect 19854 17614 19906 17666
rect 20526 17614 20578 17666
rect 25230 17614 25282 17666
rect 27134 17614 27186 17666
rect 27806 17614 27858 17666
rect 28478 17614 28530 17666
rect 37662 17614 37714 17666
rect 15934 17502 15986 17554
rect 18062 17502 18114 17554
rect 22990 17502 23042 17554
rect 27582 17502 27634 17554
rect 29150 17502 29202 17554
rect 14590 17390 14642 17442
rect 18398 17390 18450 17442
rect 18734 17390 18786 17442
rect 19518 17390 19570 17442
rect 20190 17390 20242 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 14814 17054 14866 17106
rect 19518 17054 19570 17106
rect 23550 17054 23602 17106
rect 23774 17054 23826 17106
rect 25566 17054 25618 17106
rect 16046 16942 16098 16994
rect 17502 16942 17554 16994
rect 17614 16942 17666 16994
rect 18622 16942 18674 16994
rect 20638 16942 20690 16994
rect 23438 16942 23490 16994
rect 25790 16942 25842 16994
rect 27022 16942 27074 16994
rect 14366 16830 14418 16882
rect 16606 16830 16658 16882
rect 17278 16830 17330 16882
rect 18062 16830 18114 16882
rect 20190 16830 20242 16882
rect 25230 16830 25282 16882
rect 26350 16830 26402 16882
rect 37662 16830 37714 16882
rect 11454 16718 11506 16770
rect 13582 16718 13634 16770
rect 16270 16718 16322 16770
rect 25678 16718 25730 16770
rect 29150 16718 29202 16770
rect 40014 16718 40066 16770
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 17278 16158 17330 16210
rect 21310 16158 21362 16210
rect 23774 16158 23826 16210
rect 25902 16158 25954 16210
rect 13806 16046 13858 16098
rect 15822 16046 15874 16098
rect 16270 16046 16322 16098
rect 16718 16046 16770 16098
rect 17614 16046 17666 16098
rect 18846 16046 18898 16098
rect 19854 16046 19906 16098
rect 20750 16046 20802 16098
rect 21758 16046 21810 16098
rect 22990 16046 23042 16098
rect 13470 15934 13522 15986
rect 17166 15934 17218 15986
rect 20414 15934 20466 15986
rect 15486 15822 15538 15874
rect 15710 15822 15762 15874
rect 26350 15822 26402 15874
rect 26798 15822 26850 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 17390 15486 17442 15538
rect 19070 15486 19122 15538
rect 20638 15486 20690 15538
rect 25678 15486 25730 15538
rect 14366 15374 14418 15426
rect 22878 15374 22930 15426
rect 26014 15374 26066 15426
rect 13694 15262 13746 15314
rect 17950 15262 18002 15314
rect 18510 15262 18562 15314
rect 18846 15262 18898 15314
rect 19742 15262 19794 15314
rect 20190 15262 20242 15314
rect 21646 15262 21698 15314
rect 22094 15262 22146 15314
rect 22766 15262 22818 15314
rect 23326 15262 23378 15314
rect 25230 15262 25282 15314
rect 25790 15262 25842 15314
rect 16494 15150 16546 15202
rect 23102 15150 23154 15202
rect 19966 15038 20018 15090
rect 25566 15038 25618 15090
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 19854 14702 19906 14754
rect 16718 14590 16770 14642
rect 18846 14590 18898 14642
rect 24670 14590 24722 14642
rect 25790 14590 25842 14642
rect 27918 14590 27970 14642
rect 19406 14478 19458 14530
rect 20190 14478 20242 14530
rect 21870 14478 21922 14530
rect 25006 14478 25058 14530
rect 17614 14366 17666 14418
rect 17950 14366 18002 14418
rect 19182 14366 19234 14418
rect 22542 14366 22594 14418
rect 18286 14254 18338 14306
rect 19966 14254 20018 14306
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 22094 13918 22146 13970
rect 23438 13918 23490 13970
rect 24670 13918 24722 13970
rect 25342 13918 25394 13970
rect 26350 13918 26402 13970
rect 19518 13806 19570 13858
rect 23662 13806 23714 13858
rect 23774 13806 23826 13858
rect 18734 13694 18786 13746
rect 21646 13582 21698 13634
rect 26462 13582 26514 13634
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 16046 13022 16098 13074
rect 18174 13022 18226 13074
rect 18734 13022 18786 13074
rect 15374 12910 15426 12962
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 27134 4286 27186 4338
rect 28142 4062 28194 4114
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 25566 3614 25618 3666
rect 24558 3502 24610 3554
rect 12350 3278 12402 3330
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
<< metal2 >>
rect 16128 41200 16240 42000
rect 16800 41200 16912 42000
rect 19488 41200 19600 42000
rect 20160 41200 20272 42000
rect 20832 41200 20944 42000
rect 23520 41200 23632 42000
rect 24192 41200 24304 42000
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 16156 36708 16212 41200
rect 16828 37492 16884 41200
rect 19180 38276 19236 38286
rect 19516 38276 19572 41200
rect 20188 38612 20244 41200
rect 20188 38546 20244 38556
rect 19180 38274 19572 38276
rect 19180 38222 19182 38274
rect 19234 38222 19572 38274
rect 19180 38220 19572 38222
rect 20860 38276 20916 41200
rect 19180 38210 19236 38220
rect 20860 38210 20916 38220
rect 21420 38612 21476 38622
rect 19740 38052 19796 38062
rect 21084 38052 21140 38062
rect 19292 38050 19796 38052
rect 19292 37998 19742 38050
rect 19794 37998 19796 38050
rect 19292 37996 19796 37998
rect 16828 37426 16884 37436
rect 18396 37492 18452 37502
rect 18396 37398 18452 37436
rect 17724 37266 17780 37278
rect 17724 37214 17726 37266
rect 17778 37214 17780 37266
rect 16156 36642 16212 36652
rect 17388 36708 17444 36718
rect 17388 36614 17444 36652
rect 16380 36482 16436 36494
rect 16380 36430 16382 36482
rect 16434 36430 16436 36482
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 16380 31948 16436 36430
rect 15932 31892 16436 31948
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 15932 28082 15988 31892
rect 15932 28030 15934 28082
rect 15986 28030 15988 28082
rect 15708 27860 15764 27870
rect 15260 27858 15764 27860
rect 15260 27806 15710 27858
rect 15762 27806 15764 27858
rect 15260 27804 15764 27806
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 14476 27074 14532 27086
rect 14476 27022 14478 27074
rect 14530 27022 14532 27074
rect 4172 26964 4228 26974
rect 1932 24050 1988 24062
rect 1932 23998 1934 24050
rect 1986 23998 1988 24050
rect 1932 23604 1988 23998
rect 1932 23538 1988 23548
rect 1932 22932 1988 22942
rect 1932 22838 1988 22876
rect 1932 20914 1988 20926
rect 1932 20862 1934 20914
rect 1986 20862 1988 20914
rect 1932 20244 1988 20862
rect 4172 20580 4228 26908
rect 13356 26292 13412 26302
rect 13356 26198 13412 26236
rect 14476 26292 14532 27022
rect 15148 26964 15204 26974
rect 15148 26870 15204 26908
rect 14028 26178 14084 26190
rect 14028 26126 14030 26178
rect 14082 26126 14084 26178
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 14028 25732 14084 26126
rect 14028 25666 14084 25676
rect 14476 25284 14532 26236
rect 14924 25732 14980 25742
rect 14924 25506 14980 25676
rect 14924 25454 14926 25506
rect 14978 25454 14980 25506
rect 14924 25442 14980 25454
rect 15260 25506 15316 27804
rect 15708 27794 15764 27804
rect 15932 26180 15988 28030
rect 16044 27860 16100 27870
rect 16044 27766 16100 27804
rect 17388 27858 17444 27870
rect 17388 27806 17390 27858
rect 17442 27806 17444 27858
rect 17388 27412 17444 27806
rect 17164 27356 17444 27412
rect 16156 26964 16212 26974
rect 16716 26964 16772 26974
rect 16212 26908 16436 26964
rect 16156 26898 16212 26908
rect 16380 26514 16436 26908
rect 16380 26462 16382 26514
rect 16434 26462 16436 26514
rect 16380 26450 16436 26462
rect 16604 26402 16660 26414
rect 16604 26350 16606 26402
rect 16658 26350 16660 26402
rect 16156 26180 16212 26190
rect 15932 26178 16212 26180
rect 15932 26126 16158 26178
rect 16210 26126 16212 26178
rect 15932 26124 16212 26126
rect 16156 26114 16212 26124
rect 15260 25454 15262 25506
rect 15314 25454 15316 25506
rect 15260 25442 15316 25454
rect 14476 25218 14532 25228
rect 15148 25284 15204 25294
rect 16380 25284 16436 25294
rect 15148 25282 15540 25284
rect 15148 25230 15150 25282
rect 15202 25230 15540 25282
rect 15148 25228 15540 25230
rect 15148 25218 15204 25228
rect 15148 25060 15204 25070
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 14588 24052 14644 24062
rect 13468 24050 14644 24052
rect 13468 23998 14590 24050
rect 14642 23998 14644 24050
rect 13468 23996 14644 23998
rect 4284 23940 4340 23950
rect 4284 23846 4340 23884
rect 12012 23940 12068 23950
rect 4284 23156 4340 23166
rect 4284 23062 4340 23100
rect 11340 23156 11396 23166
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 11340 21474 11396 23100
rect 12012 23042 12068 23884
rect 12012 22990 12014 23042
rect 12066 22990 12068 23042
rect 12012 22978 12068 22990
rect 13468 21698 13524 23996
rect 14588 23986 14644 23996
rect 14700 23828 14756 23838
rect 14700 23734 14756 23772
rect 14924 23828 14980 23838
rect 14924 23826 15092 23828
rect 14924 23774 14926 23826
rect 14978 23774 15092 23826
rect 14924 23772 15092 23774
rect 14924 23762 14980 23772
rect 14924 23492 14980 23502
rect 14924 23156 14980 23436
rect 15036 23380 15092 23772
rect 15148 23492 15204 25004
rect 15260 23940 15316 23950
rect 15260 23846 15316 23884
rect 15372 23716 15428 23726
rect 15372 23622 15428 23660
rect 15148 23426 15204 23436
rect 15484 23380 15540 25228
rect 16380 25190 16436 25228
rect 16268 24724 16324 24734
rect 15820 23714 15876 23726
rect 15820 23662 15822 23714
rect 15874 23662 15876 23714
rect 15820 23492 15876 23662
rect 15820 23426 15876 23436
rect 15036 23314 15092 23324
rect 15372 23324 15540 23380
rect 15596 23380 15652 23390
rect 14812 23154 14980 23156
rect 14812 23102 14926 23154
rect 14978 23102 14980 23154
rect 14812 23100 14980 23102
rect 14140 23044 14196 23054
rect 13916 23042 14196 23044
rect 13916 22990 14142 23042
rect 14194 22990 14196 23042
rect 13916 22988 14196 22990
rect 13692 22370 13748 22382
rect 13692 22318 13694 22370
rect 13746 22318 13748 22370
rect 13692 22036 13748 22318
rect 13916 22258 13972 22988
rect 14140 22978 14196 22988
rect 13916 22206 13918 22258
rect 13970 22206 13972 22258
rect 13916 22194 13972 22206
rect 14700 22146 14756 22158
rect 14700 22094 14702 22146
rect 14754 22094 14756 22146
rect 14700 22036 14756 22094
rect 13692 21980 14756 22036
rect 14700 21812 14756 21822
rect 14812 21812 14868 23100
rect 14924 23090 14980 23100
rect 15260 23156 15316 23166
rect 15260 23062 15316 23100
rect 15148 23044 15204 23054
rect 15148 22370 15204 22988
rect 15372 22932 15428 23324
rect 15596 23286 15652 23324
rect 15932 23268 15988 23278
rect 15484 23156 15540 23166
rect 15484 23062 15540 23100
rect 15708 23154 15764 23166
rect 15708 23102 15710 23154
rect 15762 23102 15764 23154
rect 15372 22876 15540 22932
rect 15484 22484 15540 22876
rect 15148 22318 15150 22370
rect 15202 22318 15204 22370
rect 15148 22306 15204 22318
rect 15260 22428 15540 22484
rect 13468 21646 13470 21698
rect 13522 21646 13524 21698
rect 13468 21634 13524 21646
rect 14252 21810 14868 21812
rect 14252 21758 14702 21810
rect 14754 21758 14868 21810
rect 14252 21756 14868 21758
rect 15148 22148 15204 22158
rect 14252 21588 14308 21756
rect 14700 21746 14756 21756
rect 11340 21422 11342 21474
rect 11394 21422 11396 21474
rect 11340 21410 11396 21422
rect 13692 21586 14308 21588
rect 13692 21534 14254 21586
rect 14306 21534 14308 21586
rect 13692 21532 14308 21534
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 9996 20914 10052 20926
rect 9996 20862 9998 20914
rect 10050 20862 10052 20914
rect 4284 20804 4340 20814
rect 4284 20710 4340 20748
rect 9996 20692 10052 20862
rect 12908 20916 12964 20926
rect 12124 20804 12180 20814
rect 12124 20710 12180 20748
rect 12908 20802 12964 20860
rect 13692 20916 13748 21532
rect 14252 21522 14308 21532
rect 15148 21028 15204 22092
rect 15260 21810 15316 22428
rect 15484 22370 15540 22428
rect 15484 22318 15486 22370
rect 15538 22318 15540 22370
rect 15484 22306 15540 22318
rect 15596 22370 15652 22382
rect 15596 22318 15598 22370
rect 15650 22318 15652 22370
rect 15372 22258 15428 22270
rect 15372 22206 15374 22258
rect 15426 22206 15428 22258
rect 15372 21924 15428 22206
rect 15596 22148 15652 22318
rect 15596 22082 15652 22092
rect 15708 22036 15764 23102
rect 15932 23154 15988 23212
rect 15932 23102 15934 23154
rect 15986 23102 15988 23154
rect 15932 23090 15988 23102
rect 16268 23266 16324 24668
rect 16268 23214 16270 23266
rect 16322 23214 16324 23266
rect 16268 23156 16324 23214
rect 16268 23090 16324 23100
rect 16492 23716 16548 23726
rect 16492 23154 16548 23660
rect 16604 23604 16660 26350
rect 16716 26402 16772 26908
rect 16716 26350 16718 26402
rect 16770 26350 16772 26402
rect 16716 26338 16772 26350
rect 17164 26180 17220 27356
rect 17276 27188 17332 27198
rect 17724 27188 17780 37214
rect 17276 27186 17780 27188
rect 17276 27134 17278 27186
rect 17330 27134 17780 27186
rect 17276 27132 17780 27134
rect 17276 27122 17332 27132
rect 17500 26964 17556 26974
rect 17500 26870 17556 26908
rect 17724 26962 17780 27132
rect 17836 27860 17892 27870
rect 17836 27076 17892 27804
rect 17836 26982 17892 27020
rect 18172 27746 18228 27758
rect 19292 27748 19348 37996
rect 19740 37986 19796 37996
rect 20188 38050 21140 38052
rect 20188 37998 21086 38050
rect 21138 37998 21140 38050
rect 20188 37996 21140 37998
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 18172 27694 18174 27746
rect 18226 27694 18228 27746
rect 18172 27074 18228 27694
rect 18172 27022 18174 27074
rect 18226 27022 18228 27074
rect 18172 27010 18228 27022
rect 18956 27692 19292 27748
rect 17724 26910 17726 26962
rect 17778 26910 17780 26962
rect 17724 26898 17780 26910
rect 18508 26964 18564 26974
rect 18732 26964 18788 26974
rect 18508 26962 18788 26964
rect 18508 26910 18510 26962
rect 18562 26910 18734 26962
rect 18786 26910 18788 26962
rect 18508 26908 18788 26910
rect 18508 26898 18564 26908
rect 18732 26898 18788 26908
rect 18956 26962 19012 27692
rect 19292 27682 19348 27692
rect 19068 27076 19124 27086
rect 19068 26982 19124 27020
rect 18956 26910 18958 26962
rect 19010 26910 19012 26962
rect 18956 26898 19012 26910
rect 18396 26852 18452 26862
rect 18284 26850 18452 26852
rect 18284 26798 18398 26850
rect 18450 26798 18452 26850
rect 18284 26796 18452 26798
rect 17500 26180 17556 26190
rect 17164 26178 17556 26180
rect 17164 26126 17502 26178
rect 17554 26126 17556 26178
rect 17164 26124 17556 26126
rect 17500 25508 17556 26124
rect 17836 25508 17892 25518
rect 17500 25506 17892 25508
rect 17500 25454 17838 25506
rect 17890 25454 17892 25506
rect 17500 25452 17892 25454
rect 17836 25284 17892 25452
rect 17836 25218 17892 25228
rect 18284 24162 18340 26796
rect 18396 26786 18452 26796
rect 20188 26850 20244 37996
rect 21084 37986 21140 37996
rect 21420 37490 21476 38556
rect 22092 38276 22148 38286
rect 22092 38182 22148 38220
rect 23548 38276 23604 41200
rect 23548 38210 23604 38220
rect 21420 37438 21422 37490
rect 21474 37438 21476 37490
rect 21420 37426 21476 37438
rect 24220 37492 24276 41200
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 25564 38276 25620 38286
rect 25564 38182 25620 38220
rect 24220 37426 24276 37436
rect 24556 38050 24612 38062
rect 24556 37998 24558 38050
rect 24610 37998 24612 38050
rect 20524 37266 20580 37278
rect 20524 37214 20526 37266
rect 20578 37214 20580 37266
rect 20300 27748 20356 27758
rect 20300 27654 20356 27692
rect 20524 27188 20580 37214
rect 24556 31948 24612 37998
rect 26236 37492 26292 37502
rect 26236 37398 26292 37436
rect 23772 31892 24612 31948
rect 25228 37266 25284 37278
rect 25228 37214 25230 37266
rect 25282 37214 25284 37266
rect 21420 27858 21476 27870
rect 21420 27806 21422 27858
rect 21474 27806 21476 27858
rect 20188 26798 20190 26850
rect 20242 26798 20244 26850
rect 20188 26786 20244 26798
rect 20300 27132 20580 27188
rect 21196 27748 21252 27758
rect 21420 27748 21476 27806
rect 21196 27746 21476 27748
rect 21196 27694 21198 27746
rect 21250 27694 21476 27746
rect 21196 27692 21476 27694
rect 22204 27748 22260 27758
rect 23660 27748 23716 27758
rect 22204 27746 22820 27748
rect 22204 27694 22206 27746
rect 22258 27694 22820 27746
rect 22204 27692 22820 27694
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 20300 26290 20356 27132
rect 21196 26908 21252 27692
rect 22204 27682 22260 27692
rect 22764 27074 22820 27692
rect 23548 27300 23604 27310
rect 22764 27022 22766 27074
rect 22818 27022 22820 27074
rect 22764 27010 22820 27022
rect 23100 27298 23604 27300
rect 23100 27246 23550 27298
rect 23602 27246 23604 27298
rect 23100 27244 23604 27246
rect 23100 27074 23156 27244
rect 23548 27234 23604 27244
rect 23436 27076 23492 27086
rect 23100 27022 23102 27074
rect 23154 27022 23156 27074
rect 23100 27010 23156 27022
rect 23212 27020 23436 27076
rect 20412 26850 20468 26862
rect 20412 26798 20414 26850
rect 20466 26798 20468 26850
rect 20412 26628 20468 26798
rect 20524 26852 20580 26862
rect 20636 26852 21252 26908
rect 22988 26852 23044 26862
rect 20524 26850 20692 26852
rect 20524 26798 20526 26850
rect 20578 26798 20692 26850
rect 20524 26796 20692 26798
rect 20524 26786 20580 26796
rect 20412 26572 20580 26628
rect 20524 26514 20580 26572
rect 20524 26462 20526 26514
rect 20578 26462 20580 26514
rect 20524 26450 20580 26462
rect 20300 26238 20302 26290
rect 20354 26238 20356 26290
rect 18620 25396 18676 25406
rect 18620 25394 19124 25396
rect 18620 25342 18622 25394
rect 18674 25342 19124 25394
rect 18620 25340 19124 25342
rect 18620 25330 18676 25340
rect 19068 24946 19124 25340
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 19068 24894 19070 24946
rect 19122 24894 19124 24946
rect 19068 24882 19124 24894
rect 19292 24948 19348 24958
rect 19628 24948 19684 24958
rect 19292 24946 19684 24948
rect 19292 24894 19294 24946
rect 19346 24894 19630 24946
rect 19682 24894 19684 24946
rect 19292 24892 19684 24894
rect 19292 24882 19348 24892
rect 19628 24882 19684 24892
rect 19852 24948 19908 24958
rect 19852 24854 19908 24892
rect 20300 24948 20356 26238
rect 20300 24882 20356 24892
rect 20636 25284 20692 26796
rect 22876 26850 23044 26852
rect 22876 26798 22990 26850
rect 23042 26798 23044 26850
rect 22876 26796 23044 26798
rect 22876 25730 22932 26796
rect 22988 26786 23044 26796
rect 23100 26516 23156 26526
rect 23212 26516 23268 27020
rect 23436 26982 23492 27020
rect 23548 26964 23604 26974
rect 23660 26964 23716 27692
rect 23548 26962 23716 26964
rect 23548 26910 23550 26962
rect 23602 26910 23716 26962
rect 23548 26908 23716 26910
rect 23548 26898 23604 26908
rect 23100 26514 23268 26516
rect 23100 26462 23102 26514
rect 23154 26462 23268 26514
rect 23100 26460 23268 26462
rect 23100 26450 23156 26460
rect 22876 25678 22878 25730
rect 22930 25678 22932 25730
rect 22876 25666 22932 25678
rect 23324 26292 23380 26302
rect 19404 24724 19460 24734
rect 19964 24724 20020 24734
rect 19404 24722 19796 24724
rect 19404 24670 19406 24722
rect 19458 24670 19796 24722
rect 19404 24668 19796 24670
rect 19404 24658 19460 24668
rect 18284 24110 18286 24162
rect 18338 24110 18340 24162
rect 18284 24098 18340 24110
rect 19740 24052 19796 24668
rect 20636 24724 20692 25228
rect 20748 25618 20804 25630
rect 20748 25566 20750 25618
rect 20802 25566 20804 25618
rect 20748 24948 20804 25566
rect 22764 25396 22820 25406
rect 22540 25394 22820 25396
rect 22540 25342 22766 25394
rect 22818 25342 22820 25394
rect 22540 25340 22820 25342
rect 21420 25284 21476 25294
rect 21420 25190 21476 25228
rect 20748 24882 20804 24892
rect 20748 24724 20804 24734
rect 20636 24722 20804 24724
rect 20636 24670 20750 24722
rect 20802 24670 20804 24722
rect 20636 24668 20804 24670
rect 19964 24630 20020 24668
rect 19852 24052 19908 24062
rect 19740 24050 19908 24052
rect 19740 23998 19854 24050
rect 19906 23998 19908 24050
rect 19740 23996 19908 23998
rect 19852 23986 19908 23996
rect 19628 23938 19684 23950
rect 19628 23886 19630 23938
rect 19682 23886 19684 23938
rect 16604 23538 16660 23548
rect 16828 23828 16884 23838
rect 16492 23102 16494 23154
rect 16546 23102 16548 23154
rect 16492 23090 16548 23102
rect 16604 23268 16660 23278
rect 16380 23044 16436 23054
rect 16380 22950 16436 22988
rect 15708 21980 15988 22036
rect 15372 21868 15876 21924
rect 15260 21758 15262 21810
rect 15314 21758 15316 21810
rect 15260 21746 15316 21758
rect 15820 21810 15876 21868
rect 15820 21758 15822 21810
rect 15874 21758 15876 21810
rect 15820 21746 15876 21758
rect 15932 21812 15988 21980
rect 15932 21746 15988 21756
rect 14812 20972 15204 21028
rect 13692 20822 13748 20860
rect 14252 20914 14308 20926
rect 14252 20862 14254 20914
rect 14306 20862 14308 20914
rect 12908 20750 12910 20802
rect 12962 20750 12964 20802
rect 12908 20738 12964 20750
rect 14252 20804 14308 20862
rect 14252 20738 14308 20748
rect 14812 20802 14868 20972
rect 14812 20750 14814 20802
rect 14866 20750 14868 20802
rect 14812 20738 14868 20750
rect 9996 20626 10052 20636
rect 14140 20692 14196 20702
rect 4172 20514 4228 20524
rect 13468 20244 13524 20254
rect 1932 20178 1988 20188
rect 13356 20132 13524 20188
rect 14140 20188 14196 20636
rect 14700 20692 14756 20702
rect 14252 20578 14308 20590
rect 14252 20526 14254 20578
rect 14306 20526 14308 20578
rect 14252 20356 14308 20526
rect 14252 20290 14308 20300
rect 14364 20578 14420 20590
rect 14364 20526 14366 20578
rect 14418 20526 14420 20578
rect 14364 20188 14420 20526
rect 14588 20578 14644 20590
rect 14588 20526 14590 20578
rect 14642 20526 14644 20578
rect 14476 20356 14532 20366
rect 14476 20188 14532 20300
rect 13692 20132 13748 20142
rect 14140 20132 14308 20188
rect 13356 20130 13412 20132
rect 13356 20078 13358 20130
rect 13410 20078 13412 20130
rect 13356 20066 13412 20078
rect 13692 20038 13748 20076
rect 14252 20130 14308 20132
rect 14252 20078 14254 20130
rect 14306 20078 14308 20130
rect 14252 20066 14308 20078
rect 14364 20132 14532 20188
rect 14588 20242 14644 20526
rect 14588 20190 14590 20242
rect 14642 20190 14644 20242
rect 14588 20178 14644 20190
rect 14364 20066 14420 20076
rect 4284 20020 4340 20030
rect 4284 19926 4340 19964
rect 13916 20020 13972 20030
rect 13916 19926 13972 19964
rect 14476 20018 14532 20030
rect 14476 19966 14478 20018
rect 14530 19966 14532 20018
rect 12124 19908 12180 19918
rect 1932 19796 1988 19806
rect 1932 19702 1988 19740
rect 9996 19796 10052 19806
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 9996 19346 10052 19740
rect 9996 19294 9998 19346
rect 10050 19294 10052 19346
rect 9996 19282 10052 19294
rect 12124 19346 12180 19852
rect 13468 19908 13524 19918
rect 13468 19814 13524 19852
rect 14476 19460 14532 19966
rect 14476 19394 14532 19404
rect 14700 20018 14756 20636
rect 14812 20132 14868 20142
rect 14812 20038 14868 20076
rect 14700 19966 14702 20018
rect 14754 19966 14756 20018
rect 12124 19294 12126 19346
rect 12178 19294 12180 19346
rect 12124 19282 12180 19294
rect 12908 19236 12964 19246
rect 12908 19142 12964 19180
rect 13580 19236 13636 19246
rect 13580 19142 13636 19180
rect 14252 19236 14308 19246
rect 14308 19180 14420 19236
rect 14252 19170 14308 19180
rect 11452 18452 11508 18462
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 1932 17780 1988 17790
rect 1932 17686 1988 17724
rect 4284 17668 4340 17678
rect 4284 17574 4340 17612
rect 11452 17668 11508 18396
rect 14140 18452 14196 18462
rect 14140 18358 14196 18396
rect 14252 18338 14308 18350
rect 14252 18286 14254 18338
rect 14306 18286 14308 18338
rect 14252 18228 14308 18286
rect 14252 18162 14308 18172
rect 11452 16770 11508 17612
rect 14364 17668 14420 19180
rect 14700 18452 14756 19966
rect 15148 19234 15204 20972
rect 15372 21700 15428 21710
rect 15372 20356 15428 21644
rect 15484 21698 15540 21710
rect 15484 21646 15486 21698
rect 15538 21646 15540 21698
rect 15484 21476 15540 21646
rect 16044 21698 16100 21710
rect 16044 21646 16046 21698
rect 16098 21646 16100 21698
rect 15596 21588 15652 21598
rect 15596 21586 15876 21588
rect 15596 21534 15598 21586
rect 15650 21534 15876 21586
rect 15596 21532 15876 21534
rect 15596 21522 15652 21532
rect 15484 21410 15540 21420
rect 15372 20290 15428 20300
rect 15708 20804 15764 20814
rect 15708 20242 15764 20748
rect 15708 20190 15710 20242
rect 15762 20190 15764 20242
rect 15708 20178 15764 20190
rect 15820 20242 15876 21532
rect 15820 20190 15822 20242
rect 15874 20190 15876 20242
rect 15820 20132 15876 20190
rect 15260 20018 15316 20030
rect 15484 20020 15540 20030
rect 15260 19966 15262 20018
rect 15314 19966 15316 20018
rect 15260 19796 15316 19966
rect 15260 19730 15316 19740
rect 15372 20018 15540 20020
rect 15372 19966 15486 20018
rect 15538 19966 15540 20018
rect 15372 19964 15540 19966
rect 15260 19460 15316 19470
rect 15372 19460 15428 19964
rect 15484 19954 15540 19964
rect 15596 19908 15652 19918
rect 15596 19814 15652 19852
rect 15316 19404 15428 19460
rect 15484 19460 15540 19470
rect 15260 19394 15316 19404
rect 15484 19236 15540 19404
rect 15148 19182 15150 19234
rect 15202 19182 15204 19234
rect 15148 19170 15204 19182
rect 15260 19234 15540 19236
rect 15260 19182 15486 19234
rect 15538 19182 15540 19234
rect 15260 19180 15540 19182
rect 15260 19012 15316 19180
rect 15484 19170 15540 19180
rect 15820 19124 15876 20076
rect 15596 19122 15876 19124
rect 15596 19070 15822 19122
rect 15874 19070 15876 19122
rect 15596 19068 15876 19070
rect 15036 18956 15316 19012
rect 15372 19010 15428 19022
rect 15372 18958 15374 19010
rect 15426 18958 15428 19010
rect 14812 18452 14868 18462
rect 14700 18450 14868 18452
rect 14700 18398 14814 18450
rect 14866 18398 14868 18450
rect 14700 18396 14868 18398
rect 14476 18340 14532 18350
rect 14476 18246 14532 18284
rect 14364 17612 14756 17668
rect 14364 16884 14420 17612
rect 14588 17444 14644 17454
rect 13692 16882 14420 16884
rect 13692 16830 14366 16882
rect 14418 16830 14420 16882
rect 13692 16828 14420 16830
rect 13580 16772 13636 16782
rect 11452 16718 11454 16770
rect 11506 16718 11508 16770
rect 11452 16706 11508 16718
rect 13468 16770 13636 16772
rect 13468 16718 13582 16770
rect 13634 16718 13636 16770
rect 13468 16716 13636 16718
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 13468 15986 13524 16716
rect 13580 16706 13636 16716
rect 13468 15934 13470 15986
rect 13522 15934 13524 15986
rect 13468 15922 13524 15934
rect 13692 15314 13748 16828
rect 14364 16818 14420 16828
rect 14476 17442 14644 17444
rect 14476 17390 14590 17442
rect 14642 17390 14644 17442
rect 14476 17388 14644 17390
rect 14476 16660 14532 17388
rect 14588 17378 14644 17388
rect 14700 17108 14756 17612
rect 14812 17444 14868 18396
rect 15036 18450 15092 18956
rect 15036 18398 15038 18450
rect 15090 18398 15092 18450
rect 15036 18386 15092 18398
rect 15372 18452 15428 18958
rect 15484 18564 15540 18574
rect 15596 18564 15652 19068
rect 15820 19058 15876 19068
rect 15932 21476 15988 21486
rect 15484 18562 15652 18564
rect 15484 18510 15486 18562
rect 15538 18510 15652 18562
rect 15484 18508 15652 18510
rect 15484 18498 15540 18508
rect 15372 18386 15428 18396
rect 15820 18452 15876 18462
rect 15820 18358 15876 18396
rect 14924 18338 14980 18350
rect 14924 18286 14926 18338
rect 14978 18286 14980 18338
rect 14924 17890 14980 18286
rect 15260 18228 15316 18238
rect 15260 18134 15316 18172
rect 14924 17838 14926 17890
rect 14978 17838 14980 17890
rect 14924 17826 14980 17838
rect 15148 17668 15204 17678
rect 15708 17668 15764 17678
rect 15148 17666 15764 17668
rect 15148 17614 15150 17666
rect 15202 17614 15710 17666
rect 15762 17614 15764 17666
rect 15148 17612 15764 17614
rect 15148 17602 15204 17612
rect 15708 17602 15764 17612
rect 15932 17556 15988 21420
rect 16044 18564 16100 21646
rect 16156 21588 16212 21598
rect 16156 21494 16212 21532
rect 16492 21586 16548 21598
rect 16492 21534 16494 21586
rect 16546 21534 16548 21586
rect 16492 20804 16548 21534
rect 16492 20738 16548 20748
rect 16268 20356 16324 20366
rect 16324 20300 16436 20356
rect 16268 20290 16324 20300
rect 16156 20132 16212 20142
rect 16156 19234 16212 20076
rect 16156 19182 16158 19234
rect 16210 19182 16212 19234
rect 16156 19170 16212 19182
rect 16380 19124 16436 20300
rect 16604 20244 16660 23212
rect 16828 23266 16884 23772
rect 18172 23826 18228 23838
rect 18172 23774 18174 23826
rect 18226 23774 18228 23826
rect 16828 23214 16830 23266
rect 16882 23214 16884 23266
rect 16828 23202 16884 23214
rect 16940 23716 16996 23726
rect 16828 21812 16884 21822
rect 16940 21812 16996 23660
rect 17500 23604 17556 23614
rect 17276 23492 17332 23502
rect 17276 23268 17332 23436
rect 17276 22370 17332 23212
rect 17276 22318 17278 22370
rect 17330 22318 17332 22370
rect 17276 22306 17332 22318
rect 16828 21810 16996 21812
rect 16828 21758 16830 21810
rect 16882 21758 16996 21810
rect 16828 21756 16996 21758
rect 16828 21746 16884 21756
rect 17500 21700 17556 23548
rect 18060 22258 18116 22270
rect 18060 22206 18062 22258
rect 18114 22206 18116 22258
rect 17612 21812 17668 21822
rect 17612 21718 17668 21756
rect 18060 21810 18116 22206
rect 18060 21758 18062 21810
rect 18114 21758 18116 21810
rect 18060 21746 18116 21758
rect 17836 21700 17892 21710
rect 17276 21588 17332 21598
rect 17276 21494 17332 21532
rect 17500 21474 17556 21644
rect 17500 21422 17502 21474
rect 17554 21422 17556 21474
rect 17500 21410 17556 21422
rect 17724 21698 17892 21700
rect 17724 21646 17838 21698
rect 17890 21646 17892 21698
rect 17724 21644 17892 21646
rect 16492 20132 16548 20142
rect 16604 20132 16660 20188
rect 16492 20130 16660 20132
rect 16492 20078 16494 20130
rect 16546 20078 16660 20130
rect 16492 20076 16660 20078
rect 16716 20132 16772 20142
rect 16492 20066 16548 20076
rect 16716 20018 16772 20076
rect 16716 19966 16718 20018
rect 16770 19966 16772 20018
rect 16716 19954 16772 19966
rect 16716 19236 16772 19246
rect 16492 19124 16548 19134
rect 16380 19122 16548 19124
rect 16380 19070 16494 19122
rect 16546 19070 16548 19122
rect 16380 19068 16548 19070
rect 16492 19058 16548 19068
rect 16044 18508 16212 18564
rect 16044 18340 16100 18350
rect 16044 17666 16100 18284
rect 16044 17614 16046 17666
rect 16098 17614 16100 17666
rect 16044 17602 16100 17614
rect 15932 17462 15988 17500
rect 14812 17378 14868 17388
rect 16044 17444 16100 17454
rect 14812 17108 14868 17118
rect 14700 17106 14868 17108
rect 14700 17054 14814 17106
rect 14866 17054 14868 17106
rect 14700 17052 14868 17054
rect 14812 17042 14868 17052
rect 16044 16994 16100 17388
rect 16044 16942 16046 16994
rect 16098 16942 16100 16994
rect 16044 16930 16100 16942
rect 13804 16604 14532 16660
rect 15820 16884 15876 16894
rect 13804 16098 13860 16604
rect 13804 16046 13806 16098
rect 13858 16046 13860 16098
rect 13804 16034 13860 16046
rect 15820 16098 15876 16828
rect 16156 16324 16212 18508
rect 16716 17444 16772 19180
rect 17612 19124 17668 19134
rect 17612 19030 17668 19068
rect 16828 19010 16884 19022
rect 16828 18958 16830 19010
rect 16882 18958 16884 19010
rect 16828 18676 16884 18958
rect 17724 19012 17780 21644
rect 17836 21634 17892 21644
rect 18172 19460 18228 23774
rect 19516 23828 19572 23838
rect 18284 23716 18340 23726
rect 18284 23622 18340 23660
rect 18508 22372 18564 22382
rect 18284 21700 18340 21710
rect 18284 21606 18340 21644
rect 18396 21586 18452 21598
rect 18396 21534 18398 21586
rect 18450 21534 18452 21586
rect 18284 20132 18340 20142
rect 18396 20132 18452 21534
rect 18508 21476 18564 22316
rect 18508 21410 18564 21420
rect 18620 20244 18676 20254
rect 18620 20150 18676 20188
rect 18340 20076 18452 20132
rect 18508 20130 18564 20142
rect 18508 20078 18510 20130
rect 18562 20078 18564 20130
rect 18284 20066 18340 20076
rect 18508 20020 18564 20078
rect 19180 20130 19236 20142
rect 19180 20078 19182 20130
rect 19234 20078 19236 20130
rect 19068 20020 19124 20030
rect 18172 19366 18228 19404
rect 18396 19964 18564 20020
rect 18620 20018 19124 20020
rect 18620 19966 19070 20018
rect 19122 19966 19124 20018
rect 18620 19964 19124 19966
rect 17948 19236 18004 19246
rect 17948 19142 18004 19180
rect 17724 18900 17780 18956
rect 16828 18610 16884 18620
rect 17500 18844 17780 18900
rect 18060 19124 18116 19134
rect 16716 17378 16772 17388
rect 16604 17108 16660 17118
rect 17276 17108 17332 17118
rect 16604 16882 16660 17052
rect 16604 16830 16606 16882
rect 16658 16830 16660 16882
rect 16604 16818 16660 16830
rect 17164 17052 17276 17108
rect 16156 16100 16212 16268
rect 15820 16046 15822 16098
rect 15874 16046 15876 16098
rect 15820 16034 15876 16046
rect 15932 16044 16212 16100
rect 16268 16770 16324 16782
rect 16268 16718 16270 16770
rect 16322 16718 16324 16770
rect 16268 16100 16324 16718
rect 16716 16100 16772 16110
rect 16268 16098 16548 16100
rect 16268 16046 16270 16098
rect 16322 16046 16548 16098
rect 16268 16044 16548 16046
rect 14364 15876 14420 15886
rect 14364 15426 14420 15820
rect 15484 15876 15540 15886
rect 15484 15782 15540 15820
rect 15708 15876 15764 15886
rect 15932 15876 15988 16044
rect 16268 16034 16324 16044
rect 15708 15874 15988 15876
rect 15708 15822 15710 15874
rect 15762 15822 15988 15874
rect 15708 15820 15988 15822
rect 15708 15810 15764 15820
rect 14364 15374 14366 15426
rect 14418 15374 14420 15426
rect 14364 15362 14420 15374
rect 16492 15540 16548 16044
rect 16716 16006 16772 16044
rect 13692 15262 13694 15314
rect 13746 15262 13748 15314
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 13692 14644 13748 15262
rect 16492 15202 16548 15484
rect 16492 15150 16494 15202
rect 16546 15150 16548 15202
rect 16492 15138 16548 15150
rect 17164 15986 17220 17052
rect 17276 17042 17332 17052
rect 17500 16994 17556 18844
rect 18060 18452 18116 19068
rect 18284 19010 18340 19022
rect 18284 18958 18286 19010
rect 18338 18958 18340 19010
rect 18060 17554 18116 18396
rect 18060 17502 18062 17554
rect 18114 17502 18116 17554
rect 18060 17490 18116 17502
rect 18172 18676 18228 18686
rect 18172 18562 18228 18620
rect 18172 18510 18174 18562
rect 18226 18510 18228 18562
rect 18060 17108 18116 17118
rect 17500 16942 17502 16994
rect 17554 16942 17556 16994
rect 17276 16884 17332 16894
rect 17276 16790 17332 16828
rect 17500 16884 17556 16942
rect 17612 16996 17668 17006
rect 17612 16902 17668 16940
rect 17500 16818 17556 16828
rect 18060 16882 18116 17052
rect 18060 16830 18062 16882
rect 18114 16830 18116 16882
rect 18060 16818 18116 16830
rect 17388 16772 17444 16782
rect 17276 16324 17332 16334
rect 17388 16324 17444 16716
rect 17332 16268 17444 16324
rect 17276 16210 17332 16268
rect 17276 16158 17278 16210
rect 17330 16158 17332 16210
rect 17276 16146 17332 16158
rect 17612 16100 17668 16138
rect 17612 16034 17668 16044
rect 18172 16100 18228 18510
rect 18284 18564 18340 18958
rect 18284 18498 18340 18508
rect 18396 18674 18452 19964
rect 18508 19236 18564 19246
rect 18620 19236 18676 19964
rect 19068 19954 19124 19964
rect 19180 19908 19236 20078
rect 19292 20132 19348 20142
rect 19292 20020 19348 20076
rect 19516 20132 19572 23772
rect 19628 22372 19684 23886
rect 20076 23826 20132 23838
rect 20076 23774 20078 23826
rect 20130 23774 20132 23826
rect 20076 23716 20132 23774
rect 20300 23828 20356 23838
rect 20300 23734 20356 23772
rect 20076 23660 20244 23716
rect 20188 23604 20244 23660
rect 19836 23548 20100 23558
rect 20188 23548 20356 23604
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 20188 23268 20244 23278
rect 20188 23174 20244 23212
rect 20300 22820 20356 23548
rect 20076 22764 20356 22820
rect 20748 23268 20804 24668
rect 19740 22372 19796 22382
rect 19628 22316 19740 22372
rect 19740 22306 19796 22316
rect 20076 22260 20132 22764
rect 20188 22484 20244 22494
rect 20636 22484 20692 22494
rect 20748 22484 20804 23212
rect 20188 22482 20356 22484
rect 20188 22430 20190 22482
rect 20242 22430 20356 22482
rect 20188 22428 20356 22430
rect 20188 22418 20244 22428
rect 20076 22204 20244 22260
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 20188 21812 20244 22204
rect 20188 21718 20244 21756
rect 20300 21028 20356 22428
rect 20636 22482 20748 22484
rect 20636 22430 20638 22482
rect 20690 22430 20748 22482
rect 20636 22428 20748 22430
rect 20636 22418 20692 22428
rect 20748 22390 20804 22428
rect 21196 24724 21252 24734
rect 20412 21588 20468 21598
rect 20468 21532 20580 21588
rect 20412 21494 20468 21532
rect 20412 21028 20468 21038
rect 20300 21026 20468 21028
rect 20300 20974 20414 21026
rect 20466 20974 20468 21026
rect 20300 20972 20468 20974
rect 20188 20580 20244 20590
rect 20188 20486 20244 20524
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 20300 20188 20356 20972
rect 20412 20962 20468 20972
rect 20524 20914 20580 21532
rect 20524 20862 20526 20914
rect 20578 20862 20580 20914
rect 20524 20850 20580 20862
rect 21196 21586 21252 24668
rect 21532 24610 21588 24622
rect 21532 24558 21534 24610
rect 21586 24558 21588 24610
rect 21532 23714 21588 24558
rect 21868 24052 21924 24062
rect 21868 23958 21924 23996
rect 22204 24052 22260 24062
rect 21644 23940 21700 23950
rect 21644 23846 21700 23884
rect 22092 23938 22148 23950
rect 22092 23886 22094 23938
rect 22146 23886 22148 23938
rect 22092 23828 22148 23886
rect 22092 23762 22148 23772
rect 21532 23662 21534 23714
rect 21586 23662 21588 23714
rect 21532 23650 21588 23662
rect 21420 22484 21476 22494
rect 21420 22390 21476 22428
rect 21868 22372 21924 22382
rect 21868 22278 21924 22316
rect 22092 22146 22148 22158
rect 22092 22094 22094 22146
rect 22146 22094 22148 22146
rect 21420 21700 21476 21710
rect 21420 21606 21476 21644
rect 21196 21534 21198 21586
rect 21250 21534 21252 21586
rect 19516 20066 19572 20076
rect 19740 20132 20356 20188
rect 20636 20578 20692 20590
rect 20636 20526 20638 20578
rect 20690 20526 20692 20578
rect 20636 20132 20692 20526
rect 21196 20242 21252 21534
rect 22092 21588 22148 22094
rect 22092 21522 22148 21532
rect 21308 20802 21364 20814
rect 21308 20750 21310 20802
rect 21362 20750 21364 20802
rect 21308 20580 21364 20750
rect 21308 20514 21364 20524
rect 21196 20190 21198 20242
rect 21250 20190 21252 20242
rect 21196 20178 21252 20190
rect 19740 20130 19796 20132
rect 19740 20078 19742 20130
rect 19794 20078 19796 20130
rect 19740 20066 19796 20078
rect 19404 20020 19460 20030
rect 19292 20018 19460 20020
rect 19292 19966 19406 20018
rect 19458 19966 19460 20018
rect 19292 19964 19460 19966
rect 19404 19954 19460 19964
rect 18732 19796 18788 19806
rect 18732 19702 18788 19740
rect 19068 19796 19124 19806
rect 18564 19180 18676 19236
rect 18508 19142 18564 19180
rect 18956 19012 19012 19022
rect 18956 18918 19012 18956
rect 18396 18622 18398 18674
rect 18450 18622 18452 18674
rect 18284 18338 18340 18350
rect 18284 18286 18286 18338
rect 18338 18286 18340 18338
rect 18284 18228 18340 18286
rect 18284 18162 18340 18172
rect 18396 18116 18452 18622
rect 19068 18674 19124 19740
rect 19180 19460 19236 19852
rect 19628 19796 19684 19806
rect 19628 19702 19684 19740
rect 19740 19460 19796 19470
rect 19180 19404 19572 19460
rect 19180 19236 19236 19246
rect 19180 19142 19236 19180
rect 19404 19124 19460 19134
rect 19404 19030 19460 19068
rect 19068 18622 19070 18674
rect 19122 18622 19124 18674
rect 19068 18610 19124 18622
rect 19292 19010 19348 19022
rect 19292 18958 19294 19010
rect 19346 18958 19348 19010
rect 18844 18452 18900 18462
rect 18844 18450 19012 18452
rect 18844 18398 18846 18450
rect 18898 18398 19012 18450
rect 18844 18396 19012 18398
rect 18844 18386 18900 18396
rect 18396 18050 18452 18060
rect 18956 17780 19012 18396
rect 19292 17892 19348 18958
rect 19292 17826 19348 17836
rect 19404 18452 19460 18462
rect 18956 17714 19012 17724
rect 18844 17668 18900 17678
rect 18620 17666 18900 17668
rect 18620 17614 18846 17666
rect 18898 17614 18900 17666
rect 18620 17612 18900 17614
rect 18620 17556 18676 17612
rect 18844 17602 18900 17612
rect 18508 17500 18676 17556
rect 18956 17556 19012 17566
rect 19012 17500 19124 17556
rect 18172 16034 18228 16044
rect 18396 17444 18452 17454
rect 18508 17444 18564 17500
rect 18956 17490 19012 17500
rect 18732 17444 18788 17454
rect 18396 17442 18564 17444
rect 18396 17390 18398 17442
rect 18450 17390 18564 17442
rect 18396 17388 18564 17390
rect 18620 17442 18788 17444
rect 18620 17390 18734 17442
rect 18786 17390 18788 17442
rect 18620 17388 18788 17390
rect 17164 15934 17166 15986
rect 17218 15934 17220 15986
rect 13692 14578 13748 14588
rect 15372 14644 15428 14654
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 15372 12962 15428 14588
rect 16716 14644 16772 14654
rect 16716 14550 16772 14588
rect 16044 14308 16100 14318
rect 16044 13074 16100 14252
rect 17164 14308 17220 15934
rect 17388 15540 17444 15550
rect 17388 15446 17444 15484
rect 17948 15316 18004 15326
rect 17948 15222 18004 15260
rect 18396 15316 18452 17388
rect 18620 16996 18676 17388
rect 18732 17378 18788 17388
rect 18620 16902 18676 16940
rect 18396 15250 18452 15260
rect 18508 16100 18564 16110
rect 18508 15314 18564 16044
rect 18508 15262 18510 15314
rect 18562 15262 18564 15314
rect 18508 15250 18564 15262
rect 18844 16098 18900 16110
rect 18844 16046 18846 16098
rect 18898 16046 18900 16098
rect 18844 15314 18900 16046
rect 19068 15538 19124 17500
rect 19068 15486 19070 15538
rect 19122 15486 19124 15538
rect 19068 15474 19124 15486
rect 19180 16884 19236 16894
rect 18844 15262 18846 15314
rect 18898 15262 18900 15314
rect 18732 14644 18788 14654
rect 17164 14242 17220 14252
rect 17612 14418 17668 14430
rect 17612 14366 17614 14418
rect 17666 14366 17668 14418
rect 17612 14308 17668 14366
rect 17948 14418 18004 14430
rect 17948 14366 17950 14418
rect 18002 14366 18004 14418
rect 17948 14308 18004 14366
rect 18284 14308 18340 14318
rect 17948 14306 18340 14308
rect 17948 14254 18286 14306
rect 18338 14254 18340 14306
rect 17948 14252 18340 14254
rect 17612 14242 17668 14252
rect 16044 13022 16046 13074
rect 16098 13022 16100 13074
rect 16044 13010 16100 13022
rect 18172 13076 18228 13086
rect 18284 13076 18340 14252
rect 18172 13074 18340 13076
rect 18172 13022 18174 13074
rect 18226 13022 18340 13074
rect 18172 13020 18340 13022
rect 18732 13746 18788 14588
rect 18844 14644 18900 15262
rect 18844 14642 19124 14644
rect 18844 14590 18846 14642
rect 18898 14590 19124 14642
rect 18844 14588 19124 14590
rect 18844 14578 18900 14588
rect 19068 14196 19124 14588
rect 19180 14418 19236 16828
rect 19404 15148 19460 18396
rect 19516 17442 19572 19404
rect 19740 19346 19796 19404
rect 19740 19294 19742 19346
rect 19794 19294 19796 19346
rect 19740 19282 19796 19294
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 20188 18788 20244 20132
rect 20636 20066 20692 20076
rect 21756 20132 21812 20142
rect 21756 20038 21812 20076
rect 20860 20018 20916 20030
rect 20860 19966 20862 20018
rect 20914 19966 20916 20018
rect 20300 19236 20356 19246
rect 20300 19142 20356 19180
rect 20524 19234 20580 19246
rect 20524 19182 20526 19234
rect 20578 19182 20580 19234
rect 20524 19124 20580 19182
rect 20580 19068 20804 19124
rect 20524 19058 20580 19068
rect 20636 18788 20692 18798
rect 20188 18732 20636 18788
rect 20636 18450 20692 18732
rect 20636 18398 20638 18450
rect 20690 18398 20692 18450
rect 20636 18386 20692 18398
rect 19628 18338 19684 18350
rect 19628 18286 19630 18338
rect 19682 18286 19684 18338
rect 19628 18004 19684 18286
rect 20524 18340 20580 18350
rect 20524 18246 20580 18284
rect 20412 18116 20468 18126
rect 20468 18060 20692 18116
rect 20412 18050 20468 18060
rect 19628 17938 19684 17948
rect 20300 18004 20356 18014
rect 19852 17780 19908 17790
rect 19852 17666 19908 17724
rect 19852 17614 19854 17666
rect 19906 17614 19908 17666
rect 19852 17602 19908 17614
rect 19516 17390 19518 17442
rect 19570 17390 19572 17442
rect 19516 17378 19572 17390
rect 20188 17444 20244 17454
rect 20188 17350 20244 17388
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 19516 17108 19572 17118
rect 19516 17014 19572 17052
rect 20188 16884 20244 16894
rect 20300 16884 20356 17948
rect 20188 16882 20356 16884
rect 20188 16830 20190 16882
rect 20242 16830 20356 16882
rect 20188 16828 20356 16830
rect 20524 17666 20580 17678
rect 20524 17614 20526 17666
rect 20578 17614 20580 17666
rect 20188 16818 20244 16828
rect 19740 16212 19796 16222
rect 19628 16156 19740 16212
rect 19628 15316 19684 16156
rect 19740 16146 19796 16156
rect 19852 16098 19908 16110
rect 19852 16046 19854 16098
rect 19906 16046 19908 16098
rect 19852 15876 19908 16046
rect 20412 15986 20468 15998
rect 20412 15934 20414 15986
rect 20466 15934 20468 15986
rect 19852 15820 20244 15876
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 19740 15316 19796 15326
rect 19628 15314 19796 15316
rect 19628 15262 19742 15314
rect 19794 15262 19796 15314
rect 19628 15260 19796 15262
rect 19740 15250 19796 15260
rect 20188 15316 20244 15820
rect 20188 15222 20244 15260
rect 19404 15092 19908 15148
rect 19852 14754 19908 15092
rect 19852 14702 19854 14754
rect 19906 14702 19908 14754
rect 19852 14690 19908 14702
rect 19964 15090 20020 15102
rect 20412 15092 20468 15934
rect 20524 15540 20580 17614
rect 20636 16994 20692 18060
rect 20748 17780 20804 19068
rect 20860 18004 20916 19966
rect 21084 19906 21140 19918
rect 21084 19854 21086 19906
rect 21138 19854 21140 19906
rect 20860 17938 20916 17948
rect 20972 19012 21028 19022
rect 20972 18450 21028 18956
rect 20972 18398 20974 18450
rect 21026 18398 21028 18450
rect 20748 17686 20804 17724
rect 20636 16942 20638 16994
rect 20690 16942 20692 16994
rect 20636 16212 20692 16942
rect 20636 16146 20692 16156
rect 20748 16100 20804 16110
rect 20972 16100 21028 18398
rect 20748 16098 21028 16100
rect 20748 16046 20750 16098
rect 20802 16046 21028 16098
rect 20748 16044 21028 16046
rect 20636 15540 20692 15550
rect 20524 15484 20636 15540
rect 20636 15446 20692 15484
rect 20748 15316 20804 16044
rect 20748 15250 20804 15260
rect 19964 15038 19966 15090
rect 20018 15038 20020 15090
rect 19180 14366 19182 14418
rect 19234 14366 19236 14418
rect 19180 14354 19236 14366
rect 19404 14532 19460 14542
rect 19964 14532 20020 15038
rect 19404 14530 20020 14532
rect 19404 14478 19406 14530
rect 19458 14478 20020 14530
rect 19404 14476 20020 14478
rect 20188 15036 20412 15092
rect 20188 14530 20244 15036
rect 20412 15026 20468 15036
rect 21084 15092 21140 19854
rect 21868 19906 21924 19918
rect 21868 19854 21870 19906
rect 21922 19854 21924 19906
rect 21644 19012 21700 19022
rect 21868 19012 21924 19854
rect 21980 19236 22036 19246
rect 21980 19122 22036 19180
rect 21980 19070 21982 19122
rect 22034 19070 22036 19122
rect 21980 19058 22036 19070
rect 21700 18956 21924 19012
rect 21644 18918 21700 18956
rect 22204 18564 22260 23996
rect 22540 23940 22596 25340
rect 22764 25330 22820 25340
rect 22876 25282 22932 25294
rect 22876 25230 22878 25282
rect 22930 25230 22932 25282
rect 22876 24164 22932 25230
rect 22876 24098 22932 24108
rect 22988 24612 23044 24622
rect 22988 24050 23044 24556
rect 23324 24500 23380 26236
rect 23660 24612 23716 24622
rect 23772 24612 23828 31892
rect 24332 27748 24388 27758
rect 24332 27654 24388 27692
rect 25228 27748 25284 37214
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 25228 27682 25284 27692
rect 37884 27858 37940 27870
rect 37884 27806 37886 27858
rect 37938 27806 37940 27858
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 27580 27186 27636 27198
rect 27580 27134 27582 27186
rect 27634 27134 27636 27186
rect 24556 27074 24612 27086
rect 24556 27022 24558 27074
rect 24610 27022 24612 27074
rect 24556 26908 24612 27022
rect 26908 27076 26964 27086
rect 25340 26964 25396 26974
rect 24220 26852 24612 26908
rect 25228 26962 25396 26964
rect 25228 26910 25342 26962
rect 25394 26910 25396 26962
rect 25228 26908 25396 26910
rect 24220 26850 24276 26852
rect 24220 26798 24222 26850
rect 24274 26798 24276 26850
rect 23884 25284 23940 25294
rect 24220 25284 24276 26798
rect 23940 25228 24276 25284
rect 24556 26404 24612 26414
rect 23884 25190 23940 25228
rect 24556 24946 24612 26348
rect 25228 26068 25284 26908
rect 25340 26898 25396 26908
rect 25900 26516 25956 26526
rect 25900 26422 25956 26460
rect 26908 26516 26964 27020
rect 27580 27076 27636 27134
rect 27580 27010 27636 27020
rect 28140 27076 28196 27086
rect 28140 26982 28196 27020
rect 37660 27076 37716 27086
rect 37660 26982 37716 27020
rect 28364 26964 28420 26974
rect 28364 26870 28420 26908
rect 37884 26964 37940 27806
rect 40012 27636 40068 27646
rect 40012 27542 40068 27580
rect 37884 26898 37940 26908
rect 40012 27186 40068 27198
rect 40012 27134 40014 27186
rect 40066 27134 40068 27186
rect 25340 26404 25396 26414
rect 25340 26310 25396 26348
rect 25452 26292 25508 26302
rect 25676 26292 25732 26302
rect 25452 26290 25732 26292
rect 25452 26238 25454 26290
rect 25506 26238 25678 26290
rect 25730 26238 25732 26290
rect 25452 26236 25732 26238
rect 25452 26226 25508 26236
rect 25676 26226 25732 26236
rect 26012 26292 26068 26302
rect 26012 26198 26068 26236
rect 26908 26290 26964 26460
rect 39900 26852 39956 26862
rect 27132 26404 27188 26414
rect 27132 26310 27188 26348
rect 26908 26238 26910 26290
rect 26962 26238 26964 26290
rect 26908 26226 26964 26238
rect 37660 26292 37716 26302
rect 37660 26198 37716 26236
rect 39900 26178 39956 26796
rect 40012 26292 40068 27134
rect 40012 26226 40068 26236
rect 39900 26126 39902 26178
rect 39954 26126 39956 26178
rect 39900 26114 39956 26126
rect 25340 26068 25396 26078
rect 25228 26066 25396 26068
rect 25228 26014 25342 26066
rect 25394 26014 25396 26066
rect 25228 26012 25396 26014
rect 25340 26002 25396 26012
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 25116 25284 25172 25294
rect 25172 25228 25284 25284
rect 25116 25218 25172 25228
rect 24556 24894 24558 24946
rect 24610 24894 24612 24946
rect 24556 24882 24612 24894
rect 24332 24834 24388 24846
rect 24332 24782 24334 24834
rect 24386 24782 24388 24834
rect 23716 24556 23828 24612
rect 24220 24722 24276 24734
rect 24220 24670 24222 24722
rect 24274 24670 24276 24722
rect 23660 24518 23716 24556
rect 22988 23998 22990 24050
rect 23042 23998 23044 24050
rect 22988 23986 23044 23998
rect 23100 24444 23380 24500
rect 22540 23874 22596 23884
rect 22652 23940 22708 23950
rect 22876 23940 22932 23950
rect 22652 23938 22932 23940
rect 22652 23886 22654 23938
rect 22706 23886 22878 23938
rect 22930 23886 22932 23938
rect 22652 23884 22932 23886
rect 22652 23874 22708 23884
rect 22876 23874 22932 23884
rect 22316 23828 22372 23838
rect 22316 23734 22372 23772
rect 22428 22484 22484 22494
rect 22428 22370 22484 22428
rect 22428 22318 22430 22370
rect 22482 22318 22484 22370
rect 22428 22306 22484 22318
rect 23100 22036 23156 24444
rect 23772 24164 23828 24174
rect 23436 23940 23492 23950
rect 23212 22260 23268 22270
rect 23212 22258 23380 22260
rect 23212 22206 23214 22258
rect 23266 22206 23380 22258
rect 23212 22204 23380 22206
rect 23212 22194 23268 22204
rect 23100 21980 23268 22036
rect 23100 20132 23156 20142
rect 23100 20038 23156 20076
rect 22876 19794 22932 19806
rect 22876 19742 22878 19794
rect 22930 19742 22932 19794
rect 22540 19234 22596 19246
rect 22540 19182 22542 19234
rect 22594 19182 22596 19234
rect 22316 19124 22372 19134
rect 22316 19030 22372 19068
rect 22540 18788 22596 19182
rect 22540 18722 22596 18732
rect 22316 18564 22372 18574
rect 22204 18562 22372 18564
rect 22204 18510 22318 18562
rect 22370 18510 22372 18562
rect 22204 18508 22372 18510
rect 21980 18450 22036 18462
rect 21980 18398 21982 18450
rect 22034 18398 22036 18450
rect 21980 18340 22036 18398
rect 21980 18274 22036 18284
rect 21308 16212 21364 16222
rect 21308 16118 21364 16156
rect 21756 16100 21812 16110
rect 21084 15026 21140 15036
rect 21644 16098 21812 16100
rect 21644 16046 21758 16098
rect 21810 16046 21812 16098
rect 21644 16044 21812 16046
rect 21644 15314 21700 16044
rect 21756 16034 21812 16044
rect 21644 15262 21646 15314
rect 21698 15262 21700 15314
rect 20188 14478 20190 14530
rect 20242 14478 20244 14530
rect 19404 14196 19460 14476
rect 20188 14466 20244 14478
rect 19964 14308 20020 14318
rect 19068 14140 19460 14196
rect 19628 14306 20020 14308
rect 19628 14254 19966 14306
rect 20018 14254 20020 14306
rect 19628 14252 20020 14254
rect 19516 13860 19572 13870
rect 19628 13860 19684 14252
rect 19964 14242 20020 14252
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 19516 13858 19684 13860
rect 19516 13806 19518 13858
rect 19570 13806 19684 13858
rect 19516 13804 19684 13806
rect 19516 13794 19572 13804
rect 18732 13694 18734 13746
rect 18786 13694 18788 13746
rect 18732 13074 18788 13694
rect 21644 13634 21700 15262
rect 22092 15316 22148 15326
rect 22316 15316 22372 18508
rect 22876 18452 22932 19742
rect 23212 19794 23268 21980
rect 23324 21810 23380 22204
rect 23324 21758 23326 21810
rect 23378 21758 23380 21810
rect 23324 21746 23380 21758
rect 23436 21812 23492 23884
rect 23660 23938 23716 23950
rect 23660 23886 23662 23938
rect 23714 23886 23716 23938
rect 23660 23156 23716 23886
rect 23660 23090 23716 23100
rect 23772 21812 23828 24108
rect 24108 23938 24164 23950
rect 24108 23886 24110 23938
rect 24162 23886 24164 23938
rect 23996 23826 24052 23838
rect 23996 23774 23998 23826
rect 24050 23774 24052 23826
rect 23884 23716 23940 23726
rect 23884 23622 23940 23660
rect 23996 22596 24052 23774
rect 23996 22530 24052 22540
rect 24108 23828 24164 23886
rect 23884 21812 23940 21822
rect 23436 21756 23604 21812
rect 23772 21756 23884 21812
rect 23436 21586 23492 21598
rect 23436 21534 23438 21586
rect 23490 21534 23492 21586
rect 23436 19908 23492 21534
rect 23548 21588 23604 21756
rect 23660 21588 23716 21598
rect 23548 21532 23660 21588
rect 23660 21494 23716 21532
rect 23884 21586 23940 21756
rect 23884 21534 23886 21586
rect 23938 21534 23940 21586
rect 23884 21522 23940 21534
rect 23996 21700 24052 21710
rect 24108 21700 24164 23772
rect 24220 23604 24276 24670
rect 24332 24164 24388 24782
rect 24332 24098 24388 24108
rect 24444 24052 24500 24062
rect 24444 23938 24500 23996
rect 25228 24052 25284 25228
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 27132 24052 27188 24062
rect 25228 24050 25620 24052
rect 25228 23998 25230 24050
rect 25282 23998 25620 24050
rect 25228 23996 25620 23998
rect 25228 23986 25284 23996
rect 24444 23886 24446 23938
rect 24498 23886 24500 23938
rect 24444 23874 24500 23886
rect 25564 23938 25620 23996
rect 25564 23886 25566 23938
rect 25618 23886 25620 23938
rect 24220 23538 24276 23548
rect 24556 23714 24612 23726
rect 24556 23662 24558 23714
rect 24610 23662 24612 23714
rect 24556 23604 24612 23662
rect 24556 23538 24612 23548
rect 25228 23604 25284 23614
rect 24052 21644 24164 21700
rect 24668 23154 24724 23166
rect 24668 23102 24670 23154
rect 24722 23102 24724 23154
rect 23996 21586 24052 21644
rect 24332 21588 24388 21598
rect 23996 21534 23998 21586
rect 24050 21534 24052 21586
rect 23996 21522 24052 21534
rect 24220 21586 24388 21588
rect 24220 21534 24334 21586
rect 24386 21534 24388 21586
rect 24220 21532 24388 21534
rect 23548 20132 23604 20142
rect 23548 20038 23604 20076
rect 23884 20130 23940 20142
rect 23884 20078 23886 20130
rect 23938 20078 23940 20130
rect 23884 19908 23940 20078
rect 23436 19852 23940 19908
rect 23212 19742 23214 19794
rect 23266 19742 23268 19794
rect 23212 19460 23268 19742
rect 23884 19572 23940 19852
rect 23884 19506 23940 19516
rect 23212 19394 23268 19404
rect 24220 19458 24276 21532
rect 24332 21522 24388 21532
rect 24668 20692 24724 23102
rect 25228 21698 25284 23548
rect 25564 23380 25620 23886
rect 26348 23826 26404 23838
rect 26348 23774 26350 23826
rect 26402 23774 26404 23826
rect 26348 23716 26404 23774
rect 26348 23650 26404 23660
rect 25676 23380 25732 23390
rect 25564 23378 26068 23380
rect 25564 23326 25678 23378
rect 25730 23326 26068 23378
rect 25564 23324 26068 23326
rect 25676 23314 25732 23324
rect 26012 23154 26068 23324
rect 26012 23102 26014 23154
rect 26066 23102 26068 23154
rect 26012 23090 26068 23102
rect 26796 23044 26852 23054
rect 26236 23042 26852 23044
rect 26236 22990 26798 23042
rect 26850 22990 26852 23042
rect 26236 22988 26852 22990
rect 25340 22484 25396 22494
rect 25452 22484 25508 22494
rect 25340 22482 25452 22484
rect 25340 22430 25342 22482
rect 25394 22430 25452 22482
rect 25340 22428 25452 22430
rect 25340 22418 25396 22428
rect 25228 21646 25230 21698
rect 25282 21646 25284 21698
rect 25228 21634 25284 21646
rect 25340 21698 25396 21710
rect 25340 21646 25342 21698
rect 25394 21646 25396 21698
rect 25116 20692 25172 20702
rect 24668 20690 25172 20692
rect 24668 20638 25118 20690
rect 25170 20638 25172 20690
rect 24668 20636 25172 20638
rect 25116 20188 25172 20636
rect 24668 20132 24724 20142
rect 25116 20132 25284 20188
rect 24668 20038 24724 20076
rect 24220 19406 24222 19458
rect 24274 19406 24276 19458
rect 24220 19394 24276 19406
rect 24332 20018 24388 20030
rect 24332 19966 24334 20018
rect 24386 19966 24388 20018
rect 24332 19236 24388 19966
rect 24332 19142 24388 19180
rect 24220 19124 24276 19134
rect 24220 19030 24276 19068
rect 23436 18562 23492 18574
rect 23436 18510 23438 18562
rect 23490 18510 23492 18562
rect 23100 18452 23156 18462
rect 22876 18450 23156 18452
rect 22876 18398 23102 18450
rect 23154 18398 23156 18450
rect 22876 18396 23156 18398
rect 23100 18004 23156 18396
rect 23436 18340 23492 18510
rect 23884 18564 23940 18574
rect 23884 18562 24052 18564
rect 23884 18510 23886 18562
rect 23938 18510 24052 18562
rect 23884 18508 24052 18510
rect 23884 18498 23940 18508
rect 23772 18450 23828 18462
rect 23772 18398 23774 18450
rect 23826 18398 23828 18450
rect 23492 18284 23604 18340
rect 23436 18274 23492 18284
rect 23100 17938 23156 17948
rect 23436 17892 23492 17902
rect 22988 17554 23044 17566
rect 22988 17502 22990 17554
rect 23042 17502 23044 17554
rect 22988 16098 23044 17502
rect 23436 16994 23492 17836
rect 23548 17106 23604 18284
rect 23548 17054 23550 17106
rect 23602 17054 23604 17106
rect 23548 17042 23604 17054
rect 23772 17106 23828 18398
rect 23772 17054 23774 17106
rect 23826 17054 23828 17106
rect 23772 17042 23828 17054
rect 23884 18226 23940 18238
rect 23884 18174 23886 18226
rect 23938 18174 23940 18226
rect 23436 16942 23438 16994
rect 23490 16942 23492 16994
rect 23436 16930 23492 16942
rect 23772 16212 23828 16222
rect 23884 16212 23940 18174
rect 23996 16884 24052 18508
rect 25228 17666 25284 20132
rect 25340 19572 25396 21646
rect 25452 21588 25508 22428
rect 26236 22482 26292 22988
rect 26796 22978 26852 22988
rect 26236 22430 26238 22482
rect 26290 22430 26292 22482
rect 26236 22418 26292 22430
rect 26908 22596 26964 22606
rect 25788 22372 25844 22382
rect 26348 22372 26404 22382
rect 25788 22370 26068 22372
rect 25788 22318 25790 22370
rect 25842 22318 26068 22370
rect 25788 22316 26068 22318
rect 25788 22306 25844 22316
rect 25900 22148 25956 22158
rect 25788 22146 25956 22148
rect 25788 22094 25902 22146
rect 25954 22094 25956 22146
rect 25788 22092 25956 22094
rect 25788 21924 25844 22092
rect 25900 22082 25956 22092
rect 25564 21868 25844 21924
rect 25564 21810 25620 21868
rect 25564 21758 25566 21810
rect 25618 21758 25620 21810
rect 25564 21746 25620 21758
rect 25452 21532 25732 21588
rect 25676 21252 25732 21532
rect 25676 21196 25956 21252
rect 25452 20076 25844 20132
rect 25452 20018 25508 20076
rect 25452 19966 25454 20018
rect 25506 19966 25508 20018
rect 25452 19954 25508 19966
rect 25676 19908 25732 19918
rect 25340 19506 25396 19516
rect 25564 19852 25676 19908
rect 25564 18564 25620 19852
rect 25676 19814 25732 19852
rect 25788 18564 25844 20076
rect 25900 19124 25956 21196
rect 25900 19058 25956 19068
rect 25228 17614 25230 17666
rect 25282 17614 25284 17666
rect 25228 17602 25284 17614
rect 25340 18508 25620 18564
rect 25676 18562 25844 18564
rect 25676 18510 25790 18562
rect 25842 18510 25844 18562
rect 25676 18508 25844 18510
rect 23996 16818 24052 16828
rect 25228 17444 25284 17454
rect 25228 16882 25284 17388
rect 25228 16830 25230 16882
rect 25282 16830 25284 16882
rect 25228 16818 25284 16830
rect 23772 16210 23940 16212
rect 23772 16158 23774 16210
rect 23826 16158 23940 16210
rect 23772 16156 23940 16158
rect 23996 16660 24052 16670
rect 23772 16146 23828 16156
rect 22988 16046 22990 16098
rect 23042 16046 23044 16098
rect 22876 15540 22932 15550
rect 22876 15426 22932 15484
rect 22876 15374 22878 15426
rect 22930 15374 22932 15426
rect 22876 15362 22932 15374
rect 22764 15316 22820 15326
rect 22316 15260 22764 15316
rect 22092 15222 22148 15260
rect 22764 15222 22820 15260
rect 21868 14644 21924 14654
rect 21868 14532 21924 14588
rect 22988 14644 23044 16046
rect 23324 15314 23380 15326
rect 23324 15262 23326 15314
rect 23378 15262 23380 15314
rect 22988 14578 23044 14588
rect 23100 15202 23156 15214
rect 23100 15150 23102 15202
rect 23154 15150 23156 15202
rect 21868 14530 22148 14532
rect 21868 14478 21870 14530
rect 21922 14478 22148 14530
rect 21868 14476 22148 14478
rect 21868 14466 21924 14476
rect 22092 13970 22148 14476
rect 22540 14420 22596 14430
rect 23100 14420 23156 15150
rect 23324 15148 23380 15262
rect 23996 15148 24052 16604
rect 25340 16660 25396 18508
rect 25340 15428 25396 16604
rect 25340 15362 25396 15372
rect 25452 18338 25508 18350
rect 25452 18286 25454 18338
rect 25506 18286 25508 18338
rect 25452 15764 25508 18286
rect 25564 17668 25620 17678
rect 25564 17106 25620 17612
rect 25564 17054 25566 17106
rect 25618 17054 25620 17106
rect 25564 16100 25620 17054
rect 25676 17108 25732 18508
rect 25788 18498 25844 18508
rect 26012 18228 26068 22316
rect 26348 22278 26404 22316
rect 26908 22370 26964 22540
rect 26908 22318 26910 22370
rect 26962 22318 26964 22370
rect 26908 22306 26964 22318
rect 27132 22258 27188 23996
rect 28476 24052 28532 24062
rect 28476 23958 28532 23996
rect 40012 24050 40068 24062
rect 40012 23998 40014 24050
rect 40066 23998 40068 24050
rect 37660 23940 37716 23950
rect 37660 23846 37716 23884
rect 40012 23604 40068 23998
rect 40012 23538 40068 23548
rect 37660 23156 37716 23166
rect 37660 23062 37716 23100
rect 27916 23044 27972 23054
rect 27468 22372 27524 22382
rect 27804 22372 27860 22382
rect 27468 22278 27524 22316
rect 27580 22370 27860 22372
rect 27580 22318 27806 22370
rect 27858 22318 27860 22370
rect 27580 22316 27860 22318
rect 27132 22206 27134 22258
rect 27186 22206 27188 22258
rect 27132 22194 27188 22206
rect 27244 22258 27300 22270
rect 27244 22206 27246 22258
rect 27298 22206 27300 22258
rect 26124 22146 26180 22158
rect 26124 22094 26126 22146
rect 26178 22094 26180 22146
rect 26124 21700 26180 22094
rect 26124 21634 26180 21644
rect 27244 22148 27300 22206
rect 27580 22148 27636 22316
rect 27804 22306 27860 22316
rect 27244 22092 27636 22148
rect 27692 22148 27748 22158
rect 27916 22148 27972 22988
rect 28924 23044 28980 23054
rect 28924 22950 28980 22988
rect 40012 22932 40068 22942
rect 40012 22838 40068 22876
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 40012 22482 40068 22494
rect 40012 22430 40014 22482
rect 40066 22430 40068 22482
rect 37660 22372 37716 22382
rect 37660 22278 37716 22316
rect 27692 22146 27972 22148
rect 27692 22094 27694 22146
rect 27746 22094 27972 22146
rect 27692 22092 27972 22094
rect 27020 20578 27076 20590
rect 27020 20526 27022 20578
rect 27074 20526 27076 20578
rect 27020 20188 27076 20526
rect 26124 20132 26180 20142
rect 26124 20018 26180 20076
rect 26124 19966 26126 20018
rect 26178 19966 26180 20018
rect 26124 19954 26180 19966
rect 26684 20132 27076 20188
rect 27244 20188 27300 22092
rect 27692 22082 27748 22092
rect 37884 21586 37940 21598
rect 37884 21534 37886 21586
rect 37938 21534 37940 21586
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 37660 20802 37716 20814
rect 37660 20750 37662 20802
rect 37714 20750 37716 20802
rect 27244 20132 27860 20188
rect 26684 20018 26740 20132
rect 27244 20066 27300 20076
rect 26684 19966 26686 20018
rect 26738 19966 26740 20018
rect 26124 19796 26180 19806
rect 26124 19702 26180 19740
rect 26236 19796 26292 19806
rect 26236 19794 26628 19796
rect 26236 19742 26238 19794
rect 26290 19742 26628 19794
rect 26236 19740 26628 19742
rect 26236 19730 26292 19740
rect 26236 19572 26292 19582
rect 26124 18450 26180 18462
rect 26124 18398 26126 18450
rect 26178 18398 26180 18450
rect 26124 18340 26180 18398
rect 26124 18274 26180 18284
rect 26236 18452 26292 19516
rect 26460 19460 26516 19470
rect 26460 19234 26516 19404
rect 26572 19458 26628 19740
rect 26572 19406 26574 19458
rect 26626 19406 26628 19458
rect 26572 19394 26628 19406
rect 26460 19182 26462 19234
rect 26514 19182 26516 19234
rect 26460 19170 26516 19182
rect 26572 19124 26628 19134
rect 26572 19030 26628 19068
rect 26572 18674 26628 18686
rect 26572 18622 26574 18674
rect 26626 18622 26628 18674
rect 26348 18452 26404 18462
rect 26236 18450 26404 18452
rect 26236 18398 26350 18450
rect 26402 18398 26404 18450
rect 26236 18396 26404 18398
rect 26012 18162 26068 18172
rect 25676 17042 25732 17052
rect 25788 16996 25844 17006
rect 26236 16996 26292 18396
rect 26348 18386 26404 18396
rect 26348 18228 26404 18238
rect 26348 18134 26404 18172
rect 25788 16994 26292 16996
rect 25788 16942 25790 16994
rect 25842 16942 26292 16994
rect 25788 16940 26292 16942
rect 26572 16996 26628 18622
rect 26684 18452 26740 19966
rect 27356 19906 27412 19918
rect 27356 19854 27358 19906
rect 27410 19854 27412 19906
rect 27356 19796 27412 19854
rect 27356 19730 27412 19740
rect 26908 18452 26964 18462
rect 26684 18450 26964 18452
rect 26684 18398 26910 18450
rect 26962 18398 26964 18450
rect 26684 18396 26964 18398
rect 25788 16930 25844 16940
rect 26572 16930 26628 16940
rect 25676 16884 25732 16894
rect 25676 16770 25732 16828
rect 25676 16718 25678 16770
rect 25730 16718 25732 16770
rect 25676 16706 25732 16718
rect 26348 16882 26404 16894
rect 26348 16830 26350 16882
rect 26402 16830 26404 16882
rect 25900 16210 25956 16222
rect 25900 16158 25902 16210
rect 25954 16158 25956 16210
rect 25900 16100 25956 16158
rect 25564 16044 25956 16100
rect 26348 15876 26404 16830
rect 26796 15876 26852 18396
rect 26908 18386 26964 18396
rect 27244 18340 27300 18350
rect 27244 17892 27300 18284
rect 27244 17798 27300 17836
rect 27692 18338 27748 18350
rect 27692 18286 27694 18338
rect 27746 18286 27748 18338
rect 27692 17778 27748 18286
rect 27692 17726 27694 17778
rect 27746 17726 27748 17778
rect 27692 17714 27748 17726
rect 27132 17666 27188 17678
rect 27132 17614 27134 17666
rect 27186 17614 27188 17666
rect 27020 16996 27076 17006
rect 27020 16902 27076 16940
rect 26348 15874 26852 15876
rect 26348 15822 26350 15874
rect 26402 15822 26798 15874
rect 26850 15822 26852 15874
rect 26348 15820 26852 15822
rect 26348 15764 26404 15820
rect 26796 15810 26852 15820
rect 25452 15708 26404 15764
rect 25228 15316 25284 15326
rect 25228 15222 25284 15260
rect 25452 15148 25508 15708
rect 23324 15092 23492 15148
rect 22540 14418 23156 14420
rect 22540 14366 22542 14418
rect 22594 14366 23156 14418
rect 22540 14364 23156 14366
rect 22540 14354 22596 14364
rect 22092 13918 22094 13970
rect 22146 13918 22148 13970
rect 22092 13906 22148 13918
rect 23436 13970 23492 15092
rect 23436 13918 23438 13970
rect 23490 13918 23492 13970
rect 23436 13906 23492 13918
rect 23772 15092 24052 15148
rect 25340 15092 25508 15148
rect 25676 15538 25732 15550
rect 25676 15486 25678 15538
rect 25730 15486 25732 15538
rect 25564 15092 25620 15102
rect 21644 13582 21646 13634
rect 21698 13582 21700 13634
rect 21644 13570 21700 13582
rect 23660 13858 23716 13870
rect 23660 13806 23662 13858
rect 23714 13806 23716 13858
rect 23660 13636 23716 13806
rect 23772 13858 23828 15092
rect 24668 14642 24724 14654
rect 24668 14590 24670 14642
rect 24722 14590 24724 14642
rect 24668 14532 24724 14590
rect 23772 13806 23774 13858
rect 23826 13806 23828 13858
rect 23772 13794 23828 13806
rect 24444 14476 24724 14532
rect 24780 14644 24836 14654
rect 24780 14532 24836 14588
rect 25004 14532 25060 14542
rect 25340 14532 25396 15092
rect 25564 14998 25620 15036
rect 25676 14644 25732 15486
rect 26012 15428 26068 15438
rect 26012 15334 26068 15372
rect 25788 15314 25844 15326
rect 25788 15262 25790 15314
rect 25842 15262 25844 15314
rect 25788 15148 25844 15262
rect 25788 15092 26404 15148
rect 25788 14644 25844 14654
rect 25676 14642 25844 14644
rect 25676 14590 25790 14642
rect 25842 14590 25844 14642
rect 25676 14588 25844 14590
rect 25788 14578 25844 14588
rect 24780 14530 25396 14532
rect 24780 14478 25006 14530
rect 25058 14478 25396 14530
rect 24780 14476 25396 14478
rect 24444 13636 24500 14476
rect 24668 13972 24724 13982
rect 24780 13972 24836 14476
rect 25004 14466 25060 14476
rect 24668 13970 24836 13972
rect 24668 13918 24670 13970
rect 24722 13918 24836 13970
rect 24668 13916 24836 13918
rect 25340 13970 25396 14476
rect 25340 13918 25342 13970
rect 25394 13918 25396 13970
rect 24668 13906 24724 13916
rect 25340 13906 25396 13918
rect 26348 13970 26404 15092
rect 27132 15092 27188 17614
rect 27804 17666 27860 20132
rect 30156 20132 30212 20142
rect 30156 20038 30212 20076
rect 29820 20020 29876 20030
rect 29484 19908 29540 19918
rect 29820 19908 29876 19964
rect 37660 20020 37716 20750
rect 37884 20132 37940 21534
rect 40012 21588 40068 22430
rect 40012 21522 40068 21532
rect 39900 21474 39956 21486
rect 39900 21422 39902 21474
rect 39954 21422 39956 21474
rect 39900 20916 39956 21422
rect 39900 20850 39956 20860
rect 40012 20914 40068 20926
rect 40012 20862 40014 20914
rect 40066 20862 40068 20914
rect 40012 20244 40068 20862
rect 40012 20178 40068 20188
rect 37884 20066 37940 20076
rect 37660 19954 37716 19964
rect 29484 19906 29876 19908
rect 29484 19854 29486 19906
rect 29538 19854 29876 19906
rect 29484 19852 29876 19854
rect 29484 19124 29540 19852
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 29484 19058 29540 19068
rect 37660 18452 37716 18462
rect 37660 18358 37716 18396
rect 29260 18340 29316 18350
rect 28252 18228 28308 18238
rect 28140 17892 28196 17902
rect 28140 17798 28196 17836
rect 28252 17778 28308 18172
rect 28252 17726 28254 17778
rect 28306 17726 28308 17778
rect 28252 17714 28308 17726
rect 29260 17778 29316 18284
rect 29820 18340 29876 18350
rect 29820 18246 29876 18284
rect 40012 18228 40068 18238
rect 40012 18134 40068 18172
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 29260 17726 29262 17778
rect 29314 17726 29316 17778
rect 29260 17714 29316 17726
rect 40012 17778 40068 17790
rect 40012 17726 40014 17778
rect 40066 17726 40068 17778
rect 27804 17614 27806 17666
rect 27858 17614 27860 17666
rect 27804 17602 27860 17614
rect 28476 17666 28532 17678
rect 28476 17614 28478 17666
rect 28530 17614 28532 17666
rect 27580 17556 27636 17566
rect 27580 17462 27636 17500
rect 28476 16884 28532 17614
rect 37660 17668 37716 17678
rect 37660 17574 37716 17612
rect 29148 17556 29204 17566
rect 29148 17462 29204 17500
rect 40012 17556 40068 17726
rect 40012 17490 40068 17500
rect 28476 16818 28532 16828
rect 29148 16884 29204 16894
rect 29148 16770 29204 16828
rect 37660 16884 37716 16894
rect 37660 16790 37716 16828
rect 40012 16884 40068 16894
rect 29148 16718 29150 16770
rect 29202 16718 29204 16770
rect 29148 16706 29204 16718
rect 40012 16770 40068 16828
rect 40012 16718 40014 16770
rect 40066 16718 40068 16770
rect 40012 16706 40068 16718
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 27132 15026 27188 15036
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 26348 13918 26350 13970
rect 26402 13918 26404 13970
rect 26348 13906 26404 13918
rect 27916 14642 27972 14654
rect 27916 14590 27918 14642
rect 27970 14590 27972 14642
rect 23660 13580 24500 13636
rect 18732 13022 18734 13074
rect 18786 13022 18788 13074
rect 18172 13010 18228 13020
rect 18732 13010 18788 13022
rect 15372 12910 15374 12962
rect 15426 12910 15428 12962
rect 15372 12898 15428 12910
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 24220 3668 24276 3678
rect 12348 3332 12404 3342
rect 12124 3330 12404 3332
rect 12124 3278 12350 3330
rect 12402 3278 12404 3330
rect 12124 3276 12404 3278
rect 12124 800 12180 3276
rect 12348 3266 12404 3276
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 24220 800 24276 3612
rect 24444 3556 24500 13580
rect 26460 13636 26516 13646
rect 26460 13542 26516 13580
rect 27132 13636 27188 13646
rect 27132 4338 27188 13580
rect 27916 13636 27972 14590
rect 27916 13570 27972 13580
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 27132 4286 27134 4338
rect 27186 4286 27188 4338
rect 27132 4274 27188 4286
rect 26908 4116 26964 4126
rect 25564 3668 25620 3678
rect 25564 3574 25620 3612
rect 24556 3556 24612 3566
rect 24444 3554 24612 3556
rect 24444 3502 24558 3554
rect 24610 3502 24612 3554
rect 24444 3500 24612 3502
rect 24556 3490 24612 3500
rect 26908 800 26964 4060
rect 28140 4116 28196 4126
rect 28140 4022 28196 4060
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 12096 0 12208 800
rect 24192 0 24304 800
rect 26880 0 26992 800
<< via2 >>
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 20188 38556 20244 38612
rect 20860 38220 20916 38276
rect 21420 38556 21476 38612
rect 16828 37436 16884 37492
rect 18396 37490 18452 37492
rect 18396 37438 18398 37490
rect 18398 37438 18450 37490
rect 18450 37438 18452 37490
rect 18396 37436 18452 37438
rect 16156 36652 16212 36708
rect 17388 36706 17444 36708
rect 17388 36654 17390 36706
rect 17390 36654 17442 36706
rect 17442 36654 17444 36706
rect 17388 36652 17444 36654
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 4172 26908 4228 26964
rect 1932 23548 1988 23604
rect 1932 22930 1988 22932
rect 1932 22878 1934 22930
rect 1934 22878 1986 22930
rect 1986 22878 1988 22930
rect 1932 22876 1988 22878
rect 13356 26290 13412 26292
rect 13356 26238 13358 26290
rect 13358 26238 13410 26290
rect 13410 26238 13412 26290
rect 13356 26236 13412 26238
rect 15148 26962 15204 26964
rect 15148 26910 15150 26962
rect 15150 26910 15202 26962
rect 15202 26910 15204 26962
rect 15148 26908 15204 26910
rect 14476 26236 14532 26292
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 14028 25676 14084 25732
rect 14924 25676 14980 25732
rect 16044 27858 16100 27860
rect 16044 27806 16046 27858
rect 16046 27806 16098 27858
rect 16098 27806 16100 27858
rect 16044 27804 16100 27806
rect 16156 26908 16212 26964
rect 16716 26908 16772 26964
rect 14476 25228 14532 25284
rect 15148 25004 15204 25060
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 4284 23938 4340 23940
rect 4284 23886 4286 23938
rect 4286 23886 4338 23938
rect 4338 23886 4340 23938
rect 4284 23884 4340 23886
rect 12012 23884 12068 23940
rect 4284 23154 4340 23156
rect 4284 23102 4286 23154
rect 4286 23102 4338 23154
rect 4338 23102 4340 23154
rect 4284 23100 4340 23102
rect 11340 23100 11396 23156
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 14700 23826 14756 23828
rect 14700 23774 14702 23826
rect 14702 23774 14754 23826
rect 14754 23774 14756 23826
rect 14700 23772 14756 23774
rect 14924 23436 14980 23492
rect 15260 23938 15316 23940
rect 15260 23886 15262 23938
rect 15262 23886 15314 23938
rect 15314 23886 15316 23938
rect 15260 23884 15316 23886
rect 15372 23714 15428 23716
rect 15372 23662 15374 23714
rect 15374 23662 15426 23714
rect 15426 23662 15428 23714
rect 15372 23660 15428 23662
rect 15148 23436 15204 23492
rect 16380 25282 16436 25284
rect 16380 25230 16382 25282
rect 16382 25230 16434 25282
rect 16434 25230 16436 25282
rect 16380 25228 16436 25230
rect 16268 24668 16324 24724
rect 15820 23436 15876 23492
rect 15036 23324 15092 23380
rect 15596 23378 15652 23380
rect 15596 23326 15598 23378
rect 15598 23326 15650 23378
rect 15650 23326 15652 23378
rect 15596 23324 15652 23326
rect 15260 23154 15316 23156
rect 15260 23102 15262 23154
rect 15262 23102 15314 23154
rect 15314 23102 15316 23154
rect 15260 23100 15316 23102
rect 15148 22988 15204 23044
rect 15932 23212 15988 23268
rect 15484 23154 15540 23156
rect 15484 23102 15486 23154
rect 15486 23102 15538 23154
rect 15538 23102 15540 23154
rect 15484 23100 15540 23102
rect 15148 22092 15204 22148
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 4284 20802 4340 20804
rect 4284 20750 4286 20802
rect 4286 20750 4338 20802
rect 4338 20750 4340 20802
rect 4284 20748 4340 20750
rect 12908 20860 12964 20916
rect 12124 20802 12180 20804
rect 12124 20750 12126 20802
rect 12126 20750 12178 20802
rect 12178 20750 12180 20802
rect 12124 20748 12180 20750
rect 15596 22092 15652 22148
rect 16268 23100 16324 23156
rect 16492 23660 16548 23716
rect 17500 26962 17556 26964
rect 17500 26910 17502 26962
rect 17502 26910 17554 26962
rect 17554 26910 17556 26962
rect 17500 26908 17556 26910
rect 17836 27804 17892 27860
rect 17836 27074 17892 27076
rect 17836 27022 17838 27074
rect 17838 27022 17890 27074
rect 17890 27022 17892 27074
rect 17836 27020 17892 27022
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 19292 27692 19348 27748
rect 19068 27074 19124 27076
rect 19068 27022 19070 27074
rect 19070 27022 19122 27074
rect 19122 27022 19124 27074
rect 19068 27020 19124 27022
rect 17836 25228 17892 25284
rect 22092 38274 22148 38276
rect 22092 38222 22094 38274
rect 22094 38222 22146 38274
rect 22146 38222 22148 38274
rect 22092 38220 22148 38222
rect 23548 38220 23604 38276
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 25564 38274 25620 38276
rect 25564 38222 25566 38274
rect 25566 38222 25618 38274
rect 25618 38222 25620 38274
rect 25564 38220 25620 38222
rect 24220 37436 24276 37492
rect 20300 27746 20356 27748
rect 20300 27694 20302 27746
rect 20302 27694 20354 27746
rect 20354 27694 20356 27746
rect 20300 27692 20356 27694
rect 26236 37490 26292 37492
rect 26236 37438 26238 37490
rect 26238 37438 26290 37490
rect 26290 37438 26292 37490
rect 26236 37436 26292 37438
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 23660 27692 23716 27748
rect 23436 27074 23492 27076
rect 23436 27022 23438 27074
rect 23438 27022 23490 27074
rect 23490 27022 23492 27074
rect 23436 27020 23492 27022
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 19852 24946 19908 24948
rect 19852 24894 19854 24946
rect 19854 24894 19906 24946
rect 19906 24894 19908 24946
rect 19852 24892 19908 24894
rect 20300 24892 20356 24948
rect 23324 26290 23380 26292
rect 23324 26238 23326 26290
rect 23326 26238 23378 26290
rect 23378 26238 23380 26290
rect 23324 26236 23380 26238
rect 20636 25228 20692 25284
rect 19964 24722 20020 24724
rect 19964 24670 19966 24722
rect 19966 24670 20018 24722
rect 20018 24670 20020 24722
rect 19964 24668 20020 24670
rect 21420 25282 21476 25284
rect 21420 25230 21422 25282
rect 21422 25230 21474 25282
rect 21474 25230 21476 25282
rect 21420 25228 21476 25230
rect 20748 24892 20804 24948
rect 16604 23548 16660 23604
rect 16828 23772 16884 23828
rect 16604 23212 16660 23268
rect 16380 23042 16436 23044
rect 16380 22990 16382 23042
rect 16382 22990 16434 23042
rect 16434 22990 16436 23042
rect 16380 22988 16436 22990
rect 15932 21756 15988 21812
rect 13692 20914 13748 20916
rect 13692 20862 13694 20914
rect 13694 20862 13746 20914
rect 13746 20862 13748 20914
rect 13692 20860 13748 20862
rect 14252 20748 14308 20804
rect 9996 20636 10052 20692
rect 14140 20636 14196 20692
rect 4172 20524 4228 20580
rect 1932 20188 1988 20244
rect 13468 20188 13524 20244
rect 14700 20636 14756 20692
rect 14252 20300 14308 20356
rect 14476 20300 14532 20356
rect 13692 20130 13748 20132
rect 13692 20078 13694 20130
rect 13694 20078 13746 20130
rect 13746 20078 13748 20130
rect 13692 20076 13748 20078
rect 14364 20076 14420 20132
rect 4284 20018 4340 20020
rect 4284 19966 4286 20018
rect 4286 19966 4338 20018
rect 4338 19966 4340 20018
rect 4284 19964 4340 19966
rect 13916 20018 13972 20020
rect 13916 19966 13918 20018
rect 13918 19966 13970 20018
rect 13970 19966 13972 20018
rect 13916 19964 13972 19966
rect 12124 19852 12180 19908
rect 1932 19794 1988 19796
rect 1932 19742 1934 19794
rect 1934 19742 1986 19794
rect 1986 19742 1988 19794
rect 1932 19740 1988 19742
rect 9996 19740 10052 19796
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 13468 19906 13524 19908
rect 13468 19854 13470 19906
rect 13470 19854 13522 19906
rect 13522 19854 13524 19906
rect 13468 19852 13524 19854
rect 14476 19404 14532 19460
rect 14812 20130 14868 20132
rect 14812 20078 14814 20130
rect 14814 20078 14866 20130
rect 14866 20078 14868 20130
rect 14812 20076 14868 20078
rect 12908 19234 12964 19236
rect 12908 19182 12910 19234
rect 12910 19182 12962 19234
rect 12962 19182 12964 19234
rect 12908 19180 12964 19182
rect 13580 19234 13636 19236
rect 13580 19182 13582 19234
rect 13582 19182 13634 19234
rect 13634 19182 13636 19234
rect 13580 19180 13636 19182
rect 14252 19180 14308 19236
rect 11452 18396 11508 18452
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 1932 17778 1988 17780
rect 1932 17726 1934 17778
rect 1934 17726 1986 17778
rect 1986 17726 1988 17778
rect 1932 17724 1988 17726
rect 4284 17666 4340 17668
rect 4284 17614 4286 17666
rect 4286 17614 4338 17666
rect 4338 17614 4340 17666
rect 4284 17612 4340 17614
rect 14140 18450 14196 18452
rect 14140 18398 14142 18450
rect 14142 18398 14194 18450
rect 14194 18398 14196 18450
rect 14140 18396 14196 18398
rect 14252 18172 14308 18228
rect 11452 17612 11508 17668
rect 15372 21644 15428 21700
rect 15484 21420 15540 21476
rect 15372 20300 15428 20356
rect 15708 20748 15764 20804
rect 15820 20076 15876 20132
rect 15260 19740 15316 19796
rect 15596 19906 15652 19908
rect 15596 19854 15598 19906
rect 15598 19854 15650 19906
rect 15650 19854 15652 19906
rect 15596 19852 15652 19854
rect 15260 19404 15316 19460
rect 15484 19404 15540 19460
rect 14476 18338 14532 18340
rect 14476 18286 14478 18338
rect 14478 18286 14530 18338
rect 14530 18286 14532 18338
rect 14476 18284 14532 18286
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 15932 21420 15988 21476
rect 15372 18396 15428 18452
rect 15820 18450 15876 18452
rect 15820 18398 15822 18450
rect 15822 18398 15874 18450
rect 15874 18398 15876 18450
rect 15820 18396 15876 18398
rect 15260 18226 15316 18228
rect 15260 18174 15262 18226
rect 15262 18174 15314 18226
rect 15314 18174 15316 18226
rect 15260 18172 15316 18174
rect 16156 21586 16212 21588
rect 16156 21534 16158 21586
rect 16158 21534 16210 21586
rect 16210 21534 16212 21586
rect 16156 21532 16212 21534
rect 16492 20748 16548 20804
rect 16268 20300 16324 20356
rect 16156 20076 16212 20132
rect 16940 23660 16996 23716
rect 17500 23548 17556 23604
rect 17276 23436 17332 23492
rect 17276 23212 17332 23268
rect 17612 21810 17668 21812
rect 17612 21758 17614 21810
rect 17614 21758 17666 21810
rect 17666 21758 17668 21810
rect 17612 21756 17668 21758
rect 17500 21644 17556 21700
rect 17276 21586 17332 21588
rect 17276 21534 17278 21586
rect 17278 21534 17330 21586
rect 17330 21534 17332 21586
rect 17276 21532 17332 21534
rect 16604 20188 16660 20244
rect 16716 20076 16772 20132
rect 16716 19180 16772 19236
rect 16044 18284 16100 18340
rect 15932 17554 15988 17556
rect 15932 17502 15934 17554
rect 15934 17502 15986 17554
rect 15986 17502 15988 17554
rect 15932 17500 15988 17502
rect 14812 17388 14868 17444
rect 16044 17388 16100 17444
rect 15820 16828 15876 16884
rect 17612 19122 17668 19124
rect 17612 19070 17614 19122
rect 17614 19070 17666 19122
rect 17666 19070 17668 19122
rect 17612 19068 17668 19070
rect 19516 23772 19572 23828
rect 18284 23714 18340 23716
rect 18284 23662 18286 23714
rect 18286 23662 18338 23714
rect 18338 23662 18340 23714
rect 18284 23660 18340 23662
rect 18508 22316 18564 22372
rect 18284 21698 18340 21700
rect 18284 21646 18286 21698
rect 18286 21646 18338 21698
rect 18338 21646 18340 21698
rect 18284 21644 18340 21646
rect 18508 21420 18564 21476
rect 18620 20242 18676 20244
rect 18620 20190 18622 20242
rect 18622 20190 18674 20242
rect 18674 20190 18676 20242
rect 18620 20188 18676 20190
rect 18284 20076 18340 20132
rect 18172 19458 18228 19460
rect 18172 19406 18174 19458
rect 18174 19406 18226 19458
rect 18226 19406 18228 19458
rect 18172 19404 18228 19406
rect 17948 19234 18004 19236
rect 17948 19182 17950 19234
rect 17950 19182 18002 19234
rect 18002 19182 18004 19234
rect 17948 19180 18004 19182
rect 17724 19010 17780 19012
rect 17724 18958 17726 19010
rect 17726 18958 17778 19010
rect 17778 18958 17780 19010
rect 17724 18956 17780 18958
rect 16828 18620 16884 18676
rect 18060 19068 18116 19124
rect 16716 17388 16772 17444
rect 16604 17052 16660 17108
rect 17276 17052 17332 17108
rect 16156 16268 16212 16324
rect 14364 15820 14420 15876
rect 15484 15874 15540 15876
rect 15484 15822 15486 15874
rect 15486 15822 15538 15874
rect 15538 15822 15540 15874
rect 15484 15820 15540 15822
rect 16716 16098 16772 16100
rect 16716 16046 16718 16098
rect 16718 16046 16770 16098
rect 16770 16046 16772 16098
rect 16716 16044 16772 16046
rect 16492 15484 16548 15540
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 18060 18396 18116 18452
rect 18172 18620 18228 18676
rect 18060 17052 18116 17108
rect 17276 16882 17332 16884
rect 17276 16830 17278 16882
rect 17278 16830 17330 16882
rect 17330 16830 17332 16882
rect 17276 16828 17332 16830
rect 17612 16994 17668 16996
rect 17612 16942 17614 16994
rect 17614 16942 17666 16994
rect 17666 16942 17668 16994
rect 17612 16940 17668 16942
rect 17500 16828 17556 16884
rect 17388 16716 17444 16772
rect 17276 16268 17332 16324
rect 17612 16098 17668 16100
rect 17612 16046 17614 16098
rect 17614 16046 17666 16098
rect 17666 16046 17668 16098
rect 17612 16044 17668 16046
rect 18284 18508 18340 18564
rect 19292 20076 19348 20132
rect 20300 23826 20356 23828
rect 20300 23774 20302 23826
rect 20302 23774 20354 23826
rect 20354 23774 20356 23826
rect 20300 23772 20356 23774
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 20188 23266 20244 23268
rect 20188 23214 20190 23266
rect 20190 23214 20242 23266
rect 20242 23214 20244 23266
rect 20188 23212 20244 23214
rect 20748 23212 20804 23268
rect 19740 22316 19796 22372
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 20188 21810 20244 21812
rect 20188 21758 20190 21810
rect 20190 21758 20242 21810
rect 20242 21758 20244 21810
rect 20188 21756 20244 21758
rect 20748 22428 20804 22484
rect 21196 24668 21252 24724
rect 20412 21586 20468 21588
rect 20412 21534 20414 21586
rect 20414 21534 20466 21586
rect 20466 21534 20468 21586
rect 20412 21532 20468 21534
rect 20188 20578 20244 20580
rect 20188 20526 20190 20578
rect 20190 20526 20242 20578
rect 20242 20526 20244 20578
rect 20188 20524 20244 20526
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 21868 24050 21924 24052
rect 21868 23998 21870 24050
rect 21870 23998 21922 24050
rect 21922 23998 21924 24050
rect 21868 23996 21924 23998
rect 22204 23996 22260 24052
rect 21644 23938 21700 23940
rect 21644 23886 21646 23938
rect 21646 23886 21698 23938
rect 21698 23886 21700 23938
rect 21644 23884 21700 23886
rect 22092 23772 22148 23828
rect 21420 22482 21476 22484
rect 21420 22430 21422 22482
rect 21422 22430 21474 22482
rect 21474 22430 21476 22482
rect 21420 22428 21476 22430
rect 21868 22370 21924 22372
rect 21868 22318 21870 22370
rect 21870 22318 21922 22370
rect 21922 22318 21924 22370
rect 21868 22316 21924 22318
rect 21420 21698 21476 21700
rect 21420 21646 21422 21698
rect 21422 21646 21474 21698
rect 21474 21646 21476 21698
rect 21420 21644 21476 21646
rect 19516 20076 19572 20132
rect 22092 21532 22148 21588
rect 21308 20524 21364 20580
rect 19180 19852 19236 19908
rect 18732 19794 18788 19796
rect 18732 19742 18734 19794
rect 18734 19742 18786 19794
rect 18786 19742 18788 19794
rect 18732 19740 18788 19742
rect 19068 19740 19124 19796
rect 18508 19234 18564 19236
rect 18508 19182 18510 19234
rect 18510 19182 18562 19234
rect 18562 19182 18564 19234
rect 18508 19180 18564 19182
rect 18956 19010 19012 19012
rect 18956 18958 18958 19010
rect 18958 18958 19010 19010
rect 19010 18958 19012 19010
rect 18956 18956 19012 18958
rect 18284 18172 18340 18228
rect 19628 19794 19684 19796
rect 19628 19742 19630 19794
rect 19630 19742 19682 19794
rect 19682 19742 19684 19794
rect 19628 19740 19684 19742
rect 19180 19234 19236 19236
rect 19180 19182 19182 19234
rect 19182 19182 19234 19234
rect 19234 19182 19236 19234
rect 19180 19180 19236 19182
rect 19404 19122 19460 19124
rect 19404 19070 19406 19122
rect 19406 19070 19458 19122
rect 19458 19070 19460 19122
rect 19404 19068 19460 19070
rect 18396 18060 18452 18116
rect 19292 17836 19348 17892
rect 19404 18396 19460 18452
rect 18956 17724 19012 17780
rect 18956 17500 19012 17556
rect 18172 16044 18228 16100
rect 13692 14588 13748 14644
rect 15372 14588 15428 14644
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 16716 14642 16772 14644
rect 16716 14590 16718 14642
rect 16718 14590 16770 14642
rect 16770 14590 16772 14642
rect 16716 14588 16772 14590
rect 16044 14252 16100 14308
rect 17388 15538 17444 15540
rect 17388 15486 17390 15538
rect 17390 15486 17442 15538
rect 17442 15486 17444 15538
rect 17388 15484 17444 15486
rect 17948 15314 18004 15316
rect 17948 15262 17950 15314
rect 17950 15262 18002 15314
rect 18002 15262 18004 15314
rect 17948 15260 18004 15262
rect 18620 16994 18676 16996
rect 18620 16942 18622 16994
rect 18622 16942 18674 16994
rect 18674 16942 18676 16994
rect 18620 16940 18676 16942
rect 18396 15260 18452 15316
rect 18508 16044 18564 16100
rect 19180 16828 19236 16884
rect 18732 14588 18788 14644
rect 17164 14252 17220 14308
rect 17612 14252 17668 14308
rect 19740 19404 19796 19460
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 20636 20076 20692 20132
rect 21756 20130 21812 20132
rect 21756 20078 21758 20130
rect 21758 20078 21810 20130
rect 21810 20078 21812 20130
rect 21756 20076 21812 20078
rect 20300 19234 20356 19236
rect 20300 19182 20302 19234
rect 20302 19182 20354 19234
rect 20354 19182 20356 19234
rect 20300 19180 20356 19182
rect 20524 19068 20580 19124
rect 20636 18732 20692 18788
rect 20524 18338 20580 18340
rect 20524 18286 20526 18338
rect 20526 18286 20578 18338
rect 20578 18286 20580 18338
rect 20524 18284 20580 18286
rect 20412 18060 20468 18116
rect 19628 17948 19684 18004
rect 20300 17948 20356 18004
rect 19852 17724 19908 17780
rect 20188 17442 20244 17444
rect 20188 17390 20190 17442
rect 20190 17390 20242 17442
rect 20242 17390 20244 17442
rect 20188 17388 20244 17390
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 19516 17106 19572 17108
rect 19516 17054 19518 17106
rect 19518 17054 19570 17106
rect 19570 17054 19572 17106
rect 19516 17052 19572 17054
rect 19740 16156 19796 16212
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 20188 15314 20244 15316
rect 20188 15262 20190 15314
rect 20190 15262 20242 15314
rect 20242 15262 20244 15314
rect 20188 15260 20244 15262
rect 20860 17948 20916 18004
rect 20972 18956 21028 19012
rect 20748 17778 20804 17780
rect 20748 17726 20750 17778
rect 20750 17726 20802 17778
rect 20802 17726 20804 17778
rect 20748 17724 20804 17726
rect 20636 16156 20692 16212
rect 20636 15538 20692 15540
rect 20636 15486 20638 15538
rect 20638 15486 20690 15538
rect 20690 15486 20692 15538
rect 20636 15484 20692 15486
rect 20748 15260 20804 15316
rect 20412 15036 20468 15092
rect 21980 19180 22036 19236
rect 21644 19010 21700 19012
rect 21644 18958 21646 19010
rect 21646 18958 21698 19010
rect 21698 18958 21700 19010
rect 21644 18956 21700 18958
rect 22876 24108 22932 24164
rect 22988 24556 23044 24612
rect 24332 27746 24388 27748
rect 24332 27694 24334 27746
rect 24334 27694 24386 27746
rect 24386 27694 24388 27746
rect 24332 27692 24388 27694
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 25228 27692 25284 27748
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 26908 27020 26964 27076
rect 23884 25282 23940 25284
rect 23884 25230 23886 25282
rect 23886 25230 23938 25282
rect 23938 25230 23940 25282
rect 23884 25228 23940 25230
rect 24556 26348 24612 26404
rect 25900 26514 25956 26516
rect 25900 26462 25902 26514
rect 25902 26462 25954 26514
rect 25954 26462 25956 26514
rect 25900 26460 25956 26462
rect 27580 27020 27636 27076
rect 28140 27074 28196 27076
rect 28140 27022 28142 27074
rect 28142 27022 28194 27074
rect 28194 27022 28196 27074
rect 28140 27020 28196 27022
rect 37660 27074 37716 27076
rect 37660 27022 37662 27074
rect 37662 27022 37714 27074
rect 37714 27022 37716 27074
rect 37660 27020 37716 27022
rect 28364 26962 28420 26964
rect 28364 26910 28366 26962
rect 28366 26910 28418 26962
rect 28418 26910 28420 26962
rect 28364 26908 28420 26910
rect 40012 27634 40068 27636
rect 40012 27582 40014 27634
rect 40014 27582 40066 27634
rect 40066 27582 40068 27634
rect 40012 27580 40068 27582
rect 37884 26908 37940 26964
rect 26908 26460 26964 26516
rect 25340 26402 25396 26404
rect 25340 26350 25342 26402
rect 25342 26350 25394 26402
rect 25394 26350 25396 26402
rect 25340 26348 25396 26350
rect 26012 26290 26068 26292
rect 26012 26238 26014 26290
rect 26014 26238 26066 26290
rect 26066 26238 26068 26290
rect 26012 26236 26068 26238
rect 39900 26796 39956 26852
rect 27132 26402 27188 26404
rect 27132 26350 27134 26402
rect 27134 26350 27186 26402
rect 27186 26350 27188 26402
rect 27132 26348 27188 26350
rect 37660 26290 37716 26292
rect 37660 26238 37662 26290
rect 37662 26238 37714 26290
rect 37714 26238 37716 26290
rect 37660 26236 37716 26238
rect 40012 26236 40068 26292
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 25116 25228 25172 25284
rect 23660 24610 23716 24612
rect 23660 24558 23662 24610
rect 23662 24558 23714 24610
rect 23714 24558 23716 24610
rect 23660 24556 23716 24558
rect 22540 23884 22596 23940
rect 22316 23826 22372 23828
rect 22316 23774 22318 23826
rect 22318 23774 22370 23826
rect 22370 23774 22372 23826
rect 22316 23772 22372 23774
rect 22428 22428 22484 22484
rect 23772 24108 23828 24164
rect 23436 23938 23492 23940
rect 23436 23886 23438 23938
rect 23438 23886 23490 23938
rect 23490 23886 23492 23938
rect 23436 23884 23492 23886
rect 23100 20130 23156 20132
rect 23100 20078 23102 20130
rect 23102 20078 23154 20130
rect 23154 20078 23156 20130
rect 23100 20076 23156 20078
rect 22316 19122 22372 19124
rect 22316 19070 22318 19122
rect 22318 19070 22370 19122
rect 22370 19070 22372 19122
rect 22316 19068 22372 19070
rect 22540 18732 22596 18788
rect 21980 18284 22036 18340
rect 21308 16210 21364 16212
rect 21308 16158 21310 16210
rect 21310 16158 21362 16210
rect 21362 16158 21364 16210
rect 21308 16156 21364 16158
rect 21084 15036 21140 15092
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 22092 15314 22148 15316
rect 22092 15262 22094 15314
rect 22094 15262 22146 15314
rect 22146 15262 22148 15314
rect 22092 15260 22148 15262
rect 23660 23100 23716 23156
rect 23884 23714 23940 23716
rect 23884 23662 23886 23714
rect 23886 23662 23938 23714
rect 23938 23662 23940 23714
rect 23884 23660 23940 23662
rect 23996 22540 24052 22596
rect 24108 23772 24164 23828
rect 23884 21756 23940 21812
rect 23660 21586 23716 21588
rect 23660 21534 23662 21586
rect 23662 21534 23714 21586
rect 23714 21534 23716 21586
rect 23660 21532 23716 21534
rect 24332 24108 24388 24164
rect 24444 23996 24500 24052
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 24220 23548 24276 23604
rect 24556 23548 24612 23604
rect 25228 23548 25284 23604
rect 23996 21644 24052 21700
rect 23548 20130 23604 20132
rect 23548 20078 23550 20130
rect 23550 20078 23602 20130
rect 23602 20078 23604 20130
rect 23548 20076 23604 20078
rect 23884 19516 23940 19572
rect 23212 19404 23268 19460
rect 27132 23996 27188 24052
rect 26348 23660 26404 23716
rect 25452 22428 25508 22484
rect 24668 20130 24724 20132
rect 24668 20078 24670 20130
rect 24670 20078 24722 20130
rect 24722 20078 24724 20130
rect 24668 20076 24724 20078
rect 24332 19234 24388 19236
rect 24332 19182 24334 19234
rect 24334 19182 24386 19234
rect 24386 19182 24388 19234
rect 24332 19180 24388 19182
rect 24220 19122 24276 19124
rect 24220 19070 24222 19122
rect 24222 19070 24274 19122
rect 24274 19070 24276 19122
rect 24220 19068 24276 19070
rect 23436 18284 23492 18340
rect 23100 17948 23156 18004
rect 23436 17836 23492 17892
rect 26908 22540 26964 22596
rect 25340 19516 25396 19572
rect 25676 19906 25732 19908
rect 25676 19854 25678 19906
rect 25678 19854 25730 19906
rect 25730 19854 25732 19906
rect 25676 19852 25732 19854
rect 25900 19068 25956 19124
rect 23996 16828 24052 16884
rect 25228 17388 25284 17444
rect 23996 16604 24052 16660
rect 22876 15484 22932 15540
rect 22764 15314 22820 15316
rect 22764 15262 22766 15314
rect 22766 15262 22818 15314
rect 22818 15262 22820 15314
rect 22764 15260 22820 15262
rect 21868 14588 21924 14644
rect 22988 14588 23044 14644
rect 25340 16604 25396 16660
rect 25340 15372 25396 15428
rect 25564 17612 25620 17668
rect 26348 22370 26404 22372
rect 26348 22318 26350 22370
rect 26350 22318 26402 22370
rect 26402 22318 26404 22370
rect 26348 22316 26404 22318
rect 28476 24050 28532 24052
rect 28476 23998 28478 24050
rect 28478 23998 28530 24050
rect 28530 23998 28532 24050
rect 28476 23996 28532 23998
rect 37660 23938 37716 23940
rect 37660 23886 37662 23938
rect 37662 23886 37714 23938
rect 37714 23886 37716 23938
rect 37660 23884 37716 23886
rect 40012 23548 40068 23604
rect 37660 23154 37716 23156
rect 37660 23102 37662 23154
rect 37662 23102 37714 23154
rect 37714 23102 37716 23154
rect 37660 23100 37716 23102
rect 27916 22988 27972 23044
rect 27468 22370 27524 22372
rect 27468 22318 27470 22370
rect 27470 22318 27522 22370
rect 27522 22318 27524 22370
rect 27468 22316 27524 22318
rect 26124 21644 26180 21700
rect 28924 23042 28980 23044
rect 28924 22990 28926 23042
rect 28926 22990 28978 23042
rect 28978 22990 28980 23042
rect 28924 22988 28980 22990
rect 40012 22930 40068 22932
rect 40012 22878 40014 22930
rect 40014 22878 40066 22930
rect 40066 22878 40068 22930
rect 40012 22876 40068 22878
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 37660 22370 37716 22372
rect 37660 22318 37662 22370
rect 37662 22318 37714 22370
rect 37714 22318 37716 22370
rect 37660 22316 37716 22318
rect 26124 20076 26180 20132
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 27244 20076 27300 20132
rect 26124 19794 26180 19796
rect 26124 19742 26126 19794
rect 26126 19742 26178 19794
rect 26178 19742 26180 19794
rect 26124 19740 26180 19742
rect 26236 19516 26292 19572
rect 26124 18284 26180 18340
rect 26460 19404 26516 19460
rect 26572 19122 26628 19124
rect 26572 19070 26574 19122
rect 26574 19070 26626 19122
rect 26626 19070 26628 19122
rect 26572 19068 26628 19070
rect 26012 18172 26068 18228
rect 25676 17052 25732 17108
rect 26348 18226 26404 18228
rect 26348 18174 26350 18226
rect 26350 18174 26402 18226
rect 26402 18174 26404 18226
rect 26348 18172 26404 18174
rect 27356 19740 27412 19796
rect 26572 16940 26628 16996
rect 25676 16828 25732 16884
rect 27244 18284 27300 18340
rect 27244 17890 27300 17892
rect 27244 17838 27246 17890
rect 27246 17838 27298 17890
rect 27298 17838 27300 17890
rect 27244 17836 27300 17838
rect 27020 16994 27076 16996
rect 27020 16942 27022 16994
rect 27022 16942 27074 16994
rect 27074 16942 27076 16994
rect 27020 16940 27076 16942
rect 25228 15314 25284 15316
rect 25228 15262 25230 15314
rect 25230 15262 25282 15314
rect 25282 15262 25284 15314
rect 25228 15260 25284 15262
rect 24780 14588 24836 14644
rect 25564 15090 25620 15092
rect 25564 15038 25566 15090
rect 25566 15038 25618 15090
rect 25618 15038 25620 15090
rect 25564 15036 25620 15038
rect 26012 15426 26068 15428
rect 26012 15374 26014 15426
rect 26014 15374 26066 15426
rect 26066 15374 26068 15426
rect 26012 15372 26068 15374
rect 30156 20130 30212 20132
rect 30156 20078 30158 20130
rect 30158 20078 30210 20130
rect 30210 20078 30212 20130
rect 30156 20076 30212 20078
rect 29820 20018 29876 20020
rect 29820 19966 29822 20018
rect 29822 19966 29874 20018
rect 29874 19966 29876 20018
rect 29820 19964 29876 19966
rect 40012 21532 40068 21588
rect 39900 20860 39956 20916
rect 40012 20188 40068 20244
rect 37884 20076 37940 20132
rect 37660 19964 37716 20020
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 29484 19068 29540 19124
rect 37660 18450 37716 18452
rect 37660 18398 37662 18450
rect 37662 18398 37714 18450
rect 37714 18398 37716 18450
rect 37660 18396 37716 18398
rect 29260 18284 29316 18340
rect 28252 18172 28308 18228
rect 28140 17890 28196 17892
rect 28140 17838 28142 17890
rect 28142 17838 28194 17890
rect 28194 17838 28196 17890
rect 28140 17836 28196 17838
rect 29820 18338 29876 18340
rect 29820 18286 29822 18338
rect 29822 18286 29874 18338
rect 29874 18286 29876 18338
rect 29820 18284 29876 18286
rect 40012 18226 40068 18228
rect 40012 18174 40014 18226
rect 40014 18174 40066 18226
rect 40066 18174 40068 18226
rect 40012 18172 40068 18174
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 27580 17554 27636 17556
rect 27580 17502 27582 17554
rect 27582 17502 27634 17554
rect 27634 17502 27636 17554
rect 27580 17500 27636 17502
rect 37660 17666 37716 17668
rect 37660 17614 37662 17666
rect 37662 17614 37714 17666
rect 37714 17614 37716 17666
rect 37660 17612 37716 17614
rect 29148 17554 29204 17556
rect 29148 17502 29150 17554
rect 29150 17502 29202 17554
rect 29202 17502 29204 17554
rect 29148 17500 29204 17502
rect 40012 17500 40068 17556
rect 28476 16828 28532 16884
rect 29148 16828 29204 16884
rect 37660 16882 37716 16884
rect 37660 16830 37662 16882
rect 37662 16830 37714 16882
rect 37714 16830 37716 16882
rect 37660 16828 37716 16830
rect 40012 16828 40068 16884
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 27132 15036 27188 15092
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 24220 3612 24276 3668
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 26460 13634 26516 13636
rect 26460 13582 26462 13634
rect 26462 13582 26514 13634
rect 26514 13582 26516 13634
rect 26460 13580 26516 13582
rect 27132 13580 27188 13636
rect 27916 13580 27972 13636
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 26908 4060 26964 4116
rect 25564 3666 25620 3668
rect 25564 3614 25566 3666
rect 25566 3614 25618 3666
rect 25618 3614 25620 3666
rect 25564 3612 25620 3614
rect 28140 4114 28196 4116
rect 28140 4062 28142 4114
rect 28142 4062 28194 4114
rect 28194 4062 28196 4114
rect 28140 4060 28196 4062
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
<< metal3 >>
rect 20178 38556 20188 38612
rect 20244 38556 21420 38612
rect 21476 38556 21486 38612
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 20850 38220 20860 38276
rect 20916 38220 22092 38276
rect 22148 38220 22158 38276
rect 23538 38220 23548 38276
rect 23604 38220 25564 38276
rect 25620 38220 25630 38276
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 16818 37436 16828 37492
rect 16884 37436 18396 37492
rect 18452 37436 18462 37492
rect 24210 37436 24220 37492
rect 24276 37436 26236 37492
rect 26292 37436 26302 37492
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 16146 36652 16156 36708
rect 16212 36652 17388 36708
rect 17444 36652 17454 36708
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 16034 27804 16044 27860
rect 16100 27804 17836 27860
rect 17892 27804 17902 27860
rect 19282 27692 19292 27748
rect 19348 27692 20300 27748
rect 20356 27692 20366 27748
rect 23650 27692 23660 27748
rect 23716 27692 24332 27748
rect 24388 27692 25228 27748
rect 25284 27692 25294 27748
rect 41200 27636 42000 27664
rect 40002 27580 40012 27636
rect 40068 27580 42000 27636
rect 41200 27552 42000 27580
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 17826 27020 17836 27076
rect 17892 27020 19068 27076
rect 19124 27020 23436 27076
rect 23492 27020 23502 27076
rect 26898 27020 26908 27076
rect 26964 27020 27580 27076
rect 27636 27020 28140 27076
rect 28196 27020 37660 27076
rect 37716 27020 37726 27076
rect 0 26964 800 26992
rect 41200 26964 42000 26992
rect 0 26908 4172 26964
rect 4228 26908 4238 26964
rect 15138 26908 15148 26964
rect 15204 26908 16156 26964
rect 16212 26908 16222 26964
rect 16706 26908 16716 26964
rect 16772 26908 17500 26964
rect 17556 26908 17566 26964
rect 28354 26908 28364 26964
rect 28420 26908 37884 26964
rect 37940 26908 37950 26964
rect 39900 26908 42000 26964
rect 0 26880 800 26908
rect 39900 26852 39956 26908
rect 41200 26880 42000 26908
rect 39890 26796 39900 26852
rect 39956 26796 39966 26852
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 25890 26460 25900 26516
rect 25956 26460 26908 26516
rect 26964 26460 26974 26516
rect 24546 26348 24556 26404
rect 24612 26348 25340 26404
rect 25396 26348 25406 26404
rect 27122 26348 27132 26404
rect 27188 26348 31948 26404
rect 31892 26292 31948 26348
rect 41200 26292 42000 26320
rect 13346 26236 13356 26292
rect 13412 26236 14476 26292
rect 14532 26236 14542 26292
rect 23314 26236 23324 26292
rect 23380 26236 26012 26292
rect 26068 26236 26078 26292
rect 31892 26236 37660 26292
rect 37716 26236 37726 26292
rect 40002 26236 40012 26292
rect 40068 26236 42000 26292
rect 41200 26208 42000 26236
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 14018 25676 14028 25732
rect 14084 25676 14924 25732
rect 14980 25676 14990 25732
rect 14466 25228 14476 25284
rect 14532 25228 16380 25284
rect 16436 25228 17836 25284
rect 17892 25228 17902 25284
rect 20626 25228 20636 25284
rect 20692 25228 21420 25284
rect 21476 25228 23884 25284
rect 23940 25228 25116 25284
rect 25172 25228 25182 25284
rect 15148 25060 15204 25228
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 15138 25004 15148 25060
rect 15204 25004 15214 25060
rect 19842 24892 19852 24948
rect 19908 24892 20300 24948
rect 20356 24892 20748 24948
rect 20804 24892 20814 24948
rect 16258 24668 16268 24724
rect 16324 24668 19964 24724
rect 20020 24668 21196 24724
rect 21252 24668 21262 24724
rect 22978 24556 22988 24612
rect 23044 24556 23660 24612
rect 23716 24556 23726 24612
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 22866 24108 22876 24164
rect 22932 24108 23772 24164
rect 23828 24108 24332 24164
rect 24388 24108 24398 24164
rect 21858 23996 21868 24052
rect 21924 23996 22204 24052
rect 22260 23996 24444 24052
rect 24500 23996 24510 24052
rect 27122 23996 27132 24052
rect 27188 23996 28476 24052
rect 28532 23996 31948 24052
rect 31892 23940 31948 23996
rect 4274 23884 4284 23940
rect 4340 23884 12012 23940
rect 12068 23884 15260 23940
rect 15316 23884 15326 23940
rect 21634 23884 21644 23940
rect 21700 23884 22540 23940
rect 22596 23884 23436 23940
rect 23492 23884 23502 23940
rect 31892 23884 37660 23940
rect 37716 23884 37726 23940
rect 14690 23772 14700 23828
rect 14756 23772 16828 23828
rect 16884 23772 19516 23828
rect 19572 23772 20300 23828
rect 20356 23772 22092 23828
rect 22148 23772 22158 23828
rect 22306 23772 22316 23828
rect 22372 23772 24108 23828
rect 24164 23772 24174 23828
rect 15362 23660 15372 23716
rect 15428 23660 16492 23716
rect 16548 23660 16558 23716
rect 16930 23660 16940 23716
rect 16996 23660 18284 23716
rect 18340 23660 21924 23716
rect 23874 23660 23884 23716
rect 23940 23660 26348 23716
rect 26404 23660 26414 23716
rect 0 23604 800 23632
rect 21868 23604 21924 23660
rect 41200 23604 42000 23632
rect 0 23548 1932 23604
rect 1988 23548 1998 23604
rect 16594 23548 16604 23604
rect 16660 23548 17500 23604
rect 17556 23548 17566 23604
rect 21868 23548 24220 23604
rect 24276 23548 24556 23604
rect 24612 23548 25228 23604
rect 25284 23548 25294 23604
rect 40002 23548 40012 23604
rect 40068 23548 42000 23604
rect 0 23520 800 23548
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 41200 23520 42000 23548
rect 14914 23436 14924 23492
rect 14980 23436 15148 23492
rect 15204 23436 15820 23492
rect 15876 23436 17276 23492
rect 17332 23436 17342 23492
rect 15026 23324 15036 23380
rect 15092 23324 15596 23380
rect 15652 23324 15662 23380
rect 15922 23212 15932 23268
rect 15988 23212 16604 23268
rect 16660 23212 17108 23268
rect 17266 23212 17276 23268
rect 17332 23212 20188 23268
rect 20244 23212 20748 23268
rect 20804 23212 20814 23268
rect 17052 23156 17108 23212
rect 4274 23100 4284 23156
rect 4340 23100 11340 23156
rect 11396 23100 15260 23156
rect 15316 23100 15326 23156
rect 15474 23100 15484 23156
rect 15540 23100 16268 23156
rect 16324 23100 16334 23156
rect 17052 23100 23660 23156
rect 23716 23100 23726 23156
rect 31892 23100 37660 23156
rect 37716 23100 37726 23156
rect 31892 23044 31948 23100
rect 15138 22988 15148 23044
rect 15204 22988 16380 23044
rect 16436 22988 16446 23044
rect 27906 22988 27916 23044
rect 27972 22988 28924 23044
rect 28980 22988 31948 23044
rect 0 22932 800 22960
rect 41200 22932 42000 22960
rect 0 22876 1932 22932
rect 1988 22876 1998 22932
rect 40002 22876 40012 22932
rect 40068 22876 42000 22932
rect 0 22848 800 22876
rect 41200 22848 42000 22876
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 23986 22540 23996 22596
rect 24052 22540 26908 22596
rect 26964 22540 26974 22596
rect 20738 22428 20748 22484
rect 20804 22428 21420 22484
rect 21476 22428 22428 22484
rect 22484 22428 22494 22484
rect 25442 22428 25452 22484
rect 25508 22428 31948 22484
rect 31892 22372 31948 22428
rect 18498 22316 18508 22372
rect 18564 22316 19740 22372
rect 19796 22316 21868 22372
rect 21924 22316 21934 22372
rect 26338 22316 26348 22372
rect 26404 22316 27468 22372
rect 27524 22316 27534 22372
rect 31892 22316 37660 22372
rect 37716 22316 37726 22372
rect 15138 22092 15148 22148
rect 15204 22092 15596 22148
rect 15652 22092 15662 22148
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 15922 21756 15932 21812
rect 15988 21756 17612 21812
rect 17668 21756 17678 21812
rect 20178 21756 20188 21812
rect 20244 21756 23884 21812
rect 23940 21756 23950 21812
rect 15932 21700 15988 21756
rect 15362 21644 15372 21700
rect 15428 21644 15988 21700
rect 17490 21644 17500 21700
rect 17556 21644 18284 21700
rect 18340 21644 18350 21700
rect 21410 21644 21420 21700
rect 21476 21644 23996 21700
rect 24052 21644 26124 21700
rect 26180 21644 26190 21700
rect 41200 21588 42000 21616
rect 16146 21532 16156 21588
rect 16212 21532 17276 21588
rect 17332 21532 20412 21588
rect 20468 21532 20478 21588
rect 22082 21532 22092 21588
rect 22148 21532 23660 21588
rect 23716 21532 23726 21588
rect 40002 21532 40012 21588
rect 40068 21532 42000 21588
rect 41200 21504 42000 21532
rect 15474 21420 15484 21476
rect 15540 21420 15932 21476
rect 15988 21420 18508 21476
rect 18564 21420 18574 21476
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 41200 20916 42000 20944
rect 12898 20860 12908 20916
rect 12964 20860 13692 20916
rect 13748 20860 13758 20916
rect 39890 20860 39900 20916
rect 39956 20860 42000 20916
rect 41200 20832 42000 20860
rect 4274 20748 4284 20804
rect 4340 20748 8428 20804
rect 12114 20748 12124 20804
rect 12180 20748 14252 20804
rect 14308 20748 14318 20804
rect 15092 20748 15708 20804
rect 15764 20748 16492 20804
rect 16548 20748 16558 20804
rect 8372 20692 8428 20748
rect 15092 20692 15148 20748
rect 8372 20636 9996 20692
rect 10052 20636 14140 20692
rect 14196 20636 14206 20692
rect 14690 20636 14700 20692
rect 14756 20636 15148 20692
rect 4162 20524 4172 20580
rect 4228 20524 20188 20580
rect 20244 20524 21308 20580
rect 21364 20524 21374 20580
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 14242 20300 14252 20356
rect 14308 20300 14318 20356
rect 14466 20300 14476 20356
rect 14532 20300 15372 20356
rect 15428 20300 16268 20356
rect 16324 20300 16334 20356
rect 0 20244 800 20272
rect 14252 20244 14308 20300
rect 41200 20244 42000 20272
rect 0 20188 1932 20244
rect 1988 20188 1998 20244
rect 13458 20188 13468 20244
rect 13524 20188 16604 20244
rect 16660 20188 16670 20244
rect 18060 20188 18620 20244
rect 18676 20188 18686 20244
rect 40002 20188 40012 20244
rect 40068 20188 42000 20244
rect 0 20160 800 20188
rect 18060 20132 18116 20188
rect 41200 20160 42000 20188
rect 13682 20076 13692 20132
rect 13748 20076 14364 20132
rect 14420 20076 14430 20132
rect 14802 20076 14812 20132
rect 14868 20076 15820 20132
rect 15876 20076 15886 20132
rect 16146 20076 16156 20132
rect 16212 20076 16716 20132
rect 16772 20076 18116 20132
rect 18274 20076 18284 20132
rect 18340 20076 19292 20132
rect 19348 20076 19358 20132
rect 19506 20076 19516 20132
rect 19572 20076 19610 20132
rect 20626 20076 20636 20132
rect 20692 20076 21756 20132
rect 21812 20076 23100 20132
rect 23156 20076 23548 20132
rect 23604 20076 23614 20132
rect 24658 20076 24668 20132
rect 24724 20076 26124 20132
rect 26180 20076 27244 20132
rect 27300 20076 27310 20132
rect 30146 20076 30156 20132
rect 30212 20076 37884 20132
rect 37940 20076 37950 20132
rect 4274 19964 4284 20020
rect 4340 19964 8428 20020
rect 13906 19964 13916 20020
rect 13972 19964 15148 20020
rect 29810 19964 29820 20020
rect 29876 19964 37660 20020
rect 37716 19964 37726 20020
rect 8372 19796 8428 19964
rect 15092 19908 15148 19964
rect 12114 19852 12124 19908
rect 12180 19852 13468 19908
rect 13524 19852 13534 19908
rect 15092 19852 15596 19908
rect 15652 19852 15662 19908
rect 19170 19852 19180 19908
rect 19236 19852 25676 19908
rect 25732 19852 25742 19908
rect 1922 19740 1932 19796
rect 1988 19740 1998 19796
rect 8372 19740 9996 19796
rect 10052 19740 15260 19796
rect 15316 19740 15326 19796
rect 18722 19740 18732 19796
rect 18788 19740 19068 19796
rect 19124 19740 19628 19796
rect 19684 19740 19694 19796
rect 26114 19740 26124 19796
rect 26180 19740 27356 19796
rect 27412 19740 27422 19796
rect 0 19572 800 19600
rect 1932 19572 1988 19740
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 0 19516 1988 19572
rect 23874 19516 23884 19572
rect 23940 19516 25340 19572
rect 25396 19516 26236 19572
rect 26292 19516 26302 19572
rect 0 19488 800 19516
rect 14466 19404 14476 19460
rect 14532 19404 15260 19460
rect 15316 19404 15326 19460
rect 15474 19404 15484 19460
rect 15540 19404 18172 19460
rect 18228 19404 19740 19460
rect 19796 19404 19806 19460
rect 23202 19404 23212 19460
rect 23268 19404 26460 19460
rect 26516 19404 26526 19460
rect 15092 19236 15148 19404
rect 12898 19180 12908 19236
rect 12964 19180 13580 19236
rect 13636 19180 14252 19236
rect 14308 19180 14318 19236
rect 15092 19180 16716 19236
rect 16772 19180 16782 19236
rect 17938 19180 17948 19236
rect 18004 19180 18508 19236
rect 18564 19180 18574 19236
rect 19170 19180 19180 19236
rect 19236 19180 20300 19236
rect 20356 19180 21980 19236
rect 22036 19180 24332 19236
rect 24388 19180 24398 19236
rect 17602 19068 17612 19124
rect 17668 19068 18060 19124
rect 18116 19068 19404 19124
rect 19460 19068 19470 19124
rect 20514 19068 20524 19124
rect 20580 19068 22316 19124
rect 22372 19068 22382 19124
rect 24210 19068 24220 19124
rect 24276 19068 25900 19124
rect 25956 19068 25966 19124
rect 26562 19068 26572 19124
rect 26628 19068 29484 19124
rect 29540 19068 29550 19124
rect 17714 18956 17724 19012
rect 17780 18956 18956 19012
rect 19012 18956 19022 19012
rect 20962 18956 20972 19012
rect 21028 18956 21644 19012
rect 21700 18956 21710 19012
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 20626 18732 20636 18788
rect 20692 18732 22540 18788
rect 22596 18732 22606 18788
rect 16818 18620 16828 18676
rect 16884 18620 18172 18676
rect 18228 18620 18238 18676
rect 18274 18508 18284 18564
rect 18340 18508 18350 18564
rect 18284 18452 18340 18508
rect 11442 18396 11452 18452
rect 11508 18396 14140 18452
rect 14196 18396 14206 18452
rect 15362 18396 15372 18452
rect 15428 18396 15820 18452
rect 15876 18396 18060 18452
rect 18116 18396 18126 18452
rect 18284 18396 19404 18452
rect 19460 18396 19470 18452
rect 31892 18396 37660 18452
rect 37716 18396 37726 18452
rect 31892 18340 31948 18396
rect 14466 18284 14476 18340
rect 14532 18284 15876 18340
rect 16034 18284 16044 18340
rect 16100 18284 20524 18340
rect 20580 18284 21980 18340
rect 22036 18284 22046 18340
rect 23426 18284 23436 18340
rect 23492 18284 26124 18340
rect 26180 18284 27244 18340
rect 27300 18284 27310 18340
rect 29250 18284 29260 18340
rect 29316 18284 29820 18340
rect 29876 18284 31948 18340
rect 15820 18228 15876 18284
rect 41200 18228 42000 18256
rect 14242 18172 14252 18228
rect 14308 18172 15260 18228
rect 15316 18172 15326 18228
rect 15820 18172 18284 18228
rect 18340 18172 26012 18228
rect 26068 18172 26078 18228
rect 26338 18172 26348 18228
rect 26404 18172 28252 18228
rect 28308 18172 28318 18228
rect 40002 18172 40012 18228
rect 40068 18172 42000 18228
rect 41200 18144 42000 18172
rect 18386 18060 18396 18116
rect 18452 18060 20412 18116
rect 20468 18060 20478 18116
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 19618 17948 19628 18004
rect 19684 17948 20300 18004
rect 20356 17948 20860 18004
rect 20916 17948 23100 18004
rect 23156 17948 23166 18004
rect 19282 17836 19292 17892
rect 19348 17836 23436 17892
rect 23492 17836 23502 17892
rect 27234 17836 27244 17892
rect 27300 17836 28140 17892
rect 28196 17836 28206 17892
rect 1922 17724 1932 17780
rect 1988 17724 1998 17780
rect 18946 17724 18956 17780
rect 19012 17724 19852 17780
rect 19908 17724 20748 17780
rect 20804 17724 20814 17780
rect 0 17556 800 17584
rect 1932 17556 1988 17724
rect 4274 17612 4284 17668
rect 4340 17612 11452 17668
rect 11508 17612 11518 17668
rect 25554 17612 25564 17668
rect 25620 17612 37660 17668
rect 37716 17612 37726 17668
rect 41200 17556 42000 17584
rect 0 17500 1988 17556
rect 15922 17500 15932 17556
rect 15988 17500 18956 17556
rect 19012 17500 19022 17556
rect 27570 17500 27580 17556
rect 27636 17500 29148 17556
rect 29204 17500 29214 17556
rect 40002 17500 40012 17556
rect 40068 17500 42000 17556
rect 0 17472 800 17500
rect 41200 17472 42000 17500
rect 14802 17388 14812 17444
rect 14868 17388 16044 17444
rect 16100 17388 16110 17444
rect 16706 17388 16716 17444
rect 16772 17388 20188 17444
rect 20244 17388 25228 17444
rect 25284 17388 25294 17444
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 16594 17052 16604 17108
rect 16660 17052 17276 17108
rect 17332 17052 18060 17108
rect 18116 17052 18126 17108
rect 19478 17052 19516 17108
rect 19572 17052 19582 17108
rect 25666 17052 25676 17108
rect 25732 17052 25956 17108
rect 17602 16940 17612 16996
rect 17668 16940 18620 16996
rect 18676 16940 18686 16996
rect 15810 16828 15820 16884
rect 15876 16828 17276 16884
rect 17332 16828 17342 16884
rect 17490 16828 17500 16884
rect 17556 16828 19180 16884
rect 19236 16828 19246 16884
rect 23986 16828 23996 16884
rect 24052 16828 25676 16884
rect 25732 16828 25742 16884
rect 25900 16772 25956 17052
rect 26562 16940 26572 16996
rect 26628 16940 27020 16996
rect 27076 16940 27086 16996
rect 41200 16884 42000 16912
rect 28466 16828 28476 16884
rect 28532 16828 29148 16884
rect 29204 16828 37660 16884
rect 37716 16828 37726 16884
rect 40002 16828 40012 16884
rect 40068 16828 42000 16884
rect 41200 16800 42000 16828
rect 17378 16716 17388 16772
rect 17444 16716 25956 16772
rect 23986 16604 23996 16660
rect 24052 16604 25340 16660
rect 25396 16604 25406 16660
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 16146 16268 16156 16324
rect 16212 16268 17276 16324
rect 17332 16268 17342 16324
rect 19730 16156 19740 16212
rect 19796 16156 20636 16212
rect 20692 16156 21308 16212
rect 21364 16156 21374 16212
rect 16706 16044 16716 16100
rect 16772 16044 17612 16100
rect 17668 16044 18172 16100
rect 18228 16044 18508 16100
rect 18564 16044 18574 16100
rect 14354 15820 14364 15876
rect 14420 15820 15484 15876
rect 15540 15820 15550 15876
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 16482 15484 16492 15540
rect 16548 15484 17388 15540
rect 17444 15484 17454 15540
rect 20626 15484 20636 15540
rect 20692 15484 22876 15540
rect 22932 15484 22942 15540
rect 25330 15372 25340 15428
rect 25396 15372 26012 15428
rect 26068 15372 26078 15428
rect 17938 15260 17948 15316
rect 18004 15260 18396 15316
rect 18452 15260 20188 15316
rect 20244 15260 20254 15316
rect 20738 15260 20748 15316
rect 20804 15260 22092 15316
rect 22148 15260 22158 15316
rect 22754 15260 22764 15316
rect 22820 15260 25228 15316
rect 25284 15260 25294 15316
rect 20402 15036 20412 15092
rect 20468 15036 21084 15092
rect 21140 15036 25564 15092
rect 25620 15036 27132 15092
rect 27188 15036 27198 15092
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 13682 14588 13692 14644
rect 13748 14588 15372 14644
rect 15428 14588 16716 14644
rect 16772 14588 18732 14644
rect 18788 14588 21868 14644
rect 21924 14588 22988 14644
rect 23044 14588 24780 14644
rect 24836 14588 24846 14644
rect 16034 14252 16044 14308
rect 16100 14252 17164 14308
rect 17220 14252 17612 14308
rect 17668 14252 17678 14308
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 26450 13580 26460 13636
rect 26516 13580 27132 13636
rect 27188 13580 27916 13636
rect 27972 13580 27982 13636
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 26898 4060 26908 4116
rect 26964 4060 28140 4116
rect 28196 4060 28206 4116
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 24210 3612 24220 3668
rect 24276 3612 25564 3668
rect 25620 3612 25630 3668
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
<< via3 >>
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 19516 20076 19572 20132
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 19516 17052 19572 17108
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
<< metal4 >>
rect 4448 38444 4768 38476
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 19808 37660 20128 38476
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19808 34524 20128 36036
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 19808 23548 20128 25060
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 19808 21980 20128 23492
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 19516 20132 19572 20142
rect 19516 17108 19572 20076
rect 19516 17042 19572 17052
rect 19808 18844 20128 20356
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 38444 35488 38476
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _106_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 19936 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _107_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18928 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _108_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 22960 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _109_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 18144 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _110_
timestamp 1698175906
transform 1 0 16016 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _111_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 16912 0 1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _112_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 28000 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _113_
timestamp 1698175906
transform 1 0 21392 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _114_
timestamp 1698175906
transform -1 0 22064 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _115_
timestamp 1698175906
transform 1 0 23408 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _116_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 25648 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _117_
timestamp 1698175906
transform 1 0 18144 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _118_
timestamp 1698175906
transform -1 0 19712 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _119_
timestamp 1698175906
transform -1 0 17024 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _120_
timestamp 1698175906
transform 1 0 20272 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _121_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17248 0 -1 21952
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _122_
timestamp 1698175906
transform 1 0 22736 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _123_
timestamp 1698175906
transform -1 0 23632 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _124_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 18032 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _125_
timestamp 1698175906
transform -1 0 16912 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _126_
timestamp 1698175906
transform -1 0 20720 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _127_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 19376 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _128_
timestamp 1698175906
transform 1 0 21616 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _129_
timestamp 1698175906
transform 1 0 22624 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _130_
timestamp 1698175906
transform 1 0 23296 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _131_
timestamp 1698175906
transform -1 0 23296 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _132_
timestamp 1698175906
transform 1 0 17248 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _133_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 19040 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _134_
timestamp 1698175906
transform -1 0 17808 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _135_
timestamp 1698175906
transform -1 0 16016 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _136_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18256 0 1 15680
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _137_
timestamp 1698175906
transform -1 0 18592 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _138_
timestamp 1698175906
transform 1 0 17472 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _139_
timestamp 1698175906
transform 1 0 21504 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _140_
timestamp 1698175906
transform -1 0 22848 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _141_
timestamp 1698175906
transform -1 0 20720 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _142_
timestamp 1698175906
transform 1 0 18032 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _143_
timestamp 1698175906
transform 1 0 19712 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _144_
timestamp 1698175906
transform -1 0 20048 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _145_
timestamp 1698175906
transform 1 0 18928 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _146_
timestamp 1698175906
transform -1 0 18592 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _147_
timestamp 1698175906
transform -1 0 26656 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _148_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 21728 0 -1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _149_
timestamp 1698175906
transform 1 0 21840 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _150_
timestamp 1698175906
transform -1 0 26208 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _151_
timestamp 1698175906
transform -1 0 22064 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _152_
timestamp 1698175906
transform -1 0 18928 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _153_
timestamp 1698175906
transform -1 0 16352 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _154_
timestamp 1698175906
transform -1 0 15792 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _155_
timestamp 1698175906
transform -1 0 16240 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _156_
timestamp 1698175906
transform -1 0 15456 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _157_
timestamp 1698175906
transform 1 0 24192 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _158_
timestamp 1698175906
transform 1 0 26320 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _159_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 26432 0 -1 20384
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _160_
timestamp 1698175906
transform -1 0 17024 0 -1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _161_
timestamp 1698175906
transform 1 0 16352 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _162_
timestamp 1698175906
transform 1 0 18032 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _163_
timestamp 1698175906
transform -1 0 19264 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _164_
timestamp 1698175906
transform -1 0 18704 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _165_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19600 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _166_
timestamp 1698175906
transform -1 0 23968 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _167_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 23408 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _168_
timestamp 1698175906
transform -1 0 16240 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _169_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18032 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _170_
timestamp 1698175906
transform -1 0 14672 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _171_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 15904 0 -1 18816
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _172_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 15344 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _173_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 14000 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _174_
timestamp 1698175906
transform -1 0 17024 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _175_
timestamp 1698175906
transform -1 0 20944 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _176_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 14112 0 -1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _177_
timestamp 1698175906
transform -1 0 15680 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _178_
timestamp 1698175906
transform -1 0 15008 0 1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _179_
timestamp 1698175906
transform -1 0 25984 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _180_
timestamp 1698175906
transform -1 0 19600 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _181_
timestamp 1698175906
transform 1 0 23296 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _182_
timestamp 1698175906
transform 1 0 23632 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _183_
timestamp 1698175906
transform 1 0 24080 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _184_
timestamp 1698175906
transform -1 0 26208 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _185_
timestamp 1698175906
transform -1 0 25648 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _186_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17920 0 -1 17248
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _187_
timestamp 1698175906
transform -1 0 21504 0 -1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _188_
timestamp 1698175906
transform 1 0 15120 0 -1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _189_
timestamp 1698175906
transform -1 0 15120 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _190_
timestamp 1698175906
transform -1 0 29456 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _191_
timestamp 1698175906
transform -1 0 28000 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _192_
timestamp 1698175906
transform -1 0 20160 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _193_
timestamp 1698175906
transform 1 0 19600 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _194_
timestamp 1698175906
transform -1 0 19600 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _195_
timestamp 1698175906
transform 1 0 20944 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _196_
timestamp 1698175906
transform -1 0 28000 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _197_
timestamp 1698175906
transform 1 0 25088 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _198_
timestamp 1698175906
transform 1 0 25536 0 1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _199_
timestamp 1698175906
transform -1 0 16352 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _200_
timestamp 1698175906
transform 1 0 15120 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _201_
timestamp 1698175906
transform 1 0 16128 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _202_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 15904 0 1 21952
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _203_
timestamp 1698175906
transform 1 0 13440 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _204_
timestamp 1698175906
transform -1 0 23184 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _205_
timestamp 1698175906
transform -1 0 22736 0 1 23520
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _206_
timestamp 1698175906
transform -1 0 27440 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  _207_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 24864 0 1 23520
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _208_
timestamp 1698175906
transform -1 0 24528 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _209_
timestamp 1698175906
transform -1 0 24528 0 -1 21952
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _210_
timestamp 1698175906
transform 1 0 15120 0 -1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _211_
timestamp 1698175906
transform 1 0 13216 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _212_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 26096 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _213_
timestamp 1698175906
transform 1 0 14224 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _214_
timestamp 1698175906
transform 1 0 21280 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _215_
timestamp 1698175906
transform 1 0 15120 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _216_
timestamp 1698175906
transform 1 0 13440 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _217_
timestamp 1698175906
transform 1 0 18592 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _218_
timestamp 1698175906
transform 1 0 17136 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _219_
timestamp 1698175906
transform 1 0 24864 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _220_
timestamp 1698175906
transform 1 0 13104 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _221_
timestamp 1698175906
transform 1 0 26432 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _222_
timestamp 1698175906
transform 1 0 17248 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _223_
timestamp 1698175906
transform 1 0 21616 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _224_
timestamp 1698175906
transform -1 0 14560 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _225_
timestamp 1698175906
transform -1 0 13104 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _226_
timestamp 1698175906
transform 1 0 22848 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _227_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 24416 0 1 26656
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _228_
timestamp 1698175906
transform -1 0 14448 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _229_
timestamp 1698175906
transform 1 0 26768 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _230_
timestamp 1698175906
transform 1 0 17696 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _231_
timestamp 1698175906
transform 1 0 25872 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _232_
timestamp 1698175906
transform -1 0 15120 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _233_
timestamp 1698175906
transform 1 0 20608 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _234_
timestamp 1698175906
transform 1 0 25424 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _235_
timestamp 1698175906
transform 1 0 22288 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _236_
timestamp 1698175906
transform -1 0 13104 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _238_
timestamp 1698175906
transform 1 0 27888 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _239_
timestamp 1698175906
transform 1 0 20048 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _240_
timestamp 1698175906
transform 1 0 29680 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _241_
timestamp 1698175906
transform 1 0 26656 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__212__CLK dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 26320 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__213__CLK
timestamp 1698175906
transform 1 0 17472 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__214__CLK
timestamp 1698175906
transform -1 0 21280 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__215__CLK
timestamp 1698175906
transform -1 0 18816 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__216__CLK
timestamp 1698175906
transform 1 0 16688 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__217__CLK
timestamp 1698175906
transform 1 0 22064 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__218__CLK
timestamp 1698175906
transform 1 0 20608 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__219__CLK
timestamp 1698175906
transform 1 0 24640 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__220__CLK
timestamp 1698175906
transform 1 0 16352 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__221__CLK
timestamp 1698175906
transform 1 0 26992 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__222__CLK
timestamp 1698175906
transform 1 0 20496 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__223__CLK
timestamp 1698175906
transform 1 0 25312 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__224__CLK
timestamp 1698175906
transform 1 0 14784 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__225__CLK
timestamp 1698175906
transform -1 0 13776 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__226__CLK
timestamp 1698175906
transform 1 0 26768 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__227__CLK
timestamp 1698175906
transform 1 0 24192 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__228__CLK
timestamp 1698175906
transform 1 0 14672 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__229__CLK
timestamp 1698175906
transform 1 0 25424 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__230__CLK
timestamp 1698175906
transform 1 0 21392 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__231__CLK
timestamp 1698175906
transform 1 0 25648 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__232__CLK
timestamp 1698175906
transform 1 0 15792 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__233__CLK
timestamp 1698175906
transform 1 0 23856 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__234__CLK
timestamp 1698175906
transform 1 0 25200 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__235__CLK
timestamp 1698175906
transform 1 0 21392 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__236__CLK
timestamp 1698175906
transform 1 0 13552 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1698175906
transform -1 0 20272 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21168 0 1 20384
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1698175906
transform -1 0 26768 0 1 17248
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1698175906
transform -1 0 24864 0 -1 23520
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1568 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698175906
transform 1 0 5376 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_70 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9184 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_86 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10976 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_94 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 11872 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_96 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 12096 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_101
timestamp 1698175906
transform 1 0 12656 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698175906
transform 1 0 12992 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_138
timestamp 1698175906
transform 1 0 16800 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_172
timestamp 1698175906
transform 1 0 20608 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_232 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 27328 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_236
timestamp 1698175906
transform 1 0 27776 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_240
timestamp 1698175906
transform 1 0 28224 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_274
timestamp 1698175906
transform 1 0 32032 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_308
timestamp 1698175906
transform 1 0 35840 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_342
timestamp 1698175906
transform 1 0 39648 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_346
timestamp 1698175906
transform 1 0 40096 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_348
timestamp 1698175906
transform 1 0 40320 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1568 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698175906
transform 1 0 8736 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698175906
transform 1 0 9408 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698175906
transform 1 0 16576 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_142
timestamp 1698175906
transform 1 0 17248 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_206
timestamp 1698175906
transform 1 0 24416 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_212
timestamp 1698175906
transform 1 0 25088 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_228
timestamp 1698175906
transform 1 0 26880 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_255
timestamp 1698175906
transform 1 0 29904 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_271
timestamp 1698175906
transform 1 0 31696 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_279
timestamp 1698175906
transform 1 0 32592 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_282
timestamp 1698175906
transform 1 0 32928 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_346
timestamp 1698175906
transform 1 0 40096 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_348
timestamp 1698175906
transform 1 0 40320 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698175906
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698175906
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698175906
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698175906
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_107
timestamp 1698175906
transform 1 0 13328 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_171
timestamp 1698175906
transform 1 0 20496 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_177
timestamp 1698175906
transform 1 0 21168 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_241
timestamp 1698175906
transform 1 0 28336 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698175906
transform 1 0 29008 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698175906
transform 1 0 36176 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_317
timestamp 1698175906
transform 1 0 36848 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698175906
transform 1 0 1568 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698175906
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698175906
transform 1 0 9408 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698175906
transform 1 0 16576 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_142
timestamp 1698175906
transform 1 0 17248 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_206
timestamp 1698175906
transform 1 0 24416 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_212
timestamp 1698175906
transform 1 0 25088 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_276
timestamp 1698175906
transform 1 0 32256 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_282
timestamp 1698175906
transform 1 0 32928 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_346
timestamp 1698175906
transform 1 0 40096 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_348
timestamp 1698175906
transform 1 0 40320 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698175906
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698175906
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698175906
transform 1 0 5488 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698175906
transform 1 0 12656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_107
timestamp 1698175906
transform 1 0 13328 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698175906
transform 1 0 20496 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_177
timestamp 1698175906
transform 1 0 21168 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_241
timestamp 1698175906
transform 1 0 28336 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698175906
transform 1 0 29008 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698175906
transform 1 0 36176 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_317
timestamp 1698175906
transform 1 0 36848 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698175906
transform 1 0 1568 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698175906
transform 1 0 8736 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698175906
transform 1 0 9408 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698175906
transform 1 0 16576 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_142
timestamp 1698175906
transform 1 0 17248 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_206
timestamp 1698175906
transform 1 0 24416 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_212
timestamp 1698175906
transform 1 0 25088 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698175906
transform 1 0 32256 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_282
timestamp 1698175906
transform 1 0 32928 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_346
timestamp 1698175906
transform 1 0 40096 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_348
timestamp 1698175906
transform 1 0 40320 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698175906
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698175906
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698175906
transform 1 0 5488 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698175906
transform 1 0 12656 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_107
timestamp 1698175906
transform 1 0 13328 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_171
timestamp 1698175906
transform 1 0 20496 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_177
timestamp 1698175906
transform 1 0 21168 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_241
timestamp 1698175906
transform 1 0 28336 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_247
timestamp 1698175906
transform 1 0 29008 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_311
timestamp 1698175906
transform 1 0 36176 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_317
timestamp 1698175906
transform 1 0 36848 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698175906
transform 1 0 1568 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698175906
transform 1 0 8736 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_72
timestamp 1698175906
transform 1 0 9408 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698175906
transform 1 0 16576 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_142
timestamp 1698175906
transform 1 0 17248 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_206
timestamp 1698175906
transform 1 0 24416 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_212
timestamp 1698175906
transform 1 0 25088 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_276
timestamp 1698175906
transform 1 0 32256 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_282
timestamp 1698175906
transform 1 0 32928 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_346
timestamp 1698175906
transform 1 0 40096 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_348
timestamp 1698175906
transform 1 0 40320 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698175906
transform 1 0 1568 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698175906
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_37
timestamp 1698175906
transform 1 0 5488 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_101
timestamp 1698175906
transform 1 0 12656 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_107
timestamp 1698175906
transform 1 0 13328 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_171
timestamp 1698175906
transform 1 0 20496 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_177
timestamp 1698175906
transform 1 0 21168 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_241
timestamp 1698175906
transform 1 0 28336 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_247
timestamp 1698175906
transform 1 0 29008 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_311
timestamp 1698175906
transform 1 0 36176 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_317
timestamp 1698175906
transform 1 0 36848 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698175906
transform 1 0 1568 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698175906
transform 1 0 8736 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_72
timestamp 1698175906
transform 1 0 9408 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_136
timestamp 1698175906
transform 1 0 16576 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_142
timestamp 1698175906
transform 1 0 17248 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_206
timestamp 1698175906
transform 1 0 24416 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_212
timestamp 1698175906
transform 1 0 25088 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_276
timestamp 1698175906
transform 1 0 32256 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_282
timestamp 1698175906
transform 1 0 32928 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_346
timestamp 1698175906
transform 1 0 40096 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_348
timestamp 1698175906
transform 1 0 40320 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698175906
transform 1 0 1568 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698175906
transform 1 0 5152 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_37
timestamp 1698175906
transform 1 0 5488 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698175906
transform 1 0 12656 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_107
timestamp 1698175906
transform 1 0 13328 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_171
timestamp 1698175906
transform 1 0 20496 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_177
timestamp 1698175906
transform 1 0 21168 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_241
timestamp 1698175906
transform 1 0 28336 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_247
timestamp 1698175906
transform 1 0 29008 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_311
timestamp 1698175906
transform 1 0 36176 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_317
timestamp 1698175906
transform 1 0 36848 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2
timestamp 1698175906
transform 1 0 1568 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698175906
transform 1 0 8736 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_72
timestamp 1698175906
transform 1 0 9408 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698175906
transform 1 0 16576 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_142
timestamp 1698175906
transform 1 0 17248 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_206
timestamp 1698175906
transform 1 0 24416 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_212
timestamp 1698175906
transform 1 0 25088 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_276
timestamp 1698175906
transform 1 0 32256 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_282
timestamp 1698175906
transform 1 0 32928 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_346
timestamp 1698175906
transform 1 0 40096 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_348
timestamp 1698175906
transform 1 0 40320 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698175906
transform 1 0 1568 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698175906
transform 1 0 5152 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_37
timestamp 1698175906
transform 1 0 5488 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698175906
transform 1 0 12656 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_107
timestamp 1698175906
transform 1 0 13328 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_152
timestamp 1698175906
transform 1 0 18368 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_156
timestamp 1698175906
transform 1 0 18816 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_172
timestamp 1698175906
transform 1 0 20608 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_174
timestamp 1698175906
transform 1 0 20832 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_177
timestamp 1698175906
transform 1 0 21168 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_241
timestamp 1698175906
transform 1 0 28336 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_247
timestamp 1698175906
transform 1 0 29008 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_311
timestamp 1698175906
transform 1 0 36176 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_317
timestamp 1698175906
transform 1 0 36848 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_2
timestamp 1698175906
transform 1 0 1568 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_66
timestamp 1698175906
transform 1 0 8736 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_72
timestamp 1698175906
transform 1 0 9408 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_136
timestamp 1698175906
transform 1 0 16576 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_142
timestamp 1698175906
transform 1 0 17248 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_150
timestamp 1698175906
transform 1 0 18144 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_183
timestamp 1698175906
transform 1 0 21840 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_187
timestamp 1698175906
transform 1 0 22288 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_195
timestamp 1698175906
transform 1 0 23184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_202
timestamp 1698175906
transform 1 0 23968 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_206
timestamp 1698175906
transform 1 0 24416 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_212
timestamp 1698175906
transform 1 0 25088 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_216
timestamp 1698175906
transform 1 0 25536 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_220
timestamp 1698175906
transform 1 0 25984 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_226
timestamp 1698175906
transform 1 0 26656 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_258
timestamp 1698175906
transform 1 0 30240 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_274
timestamp 1698175906
transform 1 0 32032 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_278
timestamp 1698175906
transform 1 0 32480 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_282
timestamp 1698175906
transform 1 0 32928 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_346
timestamp 1698175906
transform 1 0 40096 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_348
timestamp 1698175906
transform 1 0 40320 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698175906
transform 1 0 1568 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698175906
transform 1 0 5152 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_37
timestamp 1698175906
transform 1 0 5488 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_101
timestamp 1698175906
transform 1 0 12656 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_107
timestamp 1698175906
transform 1 0 13328 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_123
timestamp 1698175906
transform 1 0 15120 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_131
timestamp 1698175906
transform 1 0 16016 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_135
timestamp 1698175906
transform 1 0 16464 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_139
timestamp 1698175906
transform 1 0 16912 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_143
timestamp 1698175906
transform 1 0 17360 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_170
timestamp 1698175906
transform 1 0 20384 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_174
timestamp 1698175906
transform 1 0 20832 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_177
timestamp 1698175906
transform 1 0 21168 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_239
timestamp 1698175906
transform 1 0 28112 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_243
timestamp 1698175906
transform 1 0 28560 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_247
timestamp 1698175906
transform 1 0 29008 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_311
timestamp 1698175906
transform 1 0 36176 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_317
timestamp 1698175906
transform 1 0 36848 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_2
timestamp 1698175906
transform 1 0 1568 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_66
timestamp 1698175906
transform 1 0 8736 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_72
timestamp 1698175906
transform 1 0 9408 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_104
timestamp 1698175906
transform 1 0 12992 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_137
timestamp 1698175906
transform 1 0 16688 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_139
timestamp 1698175906
transform 1 0 16912 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_150
timestamp 1698175906
transform 1 0 18144 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_161
timestamp 1698175906
transform 1 0 19376 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_173
timestamp 1698175906
transform 1 0 20720 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_177
timestamp 1698175906
transform 1 0 21168 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_187
timestamp 1698175906
transform 1 0 22288 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_197
timestamp 1698175906
transform 1 0 23408 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_205
timestamp 1698175906
transform 1 0 24304 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_209
timestamp 1698175906
transform 1 0 24752 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_222
timestamp 1698175906
transform 1 0 26208 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_254
timestamp 1698175906
transform 1 0 29792 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_270
timestamp 1698175906
transform 1 0 31584 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_278
timestamp 1698175906
transform 1 0 32480 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_282
timestamp 1698175906
transform 1 0 32928 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_346
timestamp 1698175906
transform 1 0 40096 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_348
timestamp 1698175906
transform 1 0 40320 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_2
timestamp 1698175906
transform 1 0 1568 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698175906
transform 1 0 5152 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_37
timestamp 1698175906
transform 1 0 5488 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_101
timestamp 1698175906
transform 1 0 12656 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_113
timestamp 1698175906
transform 1 0 14000 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_121
timestamp 1698175906
transform 1 0 14896 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_125
timestamp 1698175906
transform 1 0 15344 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_148
timestamp 1698175906
transform 1 0 17920 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_150
timestamp 1698175906
transform 1 0 18144 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_185
timestamp 1698175906
transform 1 0 22064 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_189
timestamp 1698175906
transform 1 0 22512 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_191
timestamp 1698175906
transform 1 0 22736 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_221
timestamp 1698175906
transform 1 0 26096 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_225
timestamp 1698175906
transform 1 0 26544 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_229
timestamp 1698175906
transform 1 0 26992 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_247
timestamp 1698175906
transform 1 0 29008 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_311
timestamp 1698175906
transform 1 0 36176 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_317
timestamp 1698175906
transform 1 0 36848 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_2
timestamp 1698175906
transform 1 0 1568 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_66
timestamp 1698175906
transform 1 0 8736 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_72
timestamp 1698175906
transform 1 0 9408 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_88
timestamp 1698175906
transform 1 0 11200 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_118
timestamp 1698175906
transform 1 0 14560 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_122
timestamp 1698175906
transform 1 0 15008 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_147
timestamp 1698175906
transform 1 0 17808 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_185
timestamp 1698175906
transform 1 0 22064 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_193
timestamp 1698175906
transform 1 0 22960 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_195
timestamp 1698175906
transform 1 0 23184 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_201
timestamp 1698175906
transform 1 0 23856 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_209
timestamp 1698175906
transform 1 0 24752 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_220
timestamp 1698175906
transform 1 0 25984 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_250
timestamp 1698175906
transform 1 0 29344 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_266
timestamp 1698175906
transform 1 0 31136 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_274
timestamp 1698175906
transform 1 0 32032 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_278
timestamp 1698175906
transform 1 0 32480 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_282
timestamp 1698175906
transform 1 0 32928 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_314
timestamp 1698175906
transform 1 0 36512 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_322
timestamp 1698175906
transform 1 0 37408 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_28
timestamp 1698175906
transform 1 0 4480 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_32
timestamp 1698175906
transform 1 0 4928 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698175906
transform 1 0 5152 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_37
timestamp 1698175906
transform 1 0 5488 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_101
timestamp 1698175906
transform 1 0 12656 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_107
timestamp 1698175906
transform 1 0 13328 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_115
timestamp 1698175906
transform 1 0 14224 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_125
timestamp 1698175906
transform 1 0 15344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_127
timestamp 1698175906
transform 1 0 15568 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_133
timestamp 1698175906
transform 1 0 16240 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_141
timestamp 1698175906
transform 1 0 17136 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_145
timestamp 1698175906
transform 1 0 17584 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_147
timestamp 1698175906
transform 1 0 17808 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_158
timestamp 1698175906
transform 1 0 19040 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_160
timestamp 1698175906
transform 1 0 19264 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_227
timestamp 1698175906
transform 1 0 26768 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_244
timestamp 1698175906
transform 1 0 28672 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_251
timestamp 1698175906
transform 1 0 29456 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_317
timestamp 1698175906
transform 1 0 36848 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_321
timestamp 1698175906
transform 1 0 37296 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_2
timestamp 1698175906
transform 1 0 1568 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_66
timestamp 1698175906
transform 1 0 8736 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_72
timestamp 1698175906
transform 1 0 9408 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_104
timestamp 1698175906
transform 1 0 12992 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_112
timestamp 1698175906
transform 1 0 13888 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_130
timestamp 1698175906
transform 1 0 15904 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_138
timestamp 1698175906
transform 1 0 16800 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_142
timestamp 1698175906
transform 1 0 17248 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_146
timestamp 1698175906
transform 1 0 17696 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_148
timestamp 1698175906
transform 1 0 17920 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_165
timestamp 1698175906
transform 1 0 19824 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_169
timestamp 1698175906
transform 1 0 20272 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_182
timestamp 1698175906
transform 1 0 21728 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_189
timestamp 1698175906
transform 1 0 22512 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_204
timestamp 1698175906
transform 1 0 24192 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_208
timestamp 1698175906
transform 1 0 24640 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_212
timestamp 1698175906
transform 1 0 25088 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_214
timestamp 1698175906
transform 1 0 25312 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_256
timestamp 1698175906
transform 1 0 30016 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_272
timestamp 1698175906
transform 1 0 31808 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_282
timestamp 1698175906
transform 1 0 32928 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_314
timestamp 1698175906
transform 1 0 36512 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_322
timestamp 1698175906
transform 1 0 37408 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_2
timestamp 1698175906
transform 1 0 1568 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698175906
transform 1 0 5152 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_37
timestamp 1698175906
transform 1 0 5488 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_69
timestamp 1698175906
transform 1 0 9072 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_73
timestamp 1698175906
transform 1 0 9520 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_75
timestamp 1698175906
transform 1 0 9744 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_107
timestamp 1698175906
transform 1 0 13328 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_111
timestamp 1698175906
transform 1 0 13776 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_119
timestamp 1698175906
transform 1 0 14672 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_140
timestamp 1698175906
transform 1 0 17024 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_173
timestamp 1698175906
transform 1 0 20720 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_177
timestamp 1698175906
transform 1 0 21168 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_179
timestamp 1698175906
transform 1 0 21392 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_192
timestamp 1698175906
transform 1 0 22848 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_200
timestamp 1698175906
transform 1 0 23744 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_207
timestamp 1698175906
transform 1 0 24528 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_228
timestamp 1698175906
transform 1 0 26880 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_244
timestamp 1698175906
transform 1 0 28672 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_247
timestamp 1698175906
transform 1 0 29008 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_311
timestamp 1698175906
transform 1 0 36176 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_317
timestamp 1698175906
transform 1 0 36848 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_28
timestamp 1698175906
transform 1 0 4480 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_60
timestamp 1698175906
transform 1 0 8064 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_68
timestamp 1698175906
transform 1 0 8960 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_72
timestamp 1698175906
transform 1 0 9408 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_104
timestamp 1698175906
transform 1 0 12992 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_132
timestamp 1698175906
transform 1 0 16128 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_142
timestamp 1698175906
transform 1 0 17248 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_150
timestamp 1698175906
transform 1 0 18144 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_166
timestamp 1698175906
transform 1 0 19936 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_180
timestamp 1698175906
transform 1 0 21504 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_185
timestamp 1698175906
transform 1 0 22064 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_189
timestamp 1698175906
transform 1 0 22512 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_203
timestamp 1698175906
transform 1 0 24080 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_212
timestamp 1698175906
transform 1 0 25088 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_259
timestamp 1698175906
transform 1 0 30352 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_275
timestamp 1698175906
transform 1 0 32144 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_279
timestamp 1698175906
transform 1 0 32592 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_282
timestamp 1698175906
transform 1 0 32928 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_346
timestamp 1698175906
transform 1 0 40096 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_348
timestamp 1698175906
transform 1 0 40320 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_28
timestamp 1698175906
transform 1 0 4480 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_32
timestamp 1698175906
transform 1 0 4928 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698175906
transform 1 0 5152 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_37
timestamp 1698175906
transform 1 0 5488 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_69
timestamp 1698175906
transform 1 0 9072 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_73
timestamp 1698175906
transform 1 0 9520 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_75
timestamp 1698175906
transform 1 0 9744 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_107
timestamp 1698175906
transform 1 0 13328 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_111
timestamp 1698175906
transform 1 0 13776 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_122
timestamp 1698175906
transform 1 0 15008 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_154
timestamp 1698175906
transform 1 0 18592 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_162
timestamp 1698175906
transform 1 0 19488 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_166
timestamp 1698175906
transform 1 0 19936 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_227
timestamp 1698175906
transform 1 0 26768 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_231
timestamp 1698175906
transform 1 0 27216 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_239
timestamp 1698175906
transform 1 0 28112 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_243
timestamp 1698175906
transform 1 0 28560 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_247
timestamp 1698175906
transform 1 0 29008 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_311
timestamp 1698175906
transform 1 0 36176 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_317
timestamp 1698175906
transform 1 0 36848 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_321
timestamp 1698175906
transform 1 0 37296 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_2
timestamp 1698175906
transform 1 0 1568 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_66
timestamp 1698175906
transform 1 0 8736 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_72
timestamp 1698175906
transform 1 0 9408 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_117
timestamp 1698175906
transform 1 0 14448 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_121
timestamp 1698175906
transform 1 0 14896 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_123
timestamp 1698175906
transform 1 0 15120 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_154
timestamp 1698175906
transform 1 0 18592 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_162
timestamp 1698175906
transform 1 0 19488 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_166
timestamp 1698175906
transform 1 0 19936 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_173
timestamp 1698175906
transform 1 0 20720 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_181
timestamp 1698175906
transform 1 0 21616 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_189
timestamp 1698175906
transform 1 0 22512 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_193
timestamp 1698175906
transform 1 0 22960 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_195
timestamp 1698175906
transform 1 0 23184 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_207
timestamp 1698175906
transform 1 0 24528 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_209
timestamp 1698175906
transform 1 0 24752 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_217
timestamp 1698175906
transform 1 0 25648 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_249
timestamp 1698175906
transform 1 0 29232 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_265
timestamp 1698175906
transform 1 0 31024 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_273
timestamp 1698175906
transform 1 0 31920 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_277
timestamp 1698175906
transform 1 0 32368 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_279
timestamp 1698175906
transform 1 0 32592 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_282
timestamp 1698175906
transform 1 0 32928 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_314
timestamp 1698175906
transform 1 0 36512 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_322
timestamp 1698175906
transform 1 0 37408 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_2
timestamp 1698175906
transform 1 0 1568 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698175906
transform 1 0 5152 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_37
timestamp 1698175906
transform 1 0 5488 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_101
timestamp 1698175906
transform 1 0 12656 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_107
timestamp 1698175906
transform 1 0 13328 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_114
timestamp 1698175906
transform 1 0 14112 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_118
timestamp 1698175906
transform 1 0 14560 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_130
timestamp 1698175906
transform 1 0 15904 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_138
timestamp 1698175906
transform 1 0 16800 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_140
timestamp 1698175906
transform 1 0 17024 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_170
timestamp 1698175906
transform 1 0 20384 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_174
timestamp 1698175906
transform 1 0 20832 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_177
timestamp 1698175906
transform 1 0 21168 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_225
timestamp 1698175906
transform 1 0 26544 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_227
timestamp 1698175906
transform 1 0 26768 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_238
timestamp 1698175906
transform 1 0 28000 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_242
timestamp 1698175906
transform 1 0 28448 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_244
timestamp 1698175906
transform 1 0 28672 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_247
timestamp 1698175906
transform 1 0 29008 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_311
timestamp 1698175906
transform 1 0 36176 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_317
timestamp 1698175906
transform 1 0 36848 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_321
timestamp 1698175906
transform 1 0 37296 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_28
timestamp 1698175906
transform 1 0 4480 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_60
timestamp 1698175906
transform 1 0 8064 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_68
timestamp 1698175906
transform 1 0 8960 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_72
timestamp 1698175906
transform 1 0 9408 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_88
timestamp 1698175906
transform 1 0 11200 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_92
timestamp 1698175906
transform 1 0 11648 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_142
timestamp 1698175906
transform 1 0 17248 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_158
timestamp 1698175906
transform 1 0 19040 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_212
timestamp 1698175906
transform 1 0 25088 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_216
timestamp 1698175906
transform 1 0 25536 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_248
timestamp 1698175906
transform 1 0 29120 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_282
timestamp 1698175906
transform 1 0 32928 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_314
timestamp 1698175906
transform 1 0 36512 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_322
timestamp 1698175906
transform 1 0 37408 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_28
timestamp 1698175906
transform 1 0 4480 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_32
timestamp 1698175906
transform 1 0 4928 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698175906
transform 1 0 5152 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_37
timestamp 1698175906
transform 1 0 5488 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_101
timestamp 1698175906
transform 1 0 12656 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_107
timestamp 1698175906
transform 1 0 13328 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_115
timestamp 1698175906
transform 1 0 14224 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_127
timestamp 1698175906
transform 1 0 15568 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_131
timestamp 1698175906
transform 1 0 16016 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_147
timestamp 1698175906
transform 1 0 17808 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_154
timestamp 1698175906
transform 1 0 18592 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_162
timestamp 1698175906
transform 1 0 19488 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_171
timestamp 1698175906
transform 1 0 20496 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_177
timestamp 1698175906
transform 1 0 21168 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_179
timestamp 1698175906
transform 1 0 21392 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_195
timestamp 1698175906
transform 1 0 23184 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_210
timestamp 1698175906
transform 1 0 24864 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_212
timestamp 1698175906
transform 1 0 25088 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_244
timestamp 1698175906
transform 1 0 28672 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_247
timestamp 1698175906
transform 1 0 29008 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_311
timestamp 1698175906
transform 1 0 36176 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_317
timestamp 1698175906
transform 1 0 36848 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_321
timestamp 1698175906
transform 1 0 37296 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_2
timestamp 1698175906
transform 1 0 1568 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_66
timestamp 1698175906
transform 1 0 8736 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_72
timestamp 1698175906
transform 1 0 9408 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_136
timestamp 1698175906
transform 1 0 16576 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_142
timestamp 1698175906
transform 1 0 17248 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_168
timestamp 1698175906
transform 1 0 20160 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_201
timestamp 1698175906
transform 1 0 23856 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_208
timestamp 1698175906
transform 1 0 24640 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_212
timestamp 1698175906
transform 1 0 25088 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_276
timestamp 1698175906
transform 1 0 32256 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_282
timestamp 1698175906
transform 1 0 32928 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_346
timestamp 1698175906
transform 1 0 40096 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_348
timestamp 1698175906
transform 1 0 40320 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_2
timestamp 1698175906
transform 1 0 1568 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698175906
transform 1 0 5152 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_37
timestamp 1698175906
transform 1 0 5488 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_101
timestamp 1698175906
transform 1 0 12656 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_107
timestamp 1698175906
transform 1 0 13328 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_115
timestamp 1698175906
transform 1 0 14224 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_119
timestamp 1698175906
transform 1 0 14672 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_126
timestamp 1698175906
transform 1 0 15456 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_136
timestamp 1698175906
transform 1 0 16576 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_144
timestamp 1698175906
transform 1 0 17472 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_177
timestamp 1698175906
transform 1 0 21168 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_181
timestamp 1698175906
transform 1 0 21616 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_189
timestamp 1698175906
transform 1 0 22512 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_195
timestamp 1698175906
transform 1 0 23184 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_199
timestamp 1698175906
transform 1 0 23632 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_203
timestamp 1698175906
transform 1 0 24080 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_235
timestamp 1698175906
transform 1 0 27664 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_243
timestamp 1698175906
transform 1 0 28560 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_247
timestamp 1698175906
transform 1 0 29008 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_311
timestamp 1698175906
transform 1 0 36176 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_317
timestamp 1698175906
transform 1 0 36848 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_2
timestamp 1698175906
transform 1 0 1568 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_66
timestamp 1698175906
transform 1 0 8736 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_72
timestamp 1698175906
transform 1 0 9408 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_104
timestamp 1698175906
transform 1 0 12992 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_139
timestamp 1698175906
transform 1 0 16912 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_142
timestamp 1698175906
transform 1 0 17248 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_146
timestamp 1698175906
transform 1 0 17696 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_162
timestamp 1698175906
transform 1 0 19488 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_166
timestamp 1698175906
transform 1 0 19936 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_173
timestamp 1698175906
transform 1 0 20720 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_189
timestamp 1698175906
transform 1 0 22512 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_199
timestamp 1698175906
transform 1 0 23632 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_207
timestamp 1698175906
transform 1 0 24528 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_209
timestamp 1698175906
transform 1 0 24752 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_222
timestamp 1698175906
transform 1 0 26208 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_232
timestamp 1698175906
transform 1 0 27328 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_264
timestamp 1698175906
transform 1 0 30912 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_282
timestamp 1698175906
transform 1 0 32928 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_314
timestamp 1698175906
transform 1 0 36512 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_322
timestamp 1698175906
transform 1 0 37408 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_2
timestamp 1698175906
transform 1 0 1568 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698175906
transform 1 0 5152 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_37
timestamp 1698175906
transform 1 0 5488 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_101
timestamp 1698175906
transform 1 0 12656 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_107
timestamp 1698175906
transform 1 0 13328 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_149
timestamp 1698175906
transform 1 0 18032 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_160
timestamp 1698175906
transform 1 0 19264 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_168
timestamp 1698175906
transform 1 0 20160 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_170
timestamp 1698175906
transform 1 0 20384 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_173
timestamp 1698175906
transform 1 0 20720 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_177
timestamp 1698175906
transform 1 0 21168 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_185
timestamp 1698175906
transform 1 0 22064 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_189
timestamp 1698175906
transform 1 0 22512 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_201
timestamp 1698175906
transform 1 0 23856 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_203
timestamp 1698175906
transform 1 0 24080 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_243
timestamp 1698175906
transform 1 0 28560 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_247
timestamp 1698175906
transform 1 0 29008 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_311
timestamp 1698175906
transform 1 0 36176 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_317
timestamp 1698175906
transform 1 0 36848 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_321
timestamp 1698175906
transform 1 0 37296 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_2
timestamp 1698175906
transform 1 0 1568 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_66
timestamp 1698175906
transform 1 0 8736 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_72
timestamp 1698175906
transform 1 0 9408 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_104
timestamp 1698175906
transform 1 0 12992 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_120
timestamp 1698175906
transform 1 0 14784 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_133
timestamp 1698175906
transform 1 0 16240 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_137
timestamp 1698175906
transform 1 0 16688 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_139
timestamp 1698175906
transform 1 0 16912 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_171
timestamp 1698175906
transform 1 0 20496 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_175
timestamp 1698175906
transform 1 0 20944 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_207
timestamp 1698175906
transform 1 0 24528 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_209
timestamp 1698175906
transform 1 0 24752 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_212
timestamp 1698175906
transform 1 0 25088 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_276
timestamp 1698175906
transform 1 0 32256 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_282
timestamp 1698175906
transform 1 0 32928 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_314
timestamp 1698175906
transform 1 0 36512 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_322
timestamp 1698175906
transform 1 0 37408 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_2
timestamp 1698175906
transform 1 0 1568 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698175906
transform 1 0 5152 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_37
timestamp 1698175906
transform 1 0 5488 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_101
timestamp 1698175906
transform 1 0 12656 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_107
timestamp 1698175906
transform 1 0 13328 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_171
timestamp 1698175906
transform 1 0 20496 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_177
timestamp 1698175906
transform 1 0 21168 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_241
timestamp 1698175906
transform 1 0 28336 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_247
timestamp 1698175906
transform 1 0 29008 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_311
timestamp 1698175906
transform 1 0 36176 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_317
timestamp 1698175906
transform 1 0 36848 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_2
timestamp 1698175906
transform 1 0 1568 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_66
timestamp 1698175906
transform 1 0 8736 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_72
timestamp 1698175906
transform 1 0 9408 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_136
timestamp 1698175906
transform 1 0 16576 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_142
timestamp 1698175906
transform 1 0 17248 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_206
timestamp 1698175906
transform 1 0 24416 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_212
timestamp 1698175906
transform 1 0 25088 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_276
timestamp 1698175906
transform 1 0 32256 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_282
timestamp 1698175906
transform 1 0 32928 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_346
timestamp 1698175906
transform 1 0 40096 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_348
timestamp 1698175906
transform 1 0 40320 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698175906
transform 1 0 1568 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698175906
transform 1 0 5152 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_37
timestamp 1698175906
transform 1 0 5488 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_101
timestamp 1698175906
transform 1 0 12656 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_107
timestamp 1698175906
transform 1 0 13328 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_171
timestamp 1698175906
transform 1 0 20496 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_177
timestamp 1698175906
transform 1 0 21168 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_241
timestamp 1698175906
transform 1 0 28336 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_247
timestamp 1698175906
transform 1 0 29008 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_311
timestamp 1698175906
transform 1 0 36176 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_317
timestamp 1698175906
transform 1 0 36848 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2
timestamp 1698175906
transform 1 0 1568 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_66
timestamp 1698175906
transform 1 0 8736 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_72
timestamp 1698175906
transform 1 0 9408 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_136
timestamp 1698175906
transform 1 0 16576 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_142
timestamp 1698175906
transform 1 0 17248 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_206
timestamp 1698175906
transform 1 0 24416 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_212
timestamp 1698175906
transform 1 0 25088 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_276
timestamp 1698175906
transform 1 0 32256 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_282
timestamp 1698175906
transform 1 0 32928 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_346
timestamp 1698175906
transform 1 0 40096 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_348
timestamp 1698175906
transform 1 0 40320 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_2
timestamp 1698175906
transform 1 0 1568 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698175906
transform 1 0 5152 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_37
timestamp 1698175906
transform 1 0 5488 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_101
timestamp 1698175906
transform 1 0 12656 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_107
timestamp 1698175906
transform 1 0 13328 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_171
timestamp 1698175906
transform 1 0 20496 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_177
timestamp 1698175906
transform 1 0 21168 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_241
timestamp 1698175906
transform 1 0 28336 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_247
timestamp 1698175906
transform 1 0 29008 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_311
timestamp 1698175906
transform 1 0 36176 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_317
timestamp 1698175906
transform 1 0 36848 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2
timestamp 1698175906
transform 1 0 1568 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_66
timestamp 1698175906
transform 1 0 8736 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_72
timestamp 1698175906
transform 1 0 9408 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_136
timestamp 1698175906
transform 1 0 16576 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_142
timestamp 1698175906
transform 1 0 17248 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_206
timestamp 1698175906
transform 1 0 24416 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_212
timestamp 1698175906
transform 1 0 25088 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_276
timestamp 1698175906
transform 1 0 32256 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_282
timestamp 1698175906
transform 1 0 32928 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_346
timestamp 1698175906
transform 1 0 40096 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_348
timestamp 1698175906
transform 1 0 40320 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698175906
transform 1 0 1568 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698175906
transform 1 0 5152 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_37
timestamp 1698175906
transform 1 0 5488 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_101
timestamp 1698175906
transform 1 0 12656 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_107
timestamp 1698175906
transform 1 0 13328 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_171
timestamp 1698175906
transform 1 0 20496 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_177
timestamp 1698175906
transform 1 0 21168 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_241
timestamp 1698175906
transform 1 0 28336 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_247
timestamp 1698175906
transform 1 0 29008 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_311
timestamp 1698175906
transform 1 0 36176 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_317
timestamp 1698175906
transform 1 0 36848 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_2
timestamp 1698175906
transform 1 0 1568 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_66
timestamp 1698175906
transform 1 0 8736 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_72
timestamp 1698175906
transform 1 0 9408 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_136
timestamp 1698175906
transform 1 0 16576 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_142
timestamp 1698175906
transform 1 0 17248 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_206
timestamp 1698175906
transform 1 0 24416 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_212
timestamp 1698175906
transform 1 0 25088 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_276
timestamp 1698175906
transform 1 0 32256 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_282
timestamp 1698175906
transform 1 0 32928 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_346
timestamp 1698175906
transform 1 0 40096 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_348
timestamp 1698175906
transform 1 0 40320 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698175906
transform 1 0 1568 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698175906
transform 1 0 5152 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_37
timestamp 1698175906
transform 1 0 5488 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_101
timestamp 1698175906
transform 1 0 12656 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_107
timestamp 1698175906
transform 1 0 13328 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_171
timestamp 1698175906
transform 1 0 20496 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_177
timestamp 1698175906
transform 1 0 21168 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_241
timestamp 1698175906
transform 1 0 28336 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_247
timestamp 1698175906
transform 1 0 29008 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_311
timestamp 1698175906
transform 1 0 36176 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_317
timestamp 1698175906
transform 1 0 36848 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2
timestamp 1698175906
transform 1 0 1568 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1698175906
transform 1 0 8736 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_72
timestamp 1698175906
transform 1 0 9408 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_136
timestamp 1698175906
transform 1 0 16576 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_142
timestamp 1698175906
transform 1 0 17248 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_206
timestamp 1698175906
transform 1 0 24416 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_212
timestamp 1698175906
transform 1 0 25088 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_276
timestamp 1698175906
transform 1 0 32256 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_282
timestamp 1698175906
transform 1 0 32928 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_346
timestamp 1698175906
transform 1 0 40096 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_348
timestamp 1698175906
transform 1 0 40320 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_2
timestamp 1698175906
transform 1 0 1568 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698175906
transform 1 0 5152 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_37
timestamp 1698175906
transform 1 0 5488 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_101
timestamp 1698175906
transform 1 0 12656 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_107
timestamp 1698175906
transform 1 0 13328 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_123
timestamp 1698175906
transform 1 0 15120 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_131
timestamp 1698175906
transform 1 0 16016 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_159
timestamp 1698175906
transform 1 0 19152 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_177
timestamp 1698175906
transform 1 0 21168 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_241
timestamp 1698175906
transform 1 0 28336 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_247
timestamp 1698175906
transform 1 0 29008 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_311
timestamp 1698175906
transform 1 0 36176 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_317
timestamp 1698175906
transform 1 0 36848 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_2
timestamp 1698175906
transform 1 0 1568 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_66
timestamp 1698175906
transform 1 0 8736 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_72
timestamp 1698175906
transform 1 0 9408 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_136
timestamp 1698175906
transform 1 0 16576 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_168
timestamp 1698175906
transform 1 0 20160 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_195
timestamp 1698175906
transform 1 0 23184 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_203
timestamp 1698175906
transform 1 0 24080 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_207
timestamp 1698175906
transform 1 0 24528 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_209
timestamp 1698175906
transform 1 0 24752 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_238
timestamp 1698175906
transform 1 0 28000 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_270
timestamp 1698175906
transform 1 0 31584 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_278
timestamp 1698175906
transform 1 0 32480 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_282
timestamp 1698175906
transform 1 0 32928 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_346
timestamp 1698175906
transform 1 0 40096 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_348
timestamp 1698175906
transform 1 0 40320 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_2
timestamp 1698175906
transform 1 0 1568 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_36
timestamp 1698175906
transform 1 0 5376 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_70
timestamp 1698175906
transform 1 0 9184 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_104
timestamp 1698175906
transform 1 0 12992 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_138
timestamp 1698175906
transform 1 0 16800 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_142
timestamp 1698175906
transform 1 0 17248 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_172
timestamp 1698175906
transform 1 0 20608 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_174
timestamp 1698175906
transform 1 0 20832 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_201
timestamp 1698175906
transform 1 0 23856 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_203
timestamp 1698175906
transform 1 0 24080 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_232
timestamp 1698175906
transform 1 0 27328 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_236
timestamp 1698175906
transform 1 0 27776 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_240
timestamp 1698175906
transform 1 0 28224 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_274
timestamp 1698175906
transform 1 0 32032 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_308
timestamp 1698175906
transform 1 0 35840 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_342
timestamp 1698175906
transform 1 0 39648 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_346
timestamp 1698175906
transform 1 0 40096 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_348
timestamp 1698175906
transform 1 0 40320 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita26_26 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 12656 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 37520 0 -1 28224
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output2
timestamp 1698175906
transform 1 0 37520 0 1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output3
timestamp 1698175906
transform 1 0 37520 0 1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output4
timestamp 1698175906
transform -1 0 4480 0 1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output5
timestamp 1698175906
transform 1 0 37520 0 1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output6
timestamp 1698175906
transform 1 0 20944 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output7
timestamp 1698175906
transform 1 0 37520 0 1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output8
timestamp 1698175906
transform 1 0 37520 0 1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output9
timestamp 1698175906
transform 1 0 20272 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output10
timestamp 1698175906
transform 1 0 37520 0 -1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output11
timestamp 1698175906
transform -1 0 4480 0 1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output12
timestamp 1698175906
transform 1 0 24416 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output13
timestamp 1698175906
transform -1 0 4480 0 1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output14
timestamp 1698175906
transform 1 0 24416 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output15
timestamp 1698175906
transform -1 0 4480 0 -1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output16
timestamp 1698175906
transform 1 0 37520 0 -1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output17
timestamp 1698175906
transform -1 0 20384 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output18
timestamp 1698175906
transform 1 0 37520 0 -1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output19
timestamp 1698175906
transform 1 0 26992 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output20
timestamp 1698175906
transform 1 0 25088 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output21
timestamp 1698175906
transform 1 0 37520 0 -1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output22
timestamp 1698175906
transform 1 0 37520 0 -1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output23
timestamp 1698175906
transform 1 0 17248 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output24
timestamp 1698175906
transform 1 0 16240 0 1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output25
timestamp 1698175906
transform -1 0 4480 0 -1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_45 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698175906
transform -1 0 40656 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_46
timestamp 1698175906
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698175906
transform -1 0 40656 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_47
timestamp 1698175906
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698175906
transform -1 0 40656 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_48
timestamp 1698175906
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698175906
transform -1 0 40656 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_49
timestamp 1698175906
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698175906
transform -1 0 40656 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_50
timestamp 1698175906
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698175906
transform -1 0 40656 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_51
timestamp 1698175906
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698175906
transform -1 0 40656 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_52
timestamp 1698175906
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698175906
transform -1 0 40656 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_53
timestamp 1698175906
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698175906
transform -1 0 40656 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_54
timestamp 1698175906
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698175906
transform -1 0 40656 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_55
timestamp 1698175906
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698175906
transform -1 0 40656 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_56
timestamp 1698175906
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698175906
transform -1 0 40656 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_57
timestamp 1698175906
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698175906
transform -1 0 40656 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_58
timestamp 1698175906
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698175906
transform -1 0 40656 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_59
timestamp 1698175906
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698175906
transform -1 0 40656 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_60
timestamp 1698175906
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698175906
transform -1 0 40656 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_61
timestamp 1698175906
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698175906
transform -1 0 40656 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_62
timestamp 1698175906
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698175906
transform -1 0 40656 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_63
timestamp 1698175906
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698175906
transform -1 0 40656 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_64
timestamp 1698175906
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698175906
transform -1 0 40656 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_65
timestamp 1698175906
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698175906
transform -1 0 40656 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_66
timestamp 1698175906
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698175906
transform -1 0 40656 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_67
timestamp 1698175906
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698175906
transform -1 0 40656 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_68
timestamp 1698175906
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698175906
transform -1 0 40656 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_69
timestamp 1698175906
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698175906
transform -1 0 40656 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_70
timestamp 1698175906
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698175906
transform -1 0 40656 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_71
timestamp 1698175906
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698175906
transform -1 0 40656 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_72
timestamp 1698175906
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698175906
transform -1 0 40656 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_73
timestamp 1698175906
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698175906
transform -1 0 40656 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_74
timestamp 1698175906
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698175906
transform -1 0 40656 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_75
timestamp 1698175906
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698175906
transform -1 0 40656 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_76
timestamp 1698175906
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698175906
transform -1 0 40656 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_77
timestamp 1698175906
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698175906
transform -1 0 40656 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_78
timestamp 1698175906
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698175906
transform -1 0 40656 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_79
timestamp 1698175906
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698175906
transform -1 0 40656 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_80
timestamp 1698175906
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698175906
transform -1 0 40656 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_81
timestamp 1698175906
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698175906
transform -1 0 40656 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_82
timestamp 1698175906
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698175906
transform -1 0 40656 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_83
timestamp 1698175906
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698175906
transform -1 0 40656 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_84
timestamp 1698175906
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698175906
transform -1 0 40656 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_85
timestamp 1698175906
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698175906
transform -1 0 40656 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_86
timestamp 1698175906
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698175906
transform -1 0 40656 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_87
timestamp 1698175906
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698175906
transform -1 0 40656 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_88
timestamp 1698175906
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698175906
transform -1 0 40656 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_89
timestamp 1698175906
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698175906
transform -1 0 40656 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_90 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_91
timestamp 1698175906
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_92
timestamp 1698175906
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_93
timestamp 1698175906
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_94
timestamp 1698175906
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_95
timestamp 1698175906
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_96
timestamp 1698175906
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_97
timestamp 1698175906
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_98
timestamp 1698175906
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_99
timestamp 1698175906
transform 1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_100
timestamp 1698175906
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_101
timestamp 1698175906
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_102
timestamp 1698175906
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_103
timestamp 1698175906
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_104
timestamp 1698175906
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_105
timestamp 1698175906
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_106
timestamp 1698175906
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_107
timestamp 1698175906
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_108
timestamp 1698175906
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_109
timestamp 1698175906
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_110
timestamp 1698175906
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_111
timestamp 1698175906
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_112
timestamp 1698175906
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_113
timestamp 1698175906
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_114
timestamp 1698175906
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_115
timestamp 1698175906
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_116
timestamp 1698175906
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_117
timestamp 1698175906
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_118
timestamp 1698175906
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_119
timestamp 1698175906
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_120
timestamp 1698175906
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_121
timestamp 1698175906
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_122
timestamp 1698175906
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_123
timestamp 1698175906
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_124
timestamp 1698175906
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_125
timestamp 1698175906
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_126
timestamp 1698175906
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_127
timestamp 1698175906
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_128
timestamp 1698175906
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_129
timestamp 1698175906
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_130
timestamp 1698175906
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_131
timestamp 1698175906
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_132
timestamp 1698175906
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_133
timestamp 1698175906
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_134
timestamp 1698175906
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_135
timestamp 1698175906
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_136
timestamp 1698175906
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_137
timestamp 1698175906
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_138
timestamp 1698175906
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_139
timestamp 1698175906
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_140
timestamp 1698175906
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_141
timestamp 1698175906
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_142
timestamp 1698175906
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_143
timestamp 1698175906
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_144
timestamp 1698175906
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_145
timestamp 1698175906
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_146
timestamp 1698175906
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_147
timestamp 1698175906
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_148
timestamp 1698175906
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_149
timestamp 1698175906
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_150
timestamp 1698175906
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_151
timestamp 1698175906
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_152
timestamp 1698175906
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_153
timestamp 1698175906
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_154
timestamp 1698175906
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_155
timestamp 1698175906
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_156
timestamp 1698175906
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_157
timestamp 1698175906
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_158
timestamp 1698175906
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_159
timestamp 1698175906
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_160
timestamp 1698175906
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_161
timestamp 1698175906
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_162
timestamp 1698175906
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_163
timestamp 1698175906
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_164
timestamp 1698175906
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_165
timestamp 1698175906
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_166
timestamp 1698175906
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_167
timestamp 1698175906
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_168
timestamp 1698175906
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_169
timestamp 1698175906
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_170
timestamp 1698175906
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_171
timestamp 1698175906
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_172
timestamp 1698175906
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_173
timestamp 1698175906
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_174
timestamp 1698175906
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_175
timestamp 1698175906
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_176
timestamp 1698175906
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_177
timestamp 1698175906
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_178
timestamp 1698175906
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_179
timestamp 1698175906
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_180
timestamp 1698175906
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_181
timestamp 1698175906
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_182
timestamp 1698175906
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_183
timestamp 1698175906
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_184
timestamp 1698175906
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_185
timestamp 1698175906
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_186
timestamp 1698175906
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_187
timestamp 1698175906
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_188
timestamp 1698175906
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_189
timestamp 1698175906
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_190
timestamp 1698175906
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_191
timestamp 1698175906
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_192
timestamp 1698175906
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_193
timestamp 1698175906
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_194
timestamp 1698175906
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_195
timestamp 1698175906
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_196
timestamp 1698175906
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_197
timestamp 1698175906
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_198
timestamp 1698175906
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_199
timestamp 1698175906
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_200
timestamp 1698175906
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_201
timestamp 1698175906
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_202
timestamp 1698175906
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_203
timestamp 1698175906
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_204
timestamp 1698175906
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_205
timestamp 1698175906
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_206
timestamp 1698175906
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_207
timestamp 1698175906
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_208
timestamp 1698175906
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_209
timestamp 1698175906
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_210
timestamp 1698175906
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_211
timestamp 1698175906
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_212
timestamp 1698175906
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_213
timestamp 1698175906
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_214
timestamp 1698175906
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_215
timestamp 1698175906
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_216
timestamp 1698175906
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_217
timestamp 1698175906
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_218
timestamp 1698175906
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_219
timestamp 1698175906
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_220
timestamp 1698175906
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_221
timestamp 1698175906
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_222
timestamp 1698175906
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_223
timestamp 1698175906
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_224
timestamp 1698175906
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_225
timestamp 1698175906
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_226
timestamp 1698175906
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_227
timestamp 1698175906
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_228
timestamp 1698175906
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_229
timestamp 1698175906
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_230
timestamp 1698175906
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_231
timestamp 1698175906
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_232
timestamp 1698175906
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_233
timestamp 1698175906
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_234
timestamp 1698175906
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_235
timestamp 1698175906
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_236
timestamp 1698175906
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_237
timestamp 1698175906
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_238
timestamp 1698175906
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_239
timestamp 1698175906
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_240
timestamp 1698175906
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_241
timestamp 1698175906
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_242
timestamp 1698175906
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_243
timestamp 1698175906
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_244
timestamp 1698175906
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_245
timestamp 1698175906
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_246
timestamp 1698175906
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_247
timestamp 1698175906
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_248
timestamp 1698175906
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_249
timestamp 1698175906
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_250
timestamp 1698175906
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_251
timestamp 1698175906
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_252
timestamp 1698175906
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_253
timestamp 1698175906
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_254
timestamp 1698175906
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_255
timestamp 1698175906
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_256
timestamp 1698175906
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_257
timestamp 1698175906
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_258
timestamp 1698175906
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_259
timestamp 1698175906
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_260
timestamp 1698175906
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_261
timestamp 1698175906
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_262
timestamp 1698175906
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_263
timestamp 1698175906
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_264
timestamp 1698175906
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_265
timestamp 1698175906
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_266
timestamp 1698175906
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_267
timestamp 1698175906
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_268
timestamp 1698175906
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_269
timestamp 1698175906
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_270
timestamp 1698175906
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_271
timestamp 1698175906
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_272
timestamp 1698175906
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_273
timestamp 1698175906
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_274
timestamp 1698175906
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_275
timestamp 1698175906
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_276
timestamp 1698175906
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_277
timestamp 1698175906
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_278
timestamp 1698175906
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_279
timestamp 1698175906
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_280
timestamp 1698175906
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_281
timestamp 1698175906
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_282
timestamp 1698175906
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_283
timestamp 1698175906
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_284
timestamp 1698175906
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_285
timestamp 1698175906
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_286
timestamp 1698175906
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_287
timestamp 1698175906
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_288
timestamp 1698175906
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_289
timestamp 1698175906
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_290
timestamp 1698175906
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_291
timestamp 1698175906
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_292
timestamp 1698175906
transform 1 0 32704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_293
timestamp 1698175906
transform 1 0 5152 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_294
timestamp 1698175906
transform 1 0 8960 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_295
timestamp 1698175906
transform 1 0 12768 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_296
timestamp 1698175906
transform 1 0 16576 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_297
timestamp 1698175906
transform 1 0 20384 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_298
timestamp 1698175906
transform 1 0 24192 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_299
timestamp 1698175906
transform 1 0 28000 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_300
timestamp 1698175906
transform 1 0 31808 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_301
timestamp 1698175906
transform 1 0 35616 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_302
timestamp 1698175906
transform 1 0 39424 0 1 37632
box -86 -86 310 870
<< labels >>
flabel metal3 s 0 26880 800 26992 0 FreeSans 448 0 0 0 clk
port 0 nsew signal input
flabel metal3 s 41200 27552 42000 27664 0 FreeSans 448 0 0 0 segm[0]
port 1 nsew signal tristate
flabel metal3 s 41200 23520 42000 23632 0 FreeSans 448 0 0 0 segm[10]
port 2 nsew signal tristate
flabel metal3 s 41200 21504 42000 21616 0 FreeSans 448 0 0 0 segm[11]
port 3 nsew signal tristate
flabel metal3 s 0 20160 800 20272 0 FreeSans 448 0 0 0 segm[12]
port 4 nsew signal tristate
flabel metal3 s 41200 17472 42000 17584 0 FreeSans 448 0 0 0 segm[13]
port 5 nsew signal tristate
flabel metal2 s 20832 41200 20944 42000 0 FreeSans 448 90 0 0 segm[1]
port 6 nsew signal tristate
flabel metal3 s 41200 20160 42000 20272 0 FreeSans 448 0 0 0 segm[2]
port 7 nsew signal tristate
flabel metal3 s 41200 26208 42000 26320 0 FreeSans 448 0 0 0 segm[3]
port 8 nsew signal tristate
flabel metal2 s 20160 41200 20272 42000 0 FreeSans 448 90 0 0 segm[4]
port 9 nsew signal tristate
flabel metal2 s 12096 0 12208 800 0 FreeSans 448 90 0 0 segm[5]
port 10 nsew signal tristate
flabel metal3 s 41200 22848 42000 22960 0 FreeSans 448 0 0 0 segm[6]
port 11 nsew signal tristate
flabel metal3 s 0 23520 800 23632 0 FreeSans 448 0 0 0 segm[7]
port 12 nsew signal tristate
flabel metal2 s 23520 41200 23632 42000 0 FreeSans 448 90 0 0 segm[8]
port 13 nsew signal tristate
flabel metal3 s 0 17472 800 17584 0 FreeSans 448 0 0 0 segm[9]
port 14 nsew signal tristate
flabel metal2 s 24192 0 24304 800 0 FreeSans 448 90 0 0 sel[0]
port 15 nsew signal tristate
flabel metal3 s 0 22848 800 22960 0 FreeSans 448 0 0 0 sel[10]
port 16 nsew signal tristate
flabel metal3 s 41200 18144 42000 18256 0 FreeSans 448 0 0 0 sel[11]
port 17 nsew signal tristate
flabel metal2 s 19488 41200 19600 42000 0 FreeSans 448 90 0 0 sel[1]
port 18 nsew signal tristate
flabel metal3 s 41200 20832 42000 20944 0 FreeSans 448 0 0 0 sel[2]
port 19 nsew signal tristate
flabel metal2 s 26880 0 26992 800 0 FreeSans 448 90 0 0 sel[3]
port 20 nsew signal tristate
flabel metal2 s 24192 41200 24304 42000 0 FreeSans 448 90 0 0 sel[4]
port 21 nsew signal tristate
flabel metal3 s 41200 26880 42000 26992 0 FreeSans 448 0 0 0 sel[5]
port 22 nsew signal tristate
flabel metal3 s 41200 16800 42000 16912 0 FreeSans 448 0 0 0 sel[6]
port 23 nsew signal tristate
flabel metal2 s 16800 41200 16912 42000 0 FreeSans 448 90 0 0 sel[7]
port 24 nsew signal tristate
flabel metal2 s 16128 41200 16240 42000 0 FreeSans 448 90 0 0 sel[8]
port 25 nsew signal tristate
flabel metal3 s 0 19488 800 19600 0 FreeSans 448 0 0 0 sel[9]
port 26 nsew signal tristate
flabel metal4 s 4448 3076 4768 38476 0 FreeSans 1280 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 35168 3076 35488 38476 0 FreeSans 1280 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 19808 3076 20128 38476 0 FreeSans 1280 90 0 0 vss
port 28 nsew ground bidirectional
rlabel metal1 21000 38416 21000 38416 0 vdd
rlabel metal1 21000 37632 21000 37632 0 vss
rlabel metal2 26600 17808 26600 17808 0 _000_
rlabel metal2 16296 26936 16296 26936 0 _001_
rlabel metal2 22792 27384 22792 27384 0 _002_
rlabel metal2 16632 16968 16632 16968 0 _003_
rlabel metal2 14392 15624 14392 15624 0 _004_
rlabel metal2 19600 13832 19600 13832 0 _005_
rlabel metal2 18088 22008 18088 22008 0 _006_
rlabel metal2 25760 14616 25760 14616 0 _007_
rlabel metal2 14952 25592 14952 25592 0 _008_
rlabel metal2 27384 19824 27384 19824 0 _009_
rlabel metal2 18200 27384 18200 27384 0 _010_
rlabel metal2 22848 14392 22848 14392 0 _011_
rlabel metal2 13496 16352 13496 16352 0 _012_
rlabel metal2 14280 20832 14280 20832 0 _013_
rlabel metal2 23856 16184 23856 16184 0 _014_
rlabel metal2 25312 26936 25312 26936 0 _015_
rlabel metal2 13496 22848 13496 22848 0 _016_
rlabel metal2 27720 18032 27720 18032 0 _017_
rlabel metal2 19096 25144 19096 25144 0 _018_
rlabel metal2 26264 22736 26264 22736 0 _019_
rlabel metal2 13944 22624 13944 22624 0 _020_
rlabel metal2 21560 24136 21560 24136 0 _021_
rlabel metal2 26376 23744 26376 23744 0 _022_
rlabel metal2 23352 22008 23352 22008 0 _023_
rlabel metal2 12152 19600 12152 19600 0 _024_
rlabel metal2 15512 27832 15512 27832 0 _025_
rlabel metal2 27720 22344 27720 22344 0 _026_
rlabel metal2 26600 19600 26600 19600 0 _027_
rlabel metal2 14840 17920 14840 17920 0 _028_
rlabel metal3 17640 23688 17640 23688 0 _029_
rlabel metal2 18312 25480 18312 25480 0 _030_
rlabel metal2 18648 26936 18648 26936 0 _031_
rlabel metal2 20608 15512 20608 15512 0 _032_
rlabel metal2 23352 15204 23352 15204 0 _033_
rlabel metal2 15456 17640 15456 17640 0 _034_
rlabel metal2 18312 18256 18312 18256 0 _035_
rlabel metal2 14280 18256 14280 18256 0 _036_
rlabel metal2 14952 18088 14952 18088 0 _037_
rlabel metal2 13832 16352 13832 16352 0 _038_
rlabel metal2 14280 20440 14280 20440 0 _039_
rlabel metal2 14504 19712 14504 19712 0 _040_
rlabel metal2 14616 20384 14616 20384 0 _041_
rlabel metal2 14840 20888 14840 20888 0 _042_
rlabel metal2 25704 16800 25704 16800 0 _043_
rlabel metal2 23464 17416 23464 17416 0 _044_
rlabel metal2 23800 17752 23800 17752 0 _045_
rlabel metal2 24584 25648 24584 25648 0 _046_
rlabel metal2 25592 26264 25592 26264 0 _047_
rlabel metal3 19936 23800 19936 23800 0 _048_
rlabel metal2 21224 20888 21224 20888 0 _049_
rlabel metal2 15064 23576 15064 23576 0 _050_
rlabel metal3 28392 17528 28392 17528 0 _051_
rlabel metal2 19488 24920 19488 24920 0 _052_
rlabel metal2 19824 24024 19824 24024 0 _053_
rlabel metal2 24024 21616 24024 21616 0 _054_
rlabel metal3 26936 22344 26936 22344 0 _055_
rlabel metal2 25592 21840 25592 21840 0 _056_
rlabel metal2 15848 21840 15848 21840 0 _057_
rlabel metal2 16520 23408 16520 23408 0 _058_
rlabel metal2 15176 22680 15176 22680 0 _059_
rlabel metal2 13720 22176 13720 22176 0 _060_
rlabel metal2 22792 23912 22792 23912 0 _061_
rlabel metal2 26936 22456 26936 22456 0 _062_
rlabel metal2 24248 20496 24248 20496 0 _063_
rlabel metal3 14532 19992 14532 19992 0 _064_
rlabel metal3 19208 19768 19208 19768 0 _065_
rlabel metal2 19656 18144 19656 18144 0 _066_
rlabel metal2 27272 18088 27272 18088 0 _067_
rlabel metal3 18088 16072 18088 16072 0 _068_
rlabel metal2 15848 15848 15848 15848 0 _069_
rlabel metal2 28280 17976 28280 17976 0 _070_
rlabel metal2 20776 15680 20776 15680 0 _071_
rlabel metal3 21224 20104 21224 20104 0 _072_
rlabel metal2 26320 18424 26320 18424 0 _073_
rlabel metal2 19432 14336 19432 14336 0 _074_
rlabel metal2 17528 16912 17528 16912 0 _075_
rlabel metal2 14392 20356 14392 20356 0 _076_
rlabel metal3 16744 21560 16744 21560 0 _077_
rlabel metal2 17528 22512 17528 22512 0 _078_
rlabel metal2 23240 19600 23240 19600 0 _079_
rlabel metal2 23352 27048 23352 27048 0 _080_
rlabel metal3 17136 26936 17136 26936 0 _081_
rlabel metal2 23912 21672 23912 21672 0 _082_
rlabel metal2 19656 23128 19656 23128 0 _083_
rlabel metal2 22120 21840 22120 21840 0 _084_
rlabel metal2 22904 26264 22904 26264 0 _085_
rlabel metal2 23352 27272 23352 27272 0 _086_
rlabel metal2 19880 15960 19880 15960 0 _087_
rlabel metal2 18648 17192 18648 17192 0 _088_
rlabel metal2 15848 16464 15848 16464 0 _089_
rlabel metal2 27160 16352 27160 16352 0 _090_
rlabel metal3 18536 19096 18536 19096 0 _091_
rlabel metal2 18592 19208 18592 19208 0 _092_
rlabel metal2 24360 19600 24360 19600 0 _093_
rlabel metal2 20552 19152 20552 19152 0 _094_
rlabel metal2 15064 18704 15064 18704 0 _095_
rlabel metal3 18872 18424 18872 18424 0 _096_
rlabel metal2 19544 18424 19544 18424 0 _097_
rlabel metal2 19376 19992 19376 19992 0 _098_
rlabel metal2 25816 15204 25816 15204 0 _099_
rlabel metal3 18312 18312 18312 18312 0 _100_
rlabel metal3 24024 15288 24024 15288 0 _101_
rlabel metal2 18424 19320 18424 19320 0 _102_
rlabel metal2 16744 20048 16744 20048 0 _103_
rlabel metal2 15848 20888 15848 20888 0 _104_
rlabel metal2 15512 22624 15512 22624 0 _105_
rlabel metal3 2478 26936 2478 26936 0 clk
rlabel metal2 25144 20412 25144 20412 0 clknet_0_clk
rlabel metal2 27048 20356 27048 20356 0 clknet_1_0__leaf_clk
rlabel metal2 21448 27776 21448 27776 0 clknet_1_1__leaf_clk
rlabel metal2 18312 13664 18312 13664 0 dut26.count\[0\]
rlabel metal2 16296 16408 16296 16408 0 dut26.count\[1\]
rlabel metal2 21728 16072 21728 16072 0 dut26.count\[2\]
rlabel metal2 20384 21000 20384 21000 0 dut26.count\[3\]
rlabel metal2 37912 27384 37912 27384 0 net1
rlabel metal2 27832 22120 27832 22120 0 net10
rlabel metal2 12040 23464 12040 23464 0 net11
rlabel metal2 24192 31920 24192 31920 0 net12
rlabel metal2 11480 17584 11480 17584 0 net13
rlabel metal2 24696 14560 24696 14560 0 net14
rlabel metal2 11368 22288 11368 22288 0 net15
rlabel metal2 29288 18032 29288 18032 0 net16
rlabel metal2 18984 27328 18984 27328 0 net17
rlabel metal3 34048 20104 34048 20104 0 net18
rlabel metal2 27944 14112 27944 14112 0 net19
rlabel metal2 27160 23128 27160 23128 0 net2
rlabel metal3 24808 27720 24808 27720 0 net20
rlabel metal3 29540 26376 29540 26376 0 net21
rlabel metal2 29176 16800 29176 16800 0 net22
rlabel metal2 17528 27160 17528 27160 0 net23
rlabel metal2 15960 29988 15960 29988 0 net24
rlabel metal3 6356 19992 6356 19992 0 net25
rlabel metal2 12152 2030 12152 2030 0 net26
rlabel metal3 31920 22400 31920 22400 0 net3
rlabel metal3 6356 20776 6356 20776 0 net4
rlabel metal2 25592 17360 25592 17360 0 net5
rlabel metal2 20664 38024 20664 38024 0 net6
rlabel metal2 29512 19488 29512 19488 0 net7
rlabel metal2 27608 27104 27608 27104 0 net8
rlabel metal2 20440 27160 20440 27160 0 net9
rlabel metal3 40642 27608 40642 27608 0 segm[0]
rlabel metal2 40040 23800 40040 23800 0 segm[10]
rlabel metal2 40040 22008 40040 22008 0 segm[11]
rlabel metal3 1358 20216 1358 20216 0 segm[12]
rlabel metal2 40040 17640 40040 17640 0 segm[13]
rlabel metal2 20888 39746 20888 39746 0 segm[1]
rlabel metal2 40040 20552 40040 20552 0 segm[2]
rlabel metal2 40040 26712 40040 26712 0 segm[3]
rlabel metal2 20216 39914 20216 39914 0 segm[4]
rlabel metal3 40642 22904 40642 22904 0 segm[6]
rlabel metal3 1358 23576 1358 23576 0 segm[7]
rlabel metal2 23576 39746 23576 39746 0 segm[8]
rlabel metal3 1358 17528 1358 17528 0 segm[9]
rlabel metal3 24920 3640 24920 3640 0 sel[0]
rlabel metal3 1358 22904 1358 22904 0 sel[10]
rlabel metal3 40642 18200 40642 18200 0 sel[11]
rlabel metal2 19544 39746 19544 39746 0 sel[1]
rlabel metal2 39928 21168 39928 21168 0 sel[2]
rlabel metal2 26936 2422 26936 2422 0 sel[3]
rlabel metal2 24248 39354 24248 39354 0 sel[4]
rlabel metal2 39928 26488 39928 26488 0 sel[5]
rlabel metal2 40040 16800 40040 16800 0 sel[6]
rlabel metal2 16856 39354 16856 39354 0 sel[7]
rlabel metal2 16184 38962 16184 38962 0 sel[8]
rlabel metal3 1358 19544 1358 19544 0 sel[9]
<< properties >>
string FIXED_BBOX 0 0 42000 42000
<< end >>
