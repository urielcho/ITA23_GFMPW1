* NGSPICE file created from user_project_wrapper.ext - technology: gf180mcuD

* Black-box entry subcircuit for ita60 abstract view
.subckt ita60 clk segm[0] segm[10] segm[11] segm[12] segm[13] segm[1] segm[2] segm[3]
+ segm[4] segm[5] segm[6] segm[7] segm[8] segm[9] sel[0] sel[10] sel[11] sel[1] sel[2]
+ sel[3] sel[4] sel[5] sel[6] sel[7] sel[8] sel[9] vdd vss
.ends

* Black-box entry subcircuit for ita1 abstract view
.subckt ita1 clk segm[0] segm[10] segm[11] segm[12] segm[13] segm[1] segm[2] segm[3]
+ segm[4] segm[5] segm[6] segm[7] segm[8] segm[9] sel[0] sel[10] sel[11] sel[1] sel[2]
+ sel[3] sel[4] sel[5] sel[6] sel[7] sel[8] sel[9] vdd vss
.ends

* Black-box entry subcircuit for ita61 abstract view
.subckt ita61 clk segm[0] segm[10] segm[11] segm[12] segm[13] segm[1] segm[2] segm[3]
+ segm[4] segm[5] segm[6] segm[7] segm[8] segm[9] sel[0] sel[10] sel[11] sel[1] sel[2]
+ sel[3] sel[4] sel[5] sel[6] sel[7] sel[8] sel[9] vdd vss
.ends

* Black-box entry subcircuit for ita50 abstract view
.subckt ita50 clk segm[0] segm[10] segm[11] segm[12] segm[13] segm[1] segm[2] segm[3]
+ segm[4] segm[5] segm[6] segm[7] segm[8] segm[9] sel[0] sel[10] sel[11] sel[1] sel[2]
+ sel[3] sel[4] sel[5] sel[6] sel[7] sel[8] sel[9] vdd vss
.ends

* Black-box entry subcircuit for ita2 abstract view
.subckt ita2 clk segm[0] segm[10] segm[11] segm[12] segm[13] segm[1] segm[2] segm[3]
+ segm[4] segm[5] segm[6] segm[7] segm[8] segm[9] sel[0] sel[10] sel[11] sel[1] sel[2]
+ sel[3] sel[4] sel[5] sel[6] sel[7] sel[8] sel[9] vdd vss
.ends

* Black-box entry subcircuit for ita40 abstract view
.subckt ita40 clk segm[0] segm[10] segm[11] segm[12] segm[13] segm[1] segm[2] segm[3]
+ segm[4] segm[5] segm[6] segm[7] segm[8] segm[9] sel[0] sel[10] sel[11] sel[1] sel[2]
+ sel[3] sel[4] sel[5] sel[6] sel[7] sel[8] sel[9] vdd vss
.ends

* Black-box entry subcircuit for ita62 abstract view
.subckt ita62 clk segm[0] segm[10] segm[11] segm[12] segm[13] segm[1] segm[2] segm[3]
+ segm[4] segm[5] segm[6] segm[7] segm[8] segm[9] sel[0] sel[10] sel[11] sel[1] sel[2]
+ sel[3] sel[4] sel[5] sel[6] sel[7] sel[8] sel[9] vdd vss
.ends

* Black-box entry subcircuit for ita4 abstract view
.subckt ita4 clk segm[0] segm[10] segm[11] segm[12] segm[13] segm[1] segm[2] segm[3]
+ segm[4] segm[5] segm[6] segm[7] segm[8] segm[9] sel[0] sel[10] sel[11] sel[1] sel[2]
+ sel[3] sel[4] sel[5] sel[6] sel[7] sel[8] sel[9] vdd vss
.ends

* Black-box entry subcircuit for ita51 abstract view
.subckt ita51 clk segm[0] segm[10] segm[11] segm[12] segm[13] segm[1] segm[2] segm[3]
+ segm[4] segm[5] segm[6] segm[7] segm[8] segm[9] sel[0] sel[10] sel[11] sel[1] sel[2]
+ sel[3] sel[4] sel[5] sel[6] sel[7] sel[8] sel[9] vdd vss
.ends

* Black-box entry subcircuit for ita3 abstract view
.subckt ita3 clk segm[0] segm[10] segm[11] segm[12] segm[13] segm[1] segm[2] segm[3]
+ segm[4] segm[5] segm[6] segm[7] segm[8] segm[9] sel[0] sel[10] sel[11] sel[1] sel[2]
+ sel[3] sel[4] sel[5] sel[6] sel[7] sel[8] sel[9] vdd vss
.ends

* Black-box entry subcircuit for ita63 abstract view
.subckt ita63 clk segm[0] segm[10] segm[11] segm[12] segm[13] segm[1] segm[2] segm[3]
+ segm[4] segm[5] segm[6] segm[7] segm[8] segm[9] sel[0] sel[10] sel[11] sel[1] sel[2]
+ sel[3] sel[4] sel[5] sel[6] sel[7] sel[8] sel[9] vdd vss
.ends

* Black-box entry subcircuit for ita30 abstract view
.subckt ita30 clk segm[0] segm[10] segm[11] segm[12] segm[13] segm[1] segm[2] segm[3]
+ segm[4] segm[5] segm[6] segm[7] segm[8] segm[9] sel[0] sel[10] sel[11] sel[1] sel[2]
+ sel[3] sel[4] sel[5] sel[6] sel[7] sel[8] sel[9] vdd vss
.ends

* Black-box entry subcircuit for ita5 abstract view
.subckt ita5 clk segm[0] segm[10] segm[11] segm[12] segm[13] segm[1] segm[2] segm[3]
+ segm[4] segm[5] segm[6] segm[7] segm[8] segm[9] sel[0] sel[10] sel[11] sel[1] sel[2]
+ sel[3] sel[4] sel[5] sel[6] sel[7] sel[8] sel[9] vdd vss
.ends

* Black-box entry subcircuit for ita52 abstract view
.subckt ita52 clk segm[0] segm[10] segm[11] segm[12] segm[13] segm[1] segm[2] segm[3]
+ segm[4] segm[5] segm[6] segm[7] segm[8] segm[9] sel[0] sel[10] sel[11] sel[1] sel[2]
+ sel[3] sel[4] sel[5] sel[6] sel[7] sel[8] sel[9] vdd vss
.ends

* Black-box entry subcircuit for ita41 abstract view
.subckt ita41 clk segm[0] segm[10] segm[11] segm[12] segm[13] segm[1] segm[2] segm[3]
+ segm[4] segm[5] segm[6] segm[7] segm[8] segm[9] sel[0] sel[10] sel[11] sel[1] sel[2]
+ sel[3] sel[4] sel[5] sel[6] sel[7] sel[8] sel[9] vdd vss
.ends

* Black-box entry subcircuit for ita64 abstract view
.subckt ita64 clk segm[0] segm[10] segm[11] segm[12] segm[13] segm[1] segm[2] segm[3]
+ segm[4] segm[5] segm[6] segm[7] segm[8] segm[9] sel[0] sel[10] sel[11] sel[1] sel[2]
+ sel[3] sel[4] sel[5] sel[6] sel[7] sel[8] sel[9] vdd vss
.ends

* Black-box entry subcircuit for ita31 abstract view
.subckt ita31 clk segm[0] segm[10] segm[11] segm[12] segm[13] segm[1] segm[2] segm[3]
+ segm[4] segm[5] segm[6] segm[7] segm[8] segm[9] sel[0] sel[10] sel[11] sel[1] sel[2]
+ sel[3] sel[4] sel[5] sel[6] sel[7] sel[8] sel[9] vdd vss
.ends

* Black-box entry subcircuit for ita6 abstract view
.subckt ita6 clk segm[0] segm[10] segm[11] segm[12] segm[13] segm[1] segm[2] segm[3]
+ segm[4] segm[5] segm[6] segm[7] segm[8] segm[9] sel[0] sel[10] sel[11] sel[1] sel[2]
+ sel[3] sel[4] sel[5] sel[6] sel[7] sel[8] sel[9] vdd vss
.ends

* Black-box entry subcircuit for ita53 abstract view
.subckt ita53 clk segm[0] segm[10] segm[11] segm[12] segm[13] segm[1] segm[2] segm[3]
+ segm[4] segm[5] segm[6] segm[7] segm[8] segm[9] sel[0] sel[10] sel[11] sel[1] sel[2]
+ sel[3] sel[4] sel[5] sel[6] sel[7] sel[8] sel[9] vdd vss
.ends

* Black-box entry subcircuit for ita abstract view
.subckt ita clk io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14] io_oeb[15]
+ io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21] io_oeb[22]
+ io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27] io_oeb[28] io_oeb[29] io_oeb[2]
+ io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34] io_oeb[35] io_oeb[36] io_oeb[37]
+ io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9] itasegm[0]
+ itasegm[100] itasegm[101] itasegm[102] itasegm[103] itasegm[104] itasegm[105] itasegm[106]
+ itasegm[107] itasegm[108] itasegm[109] itasegm[10] itasegm[110] itasegm[111] itasegm[112]
+ itasegm[113] itasegm[114] itasegm[115] itasegm[116] itasegm[117] itasegm[118] itasegm[119]
+ itasegm[11] itasegm[120] itasegm[121] itasegm[122] itasegm[123] itasegm[124] itasegm[125]
+ itasegm[126] itasegm[127] itasegm[128] itasegm[129] itasegm[12] itasegm[130] itasegm[131]
+ itasegm[132] itasegm[133] itasegm[134] itasegm[135] itasegm[136] itasegm[137] itasegm[138]
+ itasegm[139] itasegm[13] itasegm[140] itasegm[141] itasegm[142] itasegm[143] itasegm[144]
+ itasegm[145] itasegm[146] itasegm[147] itasegm[148] itasegm[149] itasegm[14] itasegm[150]
+ itasegm[151] itasegm[152] itasegm[153] itasegm[154] itasegm[155] itasegm[156] itasegm[157]
+ itasegm[158] itasegm[159] itasegm[15] itasegm[160] itasegm[161] itasegm[162] itasegm[163]
+ itasegm[164] itasegm[165] itasegm[166] itasegm[167] itasegm[168] itasegm[169] itasegm[16]
+ itasegm[170] itasegm[171] itasegm[172] itasegm[173] itasegm[174] itasegm[175] itasegm[176]
+ itasegm[177] itasegm[178] itasegm[179] itasegm[17] itasegm[180] itasegm[181] itasegm[182]
+ itasegm[183] itasegm[184] itasegm[185] itasegm[186] itasegm[187] itasegm[188] itasegm[189]
+ itasegm[18] itasegm[190] itasegm[191] itasegm[192] itasegm[193] itasegm[194] itasegm[195]
+ itasegm[196] itasegm[197] itasegm[198] itasegm[199] itasegm[19] itasegm[1] itasegm[200]
+ itasegm[201] itasegm[202] itasegm[203] itasegm[204] itasegm[205] itasegm[206] itasegm[207]
+ itasegm[208] itasegm[209] itasegm[20] itasegm[210] itasegm[211] itasegm[212] itasegm[213]
+ itasegm[214] itasegm[215] itasegm[216] itasegm[217] itasegm[218] itasegm[219] itasegm[21]
+ itasegm[220] itasegm[221] itasegm[222] itasegm[223] itasegm[224] itasegm[225] itasegm[226]
+ itasegm[227] itasegm[228] itasegm[229] itasegm[22] itasegm[230] itasegm[231] itasegm[232]
+ itasegm[233] itasegm[234] itasegm[235] itasegm[236] itasegm[237] itasegm[238] itasegm[239]
+ itasegm[23] itasegm[240] itasegm[241] itasegm[242] itasegm[243] itasegm[244] itasegm[245]
+ itasegm[246] itasegm[247] itasegm[248] itasegm[249] itasegm[24] itasegm[250] itasegm[251]
+ itasegm[252] itasegm[253] itasegm[254] itasegm[255] itasegm[256] itasegm[257] itasegm[258]
+ itasegm[259] itasegm[25] itasegm[260] itasegm[261] itasegm[262] itasegm[263] itasegm[264]
+ itasegm[265] itasegm[266] itasegm[267] itasegm[268] itasegm[269] itasegm[26] itasegm[270]
+ itasegm[271] itasegm[272] itasegm[273] itasegm[274] itasegm[275] itasegm[276] itasegm[277]
+ itasegm[278] itasegm[279] itasegm[27] itasegm[280] itasegm[281] itasegm[282] itasegm[283]
+ itasegm[284] itasegm[285] itasegm[286] itasegm[287] itasegm[288] itasegm[289] itasegm[28]
+ itasegm[290] itasegm[291] itasegm[292] itasegm[293] itasegm[294] itasegm[295] itasegm[296]
+ itasegm[297] itasegm[298] itasegm[299] itasegm[29] itasegm[2] itasegm[300] itasegm[301]
+ itasegm[302] itasegm[303] itasegm[304] itasegm[305] itasegm[306] itasegm[307] itasegm[308]
+ itasegm[309] itasegm[30] itasegm[310] itasegm[311] itasegm[312] itasegm[313] itasegm[314]
+ itasegm[315] itasegm[316] itasegm[317] itasegm[318] itasegm[319] itasegm[31] itasegm[320]
+ itasegm[321] itasegm[322] itasegm[323] itasegm[324] itasegm[325] itasegm[326] itasegm[327]
+ itasegm[328] itasegm[329] itasegm[32] itasegm[330] itasegm[331] itasegm[332] itasegm[333]
+ itasegm[334] itasegm[335] itasegm[336] itasegm[337] itasegm[338] itasegm[339] itasegm[33]
+ itasegm[340] itasegm[341] itasegm[342] itasegm[343] itasegm[344] itasegm[345] itasegm[346]
+ itasegm[347] itasegm[348] itasegm[349] itasegm[34] itasegm[350] itasegm[351] itasegm[352]
+ itasegm[353] itasegm[354] itasegm[355] itasegm[356] itasegm[357] itasegm[358] itasegm[359]
+ itasegm[35] itasegm[360] itasegm[361] itasegm[362] itasegm[363] itasegm[364] itasegm[365]
+ itasegm[366] itasegm[367] itasegm[368] itasegm[369] itasegm[36] itasegm[370] itasegm[371]
+ itasegm[372] itasegm[373] itasegm[374] itasegm[375] itasegm[376] itasegm[377] itasegm[378]
+ itasegm[379] itasegm[37] itasegm[380] itasegm[381] itasegm[382] itasegm[383] itasegm[384]
+ itasegm[385] itasegm[386] itasegm[387] itasegm[388] itasegm[389] itasegm[38] itasegm[390]
+ itasegm[391] itasegm[392] itasegm[393] itasegm[394] itasegm[395] itasegm[396] itasegm[397]
+ itasegm[398] itasegm[399] itasegm[39] itasegm[3] itasegm[400] itasegm[401] itasegm[402]
+ itasegm[403] itasegm[404] itasegm[405] itasegm[406] itasegm[407] itasegm[408] itasegm[409]
+ itasegm[40] itasegm[410] itasegm[411] itasegm[412] itasegm[413] itasegm[414] itasegm[415]
+ itasegm[416] itasegm[417] itasegm[418] itasegm[419] itasegm[41] itasegm[420] itasegm[421]
+ itasegm[422] itasegm[423] itasegm[424] itasegm[425] itasegm[426] itasegm[427] itasegm[428]
+ itasegm[429] itasegm[42] itasegm[430] itasegm[431] itasegm[432] itasegm[433] itasegm[434]
+ itasegm[435] itasegm[436] itasegm[437] itasegm[438] itasegm[439] itasegm[43] itasegm[440]
+ itasegm[441] itasegm[442] itasegm[443] itasegm[444] itasegm[445] itasegm[446] itasegm[447]
+ itasegm[448] itasegm[449] itasegm[44] itasegm[450] itasegm[451] itasegm[452] itasegm[453]
+ itasegm[454] itasegm[455] itasegm[456] itasegm[457] itasegm[458] itasegm[459] itasegm[45]
+ itasegm[460] itasegm[461] itasegm[462] itasegm[463] itasegm[464] itasegm[465] itasegm[466]
+ itasegm[467] itasegm[468] itasegm[469] itasegm[46] itasegm[470] itasegm[471] itasegm[472]
+ itasegm[473] itasegm[474] itasegm[475] itasegm[476] itasegm[477] itasegm[478] itasegm[479]
+ itasegm[47] itasegm[480] itasegm[481] itasegm[482] itasegm[483] itasegm[484] itasegm[485]
+ itasegm[486] itasegm[487] itasegm[488] itasegm[489] itasegm[48] itasegm[490] itasegm[491]
+ itasegm[492] itasegm[493] itasegm[494] itasegm[495] itasegm[496] itasegm[497] itasegm[498]
+ itasegm[499] itasegm[49] itasegm[4] itasegm[500] itasegm[501] itasegm[502] itasegm[503]
+ itasegm[504] itasegm[505] itasegm[506] itasegm[507] itasegm[508] itasegm[509] itasegm[50]
+ itasegm[510] itasegm[511] itasegm[512] itasegm[513] itasegm[514] itasegm[515] itasegm[516]
+ itasegm[517] itasegm[518] itasegm[519] itasegm[51] itasegm[520] itasegm[521] itasegm[522]
+ itasegm[523] itasegm[524] itasegm[525] itasegm[526] itasegm[527] itasegm[528] itasegm[529]
+ itasegm[52] itasegm[530] itasegm[531] itasegm[532] itasegm[533] itasegm[534] itasegm[535]
+ itasegm[536] itasegm[537] itasegm[538] itasegm[539] itasegm[53] itasegm[540] itasegm[541]
+ itasegm[542] itasegm[543] itasegm[544] itasegm[545] itasegm[546] itasegm[547] itasegm[548]
+ itasegm[549] itasegm[54] itasegm[550] itasegm[551] itasegm[552] itasegm[553] itasegm[554]
+ itasegm[555] itasegm[556] itasegm[557] itasegm[558] itasegm[559] itasegm[55] itasegm[560]
+ itasegm[561] itasegm[562] itasegm[563] itasegm[564] itasegm[565] itasegm[566] itasegm[567]
+ itasegm[568] itasegm[569] itasegm[56] itasegm[570] itasegm[571] itasegm[572] itasegm[573]
+ itasegm[574] itasegm[575] itasegm[576] itasegm[577] itasegm[578] itasegm[579] itasegm[57]
+ itasegm[580] itasegm[581] itasegm[582] itasegm[583] itasegm[584] itasegm[585] itasegm[586]
+ itasegm[587] itasegm[588] itasegm[589] itasegm[58] itasegm[590] itasegm[591] itasegm[592]
+ itasegm[593] itasegm[594] itasegm[595] itasegm[596] itasegm[597] itasegm[598] itasegm[599]
+ itasegm[59] itasegm[5] itasegm[600] itasegm[601] itasegm[602] itasegm[603] itasegm[604]
+ itasegm[605] itasegm[606] itasegm[607] itasegm[608] itasegm[609] itasegm[60] itasegm[610]
+ itasegm[611] itasegm[612] itasegm[613] itasegm[614] itasegm[615] itasegm[616] itasegm[617]
+ itasegm[618] itasegm[619] itasegm[61] itasegm[620] itasegm[621] itasegm[622] itasegm[623]
+ itasegm[624] itasegm[625] itasegm[626] itasegm[627] itasegm[628] itasegm[629] itasegm[62]
+ itasegm[630] itasegm[631] itasegm[632] itasegm[633] itasegm[634] itasegm[635] itasegm[636]
+ itasegm[637] itasegm[638] itasegm[639] itasegm[63] itasegm[640] itasegm[641] itasegm[642]
+ itasegm[643] itasegm[644] itasegm[645] itasegm[646] itasegm[647] itasegm[648] itasegm[649]
+ itasegm[64] itasegm[650] itasegm[651] itasegm[652] itasegm[653] itasegm[654] itasegm[655]
+ itasegm[656] itasegm[657] itasegm[658] itasegm[659] itasegm[65] itasegm[660] itasegm[661]
+ itasegm[662] itasegm[663] itasegm[664] itasegm[665] itasegm[666] itasegm[667] itasegm[668]
+ itasegm[669] itasegm[66] itasegm[670] itasegm[671] itasegm[672] itasegm[673] itasegm[674]
+ itasegm[675] itasegm[676] itasegm[677] itasegm[678] itasegm[679] itasegm[67] itasegm[680]
+ itasegm[681] itasegm[682] itasegm[683] itasegm[684] itasegm[685] itasegm[686] itasegm[687]
+ itasegm[688] itasegm[689] itasegm[68] itasegm[690] itasegm[691] itasegm[692] itasegm[693]
+ itasegm[694] itasegm[695] itasegm[696] itasegm[697] itasegm[698] itasegm[699] itasegm[69]
+ itasegm[6] itasegm[700] itasegm[701] itasegm[702] itasegm[703] itasegm[704] itasegm[705]
+ itasegm[706] itasegm[707] itasegm[708] itasegm[709] itasegm[70] itasegm[710] itasegm[711]
+ itasegm[712] itasegm[713] itasegm[714] itasegm[715] itasegm[716] itasegm[717] itasegm[718]
+ itasegm[719] itasegm[71] itasegm[720] itasegm[721] itasegm[722] itasegm[723] itasegm[724]
+ itasegm[725] itasegm[726] itasegm[727] itasegm[728] itasegm[729] itasegm[72] itasegm[730]
+ itasegm[731] itasegm[732] itasegm[733] itasegm[734] itasegm[735] itasegm[736] itasegm[737]
+ itasegm[738] itasegm[739] itasegm[73] itasegm[740] itasegm[741] itasegm[742] itasegm[743]
+ itasegm[744] itasegm[745] itasegm[746] itasegm[747] itasegm[748] itasegm[749] itasegm[74]
+ itasegm[750] itasegm[751] itasegm[752] itasegm[753] itasegm[754] itasegm[755] itasegm[756]
+ itasegm[757] itasegm[758] itasegm[759] itasegm[75] itasegm[760] itasegm[761] itasegm[762]
+ itasegm[763] itasegm[764] itasegm[765] itasegm[766] itasegm[767] itasegm[768] itasegm[769]
+ itasegm[76] itasegm[770] itasegm[771] itasegm[772] itasegm[773] itasegm[774] itasegm[775]
+ itasegm[776] itasegm[777] itasegm[778] itasegm[779] itasegm[77] itasegm[780] itasegm[781]
+ itasegm[782] itasegm[783] itasegm[784] itasegm[785] itasegm[786] itasegm[787] itasegm[788]
+ itasegm[789] itasegm[78] itasegm[790] itasegm[791] itasegm[792] itasegm[793] itasegm[794]
+ itasegm[795] itasegm[796] itasegm[797] itasegm[798] itasegm[799] itasegm[79] itasegm[7]
+ itasegm[800] itasegm[801] itasegm[802] itasegm[803] itasegm[804] itasegm[805] itasegm[806]
+ itasegm[807] itasegm[808] itasegm[809] itasegm[80] itasegm[810] itasegm[811] itasegm[812]
+ itasegm[813] itasegm[814] itasegm[815] itasegm[816] itasegm[817] itasegm[818] itasegm[819]
+ itasegm[81] itasegm[820] itasegm[821] itasegm[822] itasegm[823] itasegm[824] itasegm[825]
+ itasegm[826] itasegm[827] itasegm[828] itasegm[829] itasegm[82] itasegm[830] itasegm[831]
+ itasegm[832] itasegm[833] itasegm[834] itasegm[835] itasegm[836] itasegm[837] itasegm[838]
+ itasegm[839] itasegm[83] itasegm[840] itasegm[841] itasegm[842] itasegm[843] itasegm[844]
+ itasegm[845] itasegm[846] itasegm[847] itasegm[848] itasegm[849] itasegm[84] itasegm[850]
+ itasegm[851] itasegm[852] itasegm[853] itasegm[854] itasegm[855] itasegm[856] itasegm[857]
+ itasegm[858] itasegm[859] itasegm[85] itasegm[860] itasegm[861] itasegm[862] itasegm[863]
+ itasegm[864] itasegm[865] itasegm[866] itasegm[867] itasegm[868] itasegm[869] itasegm[86]
+ itasegm[870] itasegm[871] itasegm[872] itasegm[873] itasegm[874] itasegm[875] itasegm[876]
+ itasegm[877] itasegm[878] itasegm[879] itasegm[87] itasegm[880] itasegm[881] itasegm[882]
+ itasegm[883] itasegm[884] itasegm[885] itasegm[886] itasegm[887] itasegm[888] itasegm[889]
+ itasegm[88] itasegm[890] itasegm[891] itasegm[892] itasegm[893] itasegm[894] itasegm[895]
+ itasegm[89] itasegm[8] itasegm[90] itasegm[91] itasegm[92] itasegm[93] itasegm[94]
+ itasegm[95] itasegm[96] itasegm[97] itasegm[98] itasegm[99] itasegm[9] itasel[0]
+ itasel[100] itasel[101] itasel[102] itasel[103] itasel[104] itasel[105] itasel[106]
+ itasel[107] itasel[108] itasel[109] itasel[10] itasel[110] itasel[111] itasel[112]
+ itasel[113] itasel[114] itasel[115] itasel[116] itasel[117] itasel[118] itasel[119]
+ itasel[11] itasel[120] itasel[121] itasel[122] itasel[123] itasel[124] itasel[125]
+ itasel[126] itasel[127] itasel[128] itasel[129] itasel[12] itasel[130] itasel[131]
+ itasel[132] itasel[133] itasel[134] itasel[135] itasel[136] itasel[137] itasel[138]
+ itasel[139] itasel[13] itasel[140] itasel[141] itasel[142] itasel[143] itasel[144]
+ itasel[145] itasel[146] itasel[147] itasel[148] itasel[149] itasel[14] itasel[150]
+ itasel[151] itasel[152] itasel[153] itasel[154] itasel[155] itasel[156] itasel[157]
+ itasel[158] itasel[159] itasel[15] itasel[160] itasel[161] itasel[162] itasel[163]
+ itasel[164] itasel[165] itasel[166] itasel[167] itasel[168] itasel[169] itasel[16]
+ itasel[170] itasel[171] itasel[172] itasel[173] itasel[174] itasel[175] itasel[176]
+ itasel[177] itasel[178] itasel[179] itasel[17] itasel[180] itasel[181] itasel[182]
+ itasel[183] itasel[184] itasel[185] itasel[186] itasel[187] itasel[188] itasel[189]
+ itasel[18] itasel[190] itasel[191] itasel[192] itasel[193] itasel[194] itasel[195]
+ itasel[196] itasel[197] itasel[198] itasel[199] itasel[19] itasel[1] itasel[200]
+ itasel[201] itasel[202] itasel[203] itasel[204] itasel[205] itasel[206] itasel[207]
+ itasel[208] itasel[209] itasel[20] itasel[210] itasel[211] itasel[212] itasel[213]
+ itasel[214] itasel[215] itasel[216] itasel[217] itasel[218] itasel[219] itasel[21]
+ itasel[220] itasel[221] itasel[222] itasel[223] itasel[224] itasel[225] itasel[226]
+ itasel[227] itasel[228] itasel[229] itasel[22] itasel[230] itasel[231] itasel[232]
+ itasel[233] itasel[234] itasel[235] itasel[236] itasel[237] itasel[238] itasel[239]
+ itasel[23] itasel[240] itasel[241] itasel[242] itasel[243] itasel[244] itasel[245]
+ itasel[246] itasel[247] itasel[248] itasel[249] itasel[24] itasel[250] itasel[251]
+ itasel[252] itasel[253] itasel[254] itasel[255] itasel[256] itasel[257] itasel[258]
+ itasel[259] itasel[25] itasel[260] itasel[261] itasel[262] itasel[263] itasel[264]
+ itasel[265] itasel[266] itasel[267] itasel[268] itasel[269] itasel[26] itasel[270]
+ itasel[271] itasel[272] itasel[273] itasel[274] itasel[275] itasel[276] itasel[277]
+ itasel[278] itasel[279] itasel[27] itasel[280] itasel[281] itasel[282] itasel[283]
+ itasel[284] itasel[285] itasel[286] itasel[287] itasel[288] itasel[289] itasel[28]
+ itasel[290] itasel[291] itasel[292] itasel[293] itasel[294] itasel[295] itasel[296]
+ itasel[297] itasel[298] itasel[299] itasel[29] itasel[2] itasel[300] itasel[301]
+ itasel[302] itasel[303] itasel[304] itasel[305] itasel[306] itasel[307] itasel[308]
+ itasel[309] itasel[30] itasel[310] itasel[311] itasel[312] itasel[313] itasel[314]
+ itasel[315] itasel[316] itasel[317] itasel[318] itasel[319] itasel[31] itasel[320]
+ itasel[321] itasel[322] itasel[323] itasel[324] itasel[325] itasel[326] itasel[327]
+ itasel[328] itasel[329] itasel[32] itasel[330] itasel[331] itasel[332] itasel[333]
+ itasel[334] itasel[335] itasel[336] itasel[337] itasel[338] itasel[339] itasel[33]
+ itasel[340] itasel[341] itasel[342] itasel[343] itasel[344] itasel[345] itasel[346]
+ itasel[347] itasel[348] itasel[349] itasel[34] itasel[350] itasel[351] itasel[352]
+ itasel[353] itasel[354] itasel[355] itasel[356] itasel[357] itasel[358] itasel[359]
+ itasel[35] itasel[360] itasel[361] itasel[362] itasel[363] itasel[364] itasel[365]
+ itasel[366] itasel[367] itasel[368] itasel[369] itasel[36] itasel[370] itasel[371]
+ itasel[372] itasel[373] itasel[374] itasel[375] itasel[376] itasel[377] itasel[378]
+ itasel[379] itasel[37] itasel[380] itasel[381] itasel[382] itasel[383] itasel[384]
+ itasel[385] itasel[386] itasel[387] itasel[388] itasel[389] itasel[38] itasel[390]
+ itasel[391] itasel[392] itasel[393] itasel[394] itasel[395] itasel[396] itasel[397]
+ itasel[398] itasel[399] itasel[39] itasel[3] itasel[400] itasel[401] itasel[402]
+ itasel[403] itasel[404] itasel[405] itasel[406] itasel[407] itasel[408] itasel[409]
+ itasel[40] itasel[410] itasel[411] itasel[412] itasel[413] itasel[414] itasel[415]
+ itasel[416] itasel[417] itasel[418] itasel[419] itasel[41] itasel[420] itasel[421]
+ itasel[422] itasel[423] itasel[424] itasel[425] itasel[426] itasel[427] itasel[428]
+ itasel[429] itasel[42] itasel[430] itasel[431] itasel[432] itasel[433] itasel[434]
+ itasel[435] itasel[436] itasel[437] itasel[438] itasel[439] itasel[43] itasel[440]
+ itasel[441] itasel[442] itasel[443] itasel[444] itasel[445] itasel[446] itasel[447]
+ itasel[448] itasel[449] itasel[44] itasel[450] itasel[451] itasel[452] itasel[453]
+ itasel[454] itasel[455] itasel[456] itasel[457] itasel[458] itasel[459] itasel[45]
+ itasel[460] itasel[461] itasel[462] itasel[463] itasel[464] itasel[465] itasel[466]
+ itasel[467] itasel[468] itasel[469] itasel[46] itasel[470] itasel[471] itasel[472]
+ itasel[473] itasel[474] itasel[475] itasel[476] itasel[477] itasel[478] itasel[479]
+ itasel[47] itasel[480] itasel[481] itasel[482] itasel[483] itasel[484] itasel[485]
+ itasel[486] itasel[487] itasel[488] itasel[489] itasel[48] itasel[490] itasel[491]
+ itasel[492] itasel[493] itasel[494] itasel[495] itasel[496] itasel[497] itasel[498]
+ itasel[499] itasel[49] itasel[4] itasel[500] itasel[501] itasel[502] itasel[503]
+ itasel[504] itasel[505] itasel[506] itasel[507] itasel[508] itasel[509] itasel[50]
+ itasel[510] itasel[511] itasel[512] itasel[513] itasel[514] itasel[515] itasel[516]
+ itasel[517] itasel[518] itasel[519] itasel[51] itasel[520] itasel[521] itasel[522]
+ itasel[523] itasel[524] itasel[525] itasel[526] itasel[527] itasel[528] itasel[529]
+ itasel[52] itasel[530] itasel[531] itasel[532] itasel[533] itasel[534] itasel[535]
+ itasel[536] itasel[537] itasel[538] itasel[539] itasel[53] itasel[540] itasel[541]
+ itasel[542] itasel[543] itasel[544] itasel[545] itasel[546] itasel[547] itasel[548]
+ itasel[549] itasel[54] itasel[550] itasel[551] itasel[552] itasel[553] itasel[554]
+ itasel[555] itasel[556] itasel[557] itasel[558] itasel[559] itasel[55] itasel[560]
+ itasel[561] itasel[562] itasel[563] itasel[564] itasel[565] itasel[566] itasel[567]
+ itasel[568] itasel[569] itasel[56] itasel[570] itasel[571] itasel[572] itasel[573]
+ itasel[574] itasel[575] itasel[576] itasel[577] itasel[578] itasel[579] itasel[57]
+ itasel[580] itasel[581] itasel[582] itasel[583] itasel[584] itasel[585] itasel[586]
+ itasel[587] itasel[588] itasel[589] itasel[58] itasel[590] itasel[591] itasel[592]
+ itasel[593] itasel[594] itasel[595] itasel[596] itasel[597] itasel[598] itasel[599]
+ itasel[59] itasel[5] itasel[600] itasel[601] itasel[602] itasel[603] itasel[604]
+ itasel[605] itasel[606] itasel[607] itasel[608] itasel[609] itasel[60] itasel[610]
+ itasel[611] itasel[612] itasel[613] itasel[614] itasel[615] itasel[616] itasel[617]
+ itasel[618] itasel[619] itasel[61] itasel[620] itasel[621] itasel[622] itasel[623]
+ itasel[624] itasel[625] itasel[626] itasel[627] itasel[628] itasel[629] itasel[62]
+ itasel[630] itasel[631] itasel[632] itasel[633] itasel[634] itasel[635] itasel[636]
+ itasel[637] itasel[638] itasel[639] itasel[63] itasel[640] itasel[641] itasel[642]
+ itasel[643] itasel[644] itasel[645] itasel[646] itasel[647] itasel[648] itasel[649]
+ itasel[64] itasel[650] itasel[651] itasel[652] itasel[653] itasel[654] itasel[655]
+ itasel[656] itasel[657] itasel[658] itasel[659] itasel[65] itasel[660] itasel[661]
+ itasel[662] itasel[663] itasel[664] itasel[665] itasel[666] itasel[667] itasel[668]
+ itasel[669] itasel[66] itasel[670] itasel[671] itasel[672] itasel[673] itasel[674]
+ itasel[675] itasel[676] itasel[677] itasel[678] itasel[679] itasel[67] itasel[680]
+ itasel[681] itasel[682] itasel[683] itasel[684] itasel[685] itasel[686] itasel[687]
+ itasel[688] itasel[689] itasel[68] itasel[690] itasel[691] itasel[692] itasel[693]
+ itasel[694] itasel[695] itasel[696] itasel[697] itasel[698] itasel[699] itasel[69]
+ itasel[6] itasel[700] itasel[701] itasel[702] itasel[703] itasel[704] itasel[705]
+ itasel[706] itasel[707] itasel[708] itasel[709] itasel[70] itasel[710] itasel[711]
+ itasel[712] itasel[713] itasel[714] itasel[715] itasel[716] itasel[717] itasel[718]
+ itasel[719] itasel[71] itasel[720] itasel[721] itasel[722] itasel[723] itasel[724]
+ itasel[725] itasel[726] itasel[727] itasel[728] itasel[729] itasel[72] itasel[730]
+ itasel[731] itasel[732] itasel[733] itasel[734] itasel[735] itasel[736] itasel[737]
+ itasel[738] itasel[739] itasel[73] itasel[740] itasel[741] itasel[742] itasel[743]
+ itasel[744] itasel[745] itasel[746] itasel[747] itasel[748] itasel[749] itasel[74]
+ itasel[750] itasel[751] itasel[752] itasel[753] itasel[754] itasel[755] itasel[756]
+ itasel[757] itasel[758] itasel[759] itasel[75] itasel[760] itasel[761] itasel[762]
+ itasel[763] itasel[764] itasel[765] itasel[766] itasel[767] itasel[76] itasel[77]
+ itasel[78] itasel[79] itasel[7] itasel[80] itasel[81] itasel[82] itasel[83] itasel[84]
+ itasel[85] itasel[86] itasel[87] itasel[88] itasel[89] itasel[8] itasel[90] itasel[91]
+ itasel[92] itasel[93] itasel[94] itasel[95] itasel[96] itasel[97] itasel[98] itasel[99]
+ itasel[9] nsel[0] nsel[1] nsel[2] nsel[3] nsel[4] nsel[5] segm[0] segm[10] segm[11]
+ segm[12] segm[13] segm[1] segm[2] segm[3] segm[4] segm[5] segm[6] segm[7] segm[8]
+ segm[9] sel[0] sel[10] sel[11] sel[1] sel[2] sel[3] sel[4] sel[5] sel[6] sel[7]
+ sel[8] sel[9] vdd vss
.ends

* Black-box entry subcircuit for ita20 abstract view
.subckt ita20 clk segm[0] segm[10] segm[11] segm[12] segm[13] segm[1] segm[2] segm[3]
+ segm[4] segm[5] segm[6] segm[7] segm[8] segm[9] sel[0] sel[10] sel[11] sel[1] sel[2]
+ sel[3] sel[4] sel[5] sel[6] sel[7] sel[8] sel[9] vdd vss
.ends

* Black-box entry subcircuit for ita42 abstract view
.subckt ita42 clk segm[0] segm[10] segm[11] segm[12] segm[13] segm[1] segm[2] segm[3]
+ segm[4] segm[5] segm[6] segm[7] segm[8] segm[9] sel[0] sel[10] sel[11] sel[1] sel[2]
+ sel[3] sel[4] sel[5] sel[6] sel[7] sel[8] sel[9] vdd vss
.ends

* Black-box entry subcircuit for ita32 abstract view
.subckt ita32 clk segm[0] segm[10] segm[11] segm[12] segm[13] segm[1] segm[2] segm[3]
+ segm[4] segm[5] segm[6] segm[7] segm[8] segm[9] sel[0] sel[10] sel[11] sel[1] sel[2]
+ sel[3] sel[4] sel[5] sel[6] sel[7] sel[8] sel[9] vdd vss
.ends

* Black-box entry subcircuit for ita7 abstract view
.subckt ita7 clk segm[0] segm[10] segm[11] segm[12] segm[13] segm[1] segm[2] segm[3]
+ segm[4] segm[5] segm[6] segm[7] segm[8] segm[9] sel[0] sel[10] sel[11] sel[1] sel[2]
+ sel[3] sel[4] sel[5] sel[6] sel[7] sel[8] sel[9] vdd vss
.ends

* Black-box entry subcircuit for ita54 abstract view
.subckt ita54 clk segm[0] segm[10] segm[11] segm[12] segm[13] segm[1] segm[2] segm[3]
+ segm[4] segm[5] segm[6] segm[7] segm[8] segm[9] sel[0] sel[10] sel[11] sel[1] sel[2]
+ sel[3] sel[4] sel[5] sel[6] sel[7] sel[8] sel[9] vdd vss
.ends

* Black-box entry subcircuit for ita21 abstract view
.subckt ita21 clk segm[0] segm[10] segm[11] segm[12] segm[13] segm[1] segm[2] segm[3]
+ segm[4] segm[5] segm[6] segm[7] segm[8] segm[9] sel[0] sel[10] sel[11] sel[1] sel[2]
+ sel[3] sel[4] sel[5] sel[6] sel[7] sel[8] sel[9] vdd vss
.ends

* Black-box entry subcircuit for ita43 abstract view
.subckt ita43 clk segm[0] segm[10] segm[11] segm[12] segm[13] segm[1] segm[2] segm[3]
+ segm[4] segm[5] segm[6] segm[7] segm[8] segm[9] sel[0] sel[10] sel[11] sel[1] sel[2]
+ sel[3] sel[4] sel[5] sel[6] sel[7] sel[8] sel[9] vdd vss
.ends

* Black-box entry subcircuit for ita10 abstract view
.subckt ita10 clk segm[0] segm[10] segm[11] segm[12] segm[13] segm[1] segm[2] segm[3]
+ segm[4] segm[5] segm[6] segm[7] segm[8] segm[9] sel[0] sel[10] sel[11] sel[1] sel[2]
+ sel[3] sel[4] sel[5] sel[6] sel[7] sel[8] sel[9] vdd vss
.ends

* Black-box entry subcircuit for ita8 abstract view
.subckt ita8 clk segm[0] segm[10] segm[11] segm[12] segm[13] segm[1] segm[2] segm[3]
+ segm[4] segm[5] segm[6] segm[7] segm[8] segm[9] sel[0] sel[10] sel[11] sel[1] sel[2]
+ sel[3] sel[4] sel[5] sel[6] sel[7] sel[8] sel[9] vdd vss
.ends

* Black-box entry subcircuit for ita55 abstract view
.subckt ita55 clk segm[0] segm[10] segm[11] segm[12] segm[13] segm[1] segm[2] segm[3]
+ segm[4] segm[5] segm[6] segm[7] segm[8] segm[9] sel[0] sel[10] sel[11] sel[1] sel[2]
+ sel[3] sel[4] sel[5] sel[6] sel[7] sel[8] sel[9] vdd vss
.ends

* Black-box entry subcircuit for ita22 abstract view
.subckt ita22 clk segm[0] segm[10] segm[11] segm[12] segm[13] segm[1] segm[2] segm[3]
+ segm[4] segm[5] segm[6] segm[7] segm[8] segm[9] sel[0] sel[10] sel[11] sel[1] sel[2]
+ sel[3] sel[4] sel[5] sel[6] sel[7] sel[8] sel[9] vdd vss
.ends

* Black-box entry subcircuit for ita44 abstract view
.subckt ita44 clk segm[0] segm[10] segm[11] segm[12] segm[13] segm[1] segm[2] segm[3]
+ segm[4] segm[5] segm[6] segm[7] segm[8] segm[9] sel[0] sel[10] sel[11] sel[1] sel[2]
+ sel[3] sel[4] sel[5] sel[6] sel[7] sel[8] sel[9] vdd vss
.ends

* Black-box entry subcircuit for ita11 abstract view
.subckt ita11 clk segm[0] segm[10] segm[11] segm[12] segm[13] segm[1] segm[2] segm[3]
+ segm[4] segm[5] segm[6] segm[7] segm[8] segm[9] sel[0] sel[10] sel[11] sel[1] sel[2]
+ sel[3] sel[4] sel[5] sel[6] sel[7] sel[8] sel[9] vdd vss
.ends

* Black-box entry subcircuit for ita33 abstract view
.subckt ita33 clk segm[0] segm[10] segm[11] segm[12] segm[13] segm[1] segm[2] segm[3]
+ segm[4] segm[5] segm[6] segm[7] segm[8] segm[9] sel[0] sel[10] sel[11] sel[1] sel[2]
+ sel[3] sel[4] sel[5] sel[6] sel[7] sel[8] sel[9] vdd vss
.ends

* Black-box entry subcircuit for ita56 abstract view
.subckt ita56 clk segm[0] segm[10] segm[11] segm[12] segm[13] segm[1] segm[2] segm[3]
+ segm[4] segm[5] segm[6] segm[7] segm[8] segm[9] sel[0] sel[10] sel[11] sel[1] sel[2]
+ sel[3] sel[4] sel[5] sel[6] sel[7] sel[8] sel[9] vdd vss
.ends

* Black-box entry subcircuit for ita23 abstract view
.subckt ita23 clk segm[0] segm[10] segm[11] segm[12] segm[13] segm[1] segm[2] segm[3]
+ segm[4] segm[5] segm[6] segm[7] segm[8] segm[9] sel[0] sel[10] sel[11] sel[1] sel[2]
+ sel[3] sel[4] sel[5] sel[6] sel[7] sel[8] sel[9] vdd vss
.ends

* Black-box entry subcircuit for ita45 abstract view
.subckt ita45 clk segm[0] segm[10] segm[11] segm[12] segm[13] segm[1] segm[2] segm[3]
+ segm[4] segm[5] segm[6] segm[7] segm[8] segm[9] sel[0] sel[10] sel[11] sel[1] sel[2]
+ sel[3] sel[4] sel[5] sel[6] sel[7] sel[8] sel[9] vdd vss
.ends

* Black-box entry subcircuit for ita12 abstract view
.subckt ita12 clk segm[0] segm[10] segm[11] segm[12] segm[13] segm[1] segm[2] segm[3]
+ segm[4] segm[5] segm[6] segm[7] segm[8] segm[9] sel[0] sel[10] sel[11] sel[1] sel[2]
+ sel[3] sel[4] sel[5] sel[6] sel[7] sel[8] sel[9] vdd vss
.ends

* Black-box entry subcircuit for ita34 abstract view
.subckt ita34 clk segm[0] segm[10] segm[11] segm[12] segm[13] segm[1] segm[2] segm[3]
+ segm[4] segm[5] segm[6] segm[7] segm[8] segm[9] sel[0] sel[10] sel[11] sel[1] sel[2]
+ sel[3] sel[4] sel[5] sel[6] sel[7] sel[8] sel[9] vdd vss
.ends

* Black-box entry subcircuit for ita9 abstract view
.subckt ita9 clk segm[0] segm[10] segm[11] segm[12] segm[13] segm[1] segm[2] segm[3]
+ segm[4] segm[5] segm[6] segm[7] segm[8] segm[9] sel[0] sel[10] sel[11] sel[1] sel[2]
+ sel[3] sel[4] sel[5] sel[6] sel[7] sel[8] sel[9] vdd vss
.ends

* Black-box entry subcircuit for ita24 abstract view
.subckt ita24 clk segm[0] segm[10] segm[11] segm[12] segm[13] segm[1] segm[2] segm[3]
+ segm[4] segm[5] segm[6] segm[7] segm[8] segm[9] sel[0] sel[10] sel[11] sel[1] sel[2]
+ sel[3] sel[4] sel[5] sel[6] sel[7] sel[8] sel[9] vdd vss
.ends

* Black-box entry subcircuit for ita47 abstract view
.subckt ita47 clk segm[0] segm[10] segm[11] segm[12] segm[13] segm[1] segm[2] segm[3]
+ segm[4] segm[5] segm[6] segm[7] segm[8] segm[9] sel[0] sel[10] sel[11] sel[1] sel[2]
+ sel[3] sel[4] sel[5] sel[6] sel[7] sel[8] sel[9] vdd vss
.ends

* Black-box entry subcircuit for ita46 abstract view
.subckt ita46 clk segm[0] segm[10] segm[11] segm[12] segm[13] segm[1] segm[2] segm[3]
+ segm[4] segm[5] segm[6] segm[7] segm[8] segm[9] sel[0] sel[10] sel[11] sel[1] sel[2]
+ sel[3] sel[4] sel[5] sel[6] sel[7] sel[8] sel[9] vdd vss
.ends

* Black-box entry subcircuit for ita14 abstract view
.subckt ita14 clk segm[0] segm[10] segm[11] segm[12] segm[13] segm[1] segm[2] segm[3]
+ segm[4] segm[5] segm[6] segm[7] segm[8] segm[9] sel[0] sel[10] sel[11] sel[1] sel[2]
+ sel[3] sel[4] sel[5] sel[6] sel[7] sel[8] sel[9] vdd vss
.ends

* Black-box entry subcircuit for ita13 abstract view
.subckt ita13 clk segm[0] segm[10] segm[11] segm[12] segm[13] segm[1] segm[2] segm[3]
+ segm[4] segm[5] segm[6] segm[7] segm[8] segm[9] sel[0] sel[10] sel[11] sel[1] sel[2]
+ sel[3] sel[4] sel[5] sel[6] sel[7] sel[8] sel[9] vdd vss
.ends

* Black-box entry subcircuit for ita36 abstract view
.subckt ita36 clk segm[0] segm[10] segm[11] segm[12] segm[13] segm[1] segm[2] segm[3]
+ segm[4] segm[5] segm[6] segm[7] segm[8] segm[9] sel[0] sel[10] sel[11] sel[1] sel[2]
+ sel[3] sel[4] sel[5] sel[6] sel[7] sel[8] sel[9] vdd vss
.ends

* Black-box entry subcircuit for ita35 abstract view
.subckt ita35 clk segm[0] segm[10] segm[11] segm[12] segm[13] segm[1] segm[2] segm[3]
+ segm[4] segm[5] segm[6] segm[7] segm[8] segm[9] sel[0] sel[10] sel[11] sel[1] sel[2]
+ sel[3] sel[4] sel[5] sel[6] sel[7] sel[8] sel[9] vdd vss
.ends

* Black-box entry subcircuit for ita57 abstract view
.subckt ita57 clk segm[0] segm[10] segm[11] segm[12] segm[13] segm[1] segm[2] segm[3]
+ segm[4] segm[5] segm[6] segm[7] segm[8] segm[9] sel[0] sel[10] sel[11] sel[1] sel[2]
+ sel[3] sel[4] sel[5] sel[6] sel[7] sel[8] sel[9] vdd vss
.ends

* Black-box entry subcircuit for ita58 abstract view
.subckt ita58 clk segm[0] segm[10] segm[11] segm[12] segm[13] segm[1] segm[2] segm[3]
+ segm[4] segm[5] segm[6] segm[7] segm[8] segm[9] sel[0] sel[10] sel[11] sel[1] sel[2]
+ sel[3] sel[4] sel[5] sel[6] sel[7] sel[8] sel[9] vdd vss
.ends

* Black-box entry subcircuit for ita25 abstract view
.subckt ita25 clk segm[0] segm[10] segm[11] segm[12] segm[13] segm[1] segm[2] segm[3]
+ segm[4] segm[5] segm[6] segm[7] segm[8] segm[9] sel[0] sel[10] sel[11] sel[1] sel[2]
+ sel[3] sel[4] sel[5] sel[6] sel[7] sel[8] sel[9] vdd vss
.ends

* Black-box entry subcircuit for ita48 abstract view
.subckt ita48 clk segm[0] segm[10] segm[11] segm[12] segm[13] segm[1] segm[2] segm[3]
+ segm[4] segm[5] segm[6] segm[7] segm[8] segm[9] sel[0] sel[10] sel[11] sel[1] sel[2]
+ sel[3] sel[4] sel[5] sel[6] sel[7] sel[8] sel[9] vdd vss
.ends

* Black-box entry subcircuit for ita15 abstract view
.subckt ita15 clk segm[0] segm[10] segm[11] segm[12] segm[13] segm[1] segm[2] segm[3]
+ segm[4] segm[5] segm[6] segm[7] segm[8] segm[9] sel[0] sel[10] sel[11] sel[1] sel[2]
+ sel[3] sel[4] sel[5] sel[6] sel[7] sel[8] sel[9] vdd vss
.ends

* Black-box entry subcircuit for ita37 abstract view
.subckt ita37 clk segm[0] segm[10] segm[11] segm[12] segm[13] segm[1] segm[2] segm[3]
+ segm[4] segm[5] segm[6] segm[7] segm[8] segm[9] sel[0] sel[10] sel[11] sel[1] sel[2]
+ sel[3] sel[4] sel[5] sel[6] sel[7] sel[8] sel[9] vdd vss
.ends

* Black-box entry subcircuit for ita59 abstract view
.subckt ita59 clk segm[0] segm[10] segm[11] segm[12] segm[13] segm[1] segm[2] segm[3]
+ segm[4] segm[5] segm[6] segm[7] segm[8] segm[9] sel[0] sel[10] sel[11] sel[1] sel[2]
+ sel[3] sel[4] sel[5] sel[6] sel[7] sel[8] sel[9] vdd vss
.ends

* Black-box entry subcircuit for ita26 abstract view
.subckt ita26 clk segm[0] segm[10] segm[11] segm[12] segm[13] segm[1] segm[2] segm[3]
+ segm[4] segm[5] segm[6] segm[7] segm[8] segm[9] sel[0] sel[10] sel[11] sel[1] sel[2]
+ sel[3] sel[4] sel[5] sel[6] sel[7] sel[8] sel[9] vdd vss
.ends

* Black-box entry subcircuit for ita16 abstract view
.subckt ita16 clk segm[0] segm[10] segm[11] segm[12] segm[13] segm[1] segm[2] segm[3]
+ segm[4] segm[5] segm[6] segm[7] segm[8] segm[9] sel[0] sel[10] sel[11] sel[1] sel[2]
+ sel[3] sel[4] sel[5] sel[6] sel[7] sel[8] sel[9] vdd vss
.ends

* Black-box entry subcircuit for ita38 abstract view
.subckt ita38 clk segm[0] segm[10] segm[11] segm[12] segm[13] segm[1] segm[2] segm[3]
+ segm[4] segm[5] segm[6] segm[7] segm[8] segm[9] sel[0] sel[10] sel[11] sel[1] sel[2]
+ sel[3] sel[4] sel[5] sel[6] sel[7] sel[8] sel[9] vdd vss
.ends

* Black-box entry subcircuit for ita27 abstract view
.subckt ita27 clk segm[0] segm[10] segm[11] segm[12] segm[13] segm[1] segm[2] segm[3]
+ segm[4] segm[5] segm[6] segm[7] segm[8] segm[9] sel[0] sel[10] sel[11] sel[1] sel[2]
+ sel[3] sel[4] sel[5] sel[6] sel[7] sel[8] sel[9] vdd vss
.ends

* Black-box entry subcircuit for ita49 abstract view
.subckt ita49 clk segm[0] segm[10] segm[11] segm[12] segm[13] segm[1] segm[2] segm[3]
+ segm[4] segm[5] segm[6] segm[7] segm[8] segm[9] sel[0] sel[10] sel[11] sel[1] sel[2]
+ sel[3] sel[4] sel[5] sel[6] sel[7] sel[8] sel[9] vdd vss
.ends

* Black-box entry subcircuit for ita39 abstract view
.subckt ita39 clk segm[0] segm[10] segm[11] segm[12] segm[13] segm[1] segm[2] segm[3]
+ segm[4] segm[5] segm[6] segm[7] segm[8] segm[9] sel[0] sel[10] sel[11] sel[1] sel[2]
+ sel[3] sel[4] sel[5] sel[6] sel[7] sel[8] sel[9] vdd vss
.ends

* Black-box entry subcircuit for ita28 abstract view
.subckt ita28 clk segm[0] segm[10] segm[11] segm[12] segm[13] segm[1] segm[2] segm[3]
+ segm[4] segm[5] segm[6] segm[7] segm[8] segm[9] sel[0] sel[10] sel[11] sel[1] sel[2]
+ sel[3] sel[4] sel[5] sel[6] sel[7] sel[8] sel[9] vdd vss
.ends

* Black-box entry subcircuit for ita17 abstract view
.subckt ita17 clk segm[0] segm[10] segm[11] segm[12] segm[13] segm[1] segm[2] segm[3]
+ segm[4] segm[5] segm[6] segm[7] segm[8] segm[9] sel[0] sel[10] sel[11] sel[1] sel[2]
+ sel[3] sel[4] sel[5] sel[6] sel[7] sel[8] sel[9] vdd vss
.ends

* Black-box entry subcircuit for ita29 abstract view
.subckt ita29 clk segm[0] segm[10] segm[11] segm[12] segm[13] segm[1] segm[2] segm[3]
+ segm[4] segm[5] segm[6] segm[7] segm[8] segm[9] sel[0] sel[10] sel[11] sel[1] sel[2]
+ sel[3] sel[4] sel[5] sel[6] sel[7] sel[8] sel[9] vdd vss
.ends

* Black-box entry subcircuit for ita18 abstract view
.subckt ita18 clk segm[0] segm[10] segm[11] segm[12] segm[13] segm[1] segm[2] segm[3]
+ segm[4] segm[5] segm[6] segm[7] segm[8] segm[9] sel[0] sel[10] sel[11] sel[1] sel[2]
+ sel[3] sel[4] sel[5] sel[6] sel[7] sel[8] sel[9] vdd vss
.ends

* Black-box entry subcircuit for ita19 abstract view
.subckt ita19 clk segm[0] segm[10] segm[11] segm[12] segm[13] segm[1] segm[2] segm[3]
+ segm[4] segm[5] segm[6] segm[7] segm[8] segm[9] sel[0] sel[10] sel[11] sel[1] sel[2]
+ sel[3] sel[4] sel[5] sel[6] sel[7] sel[8] sel[9] vdd vss
.ends

.subckt user_project_wrapper io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14]
+ io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22]
+ io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30]
+ io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12]
+ io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1]
+ io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27]
+ io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34]
+ io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29]
+ io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36]
+ io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9]
+ la_data_in[0] la_data_in[10] la_data_in[11] la_data_in[12] la_data_in[13] la_data_in[14]
+ la_data_in[15] la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1]
+ la_data_in[20] la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25]
+ la_data_in[26] la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30]
+ la_data_in[31] la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36]
+ la_data_in[37] la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41]
+ la_data_in[42] la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47]
+ la_data_in[48] la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52]
+ la_data_in[53] la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58]
+ la_data_in[59] la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63]
+ la_data_in[6] la_data_in[7] la_data_in[8] la_data_in[9] la_data_out[0] la_data_out[10]
+ la_data_out[11] la_data_out[12] la_data_out[13] la_data_out[14] la_data_out[15]
+ la_data_out[16] la_data_out[17] la_data_out[18] la_data_out[19] la_data_out[1] la_data_out[20]
+ la_data_out[21] la_data_out[22] la_data_out[23] la_data_out[24] la_data_out[25]
+ la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29] la_data_out[2] la_data_out[30]
+ la_data_out[31] la_data_out[32] la_data_out[33] la_data_out[34] la_data_out[35]
+ la_data_out[36] la_data_out[37] la_data_out[38] la_data_out[39] la_data_out[3] la_data_out[40]
+ la_data_out[41] la_data_out[42] la_data_out[43] la_data_out[44] la_data_out[45]
+ la_data_out[46] la_data_out[47] la_data_out[48] la_data_out[49] la_data_out[4] la_data_out[50]
+ la_data_out[51] la_data_out[52] la_data_out[53] la_data_out[54] la_data_out[55]
+ la_data_out[56] la_data_out[57] la_data_out[58] la_data_out[59] la_data_out[5] la_data_out[60]
+ la_data_out[61] la_data_out[62] la_data_out[63] la_data_out[6] la_data_out[7] la_data_out[8]
+ la_data_out[9] la_oenb[0] la_oenb[10] la_oenb[11] la_oenb[12] la_oenb[13] la_oenb[14]
+ la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20]
+ la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27]
+ la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33]
+ la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[3]
+ la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46]
+ la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52]
+ la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59]
+ la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63] la_oenb[6] la_oenb[7]
+ la_oenb[8] la_oenb[9] user_clock2 user_irq[0] user_irq[1] user_irq[2] vdd vss wb_clk_i
+ wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13]
+ wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19]
+ wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24]
+ wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2]
+ wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6]
+ wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11]
+ wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17]
+ wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22]
+ wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28]
+ wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4]
+ wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10]
+ wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16]
+ wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21]
+ wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27]
+ wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3]
+ wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0]
+ wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
Xita60 wb_clk_i itasegm1\[826\] itasegm1\[836\] itasegm1\[837\] itasegm1\[838\] itasegm1\[839\]
+ itasegm1\[827\] itasegm1\[828\] itasegm1\[829\] itasegm1\[830\] itasegm1\[831\]
+ itasegm1\[832\] itasegm1\[833\] itasegm1\[834\] itasegm1\[835\] itasel1\[708\] itasel1\[718\]
+ itasel1\[719\] itasel1\[709\] itasel1\[710\] itasel1\[711\] itasel1\[712\] itasel1\[713\]
+ itasel1\[714\] itasel1\[715\] itasel1\[716\] itasel1\[717\] vdd vss ita60
Xita1 wb_clk_i itasegm1\[0\] itasegm1\[10\] itasegm1\[11\] itasegm1\[12\] itasegm1\[13\]
+ itasegm1\[1\] itasegm1\[2\] itasegm1\[3\] itasegm1\[4\] itasegm1\[5\] itasegm1\[6\]
+ itasegm1\[7\] itasegm1\[8\] itasegm1\[9\] itasel1\[0\] itasel1\[10\] itasel1\[11\]
+ itasel1\[1\] itasel1\[2\] itasel1\[3\] itasel1\[4\] itasel1\[5\] itasel1\[6\] itasel1\[7\]
+ itasel1\[8\] itasel1\[9\] vdd vss ita1
Xita61 wb_clk_i itasegm1\[840\] itasegm1\[850\] itasegm1\[851\] itasegm1\[852\] itasegm1\[853\]
+ itasegm1\[841\] itasegm1\[842\] itasegm1\[843\] itasegm1\[844\] itasegm1\[845\]
+ itasegm1\[846\] itasegm1\[847\] itasegm1\[848\] itasegm1\[849\] itasel1\[720\] itasel1\[730\]
+ itasel1\[731\] itasel1\[721\] itasel1\[722\] itasel1\[723\] itasel1\[724\] itasel1\[725\]
+ itasel1\[726\] itasel1\[727\] itasel1\[728\] itasel1\[729\] vdd vss ita61
Xita50 wb_clk_i itasegm1\[686\] itasegm1\[696\] itasegm1\[697\] itasegm1\[698\] itasegm1\[699\]
+ itasegm1\[687\] itasegm1\[688\] itasegm1\[689\] itasegm1\[690\] itasegm1\[691\]
+ itasegm1\[692\] itasegm1\[693\] itasegm1\[694\] itasegm1\[695\] itasel1\[588\] itasel1\[598\]
+ itasel1\[599\] itasel1\[589\] itasel1\[590\] itasel1\[591\] itasel1\[592\] itasel1\[593\]
+ itasel1\[594\] itasel1\[595\] itasel1\[596\] itasel1\[597\] vdd vss ita50
Xita2 wb_clk_i itasegm1\[14\] itasegm1\[24\] itasegm1\[25\] itasegm1\[26\] itasegm1\[27\]
+ itasegm1\[15\] itasegm1\[16\] itasegm1\[17\] itasegm1\[18\] itasegm1\[19\] itasegm1\[20\]
+ itasegm1\[21\] itasegm1\[22\] itasegm1\[23\] itasel1\[12\] itasel1\[22\] itasel1\[23\]
+ itasel1\[13\] itasel1\[14\] itasel1\[15\] itasel1\[16\] itasel1\[17\] itasel1\[18\]
+ itasel1\[19\] itasel1\[20\] itasel1\[21\] vdd vss ita2
Xita40 wb_clk_i itasegm1\[546\] itasegm1\[556\] itasegm1\[557\] itasegm1\[558\] itasegm1\[559\]
+ itasegm1\[547\] itasegm1\[548\] itasegm1\[549\] itasegm1\[550\] itasegm1\[551\]
+ itasegm1\[552\] itasegm1\[553\] itasegm1\[554\] itasegm1\[555\] itasel1\[468\] itasel1\[478\]
+ itasel1\[479\] itasel1\[469\] itasel1\[470\] itasel1\[471\] itasel1\[472\] itasel1\[473\]
+ itasel1\[474\] itasel1\[475\] itasel1\[476\] itasel1\[477\] vdd vss ita40
Xita62 wb_clk_i itasegm1\[854\] itasegm1\[864\] itasegm1\[865\] itasegm1\[866\] itasegm1\[867\]
+ itasegm1\[855\] itasegm1\[856\] itasegm1\[857\] itasegm1\[858\] itasegm1\[859\]
+ itasegm1\[860\] itasegm1\[861\] itasegm1\[862\] itasegm1\[863\] itasel1\[732\] itasel1\[742\]
+ itasel1\[743\] itasel1\[733\] itasel1\[734\] itasel1\[735\] itasel1\[736\] itasel1\[737\]
+ itasel1\[738\] itasel1\[739\] itasel1\[740\] itasel1\[741\] vdd vss ita62
Xita4 wb_clk_i itasegm1\[42\] itasegm1\[52\] itasegm1\[53\] itasegm1\[54\] itasegm1\[55\]
+ itasegm1\[43\] itasegm1\[44\] itasegm1\[45\] itasegm1\[46\] itasegm1\[47\] itasegm1\[48\]
+ itasegm1\[49\] itasegm1\[50\] itasegm1\[51\] itasel1\[36\] itasel1\[46\] itasel1\[47\]
+ itasel1\[37\] itasel1\[38\] itasel1\[39\] itasel1\[40\] itasel1\[41\] itasel1\[42\]
+ itasel1\[43\] itasel1\[44\] itasel1\[45\] vdd vss ita4
Xita51 wb_clk_i itasegm1\[700\] itasegm1\[710\] itasegm1\[711\] itasegm1\[712\] itasegm1\[713\]
+ itasegm1\[701\] itasegm1\[702\] itasegm1\[703\] itasegm1\[704\] itasegm1\[705\]
+ itasegm1\[706\] itasegm1\[707\] itasegm1\[708\] itasegm1\[709\] itasel1\[600\] itasel1\[610\]
+ itasel1\[611\] itasel1\[601\] itasel1\[602\] itasel1\[603\] itasel1\[604\] itasel1\[605\]
+ itasel1\[606\] itasel1\[607\] itasel1\[608\] itasel1\[609\] vdd vss ita51
Xita3 wb_clk_i itasegm1\[28\] itasegm1\[38\] itasegm1\[39\] itasegm1\[40\] itasegm1\[41\]
+ itasegm1\[29\] itasegm1\[30\] itasegm1\[31\] itasegm1\[32\] itasegm1\[33\] itasegm1\[34\]
+ itasegm1\[35\] itasegm1\[36\] itasegm1\[37\] itasel1\[24\] itasel1\[34\] itasel1\[35\]
+ itasel1\[25\] itasel1\[26\] itasel1\[27\] itasel1\[28\] itasel1\[29\] itasel1\[30\]
+ itasel1\[31\] itasel1\[32\] itasel1\[33\] vdd vss ita3
Xita63 wb_clk_i itasegm1\[868\] itasegm1\[878\] itasegm1\[879\] itasegm1\[880\] itasegm1\[881\]
+ itasegm1\[869\] itasegm1\[870\] itasegm1\[871\] itasegm1\[872\] itasegm1\[873\]
+ itasegm1\[874\] itasegm1\[875\] itasegm1\[876\] itasegm1\[877\] itasel1\[744\] itasel1\[754\]
+ itasel1\[755\] itasel1\[745\] itasel1\[746\] itasel1\[747\] itasel1\[748\] itasel1\[749\]
+ itasel1\[750\] itasel1\[751\] itasel1\[752\] itasel1\[753\] vdd vss ita63
Xita30 wb_clk_i itasegm1\[406\] itasegm1\[416\] itasegm1\[417\] itasegm1\[418\] itasegm1\[419\]
+ itasegm1\[407\] itasegm1\[408\] itasegm1\[409\] itasegm1\[410\] itasegm1\[411\]
+ itasegm1\[412\] itasegm1\[413\] itasegm1\[414\] itasegm1\[415\] itasel1\[348\] itasel1\[358\]
+ itasel1\[359\] itasel1\[349\] itasel1\[350\] itasel1\[351\] itasel1\[352\] itasel1\[353\]
+ itasel1\[354\] itasel1\[355\] itasel1\[356\] itasel1\[357\] vdd vss ita30
Xita5 wb_clk_i itasegm1\[56\] itasegm1\[66\] itasegm1\[67\] itasegm1\[68\] itasegm1\[69\]
+ itasegm1\[57\] itasegm1\[58\] itasegm1\[59\] itasegm1\[60\] itasegm1\[61\] itasegm1\[62\]
+ itasegm1\[63\] itasegm1\[64\] itasegm1\[65\] itasel1\[48\] itasel1\[58\] itasel1\[59\]
+ itasel1\[49\] itasel1\[50\] itasel1\[51\] itasel1\[52\] itasel1\[53\] itasel1\[54\]
+ itasel1\[55\] itasel1\[56\] itasel1\[57\] vdd vss ita5
Xita52 wb_clk_i itasegm1\[714\] itasegm1\[724\] itasegm1\[725\] itasegm1\[726\] itasegm1\[727\]
+ itasegm1\[715\] itasegm1\[716\] itasegm1\[717\] itasegm1\[718\] itasegm1\[719\]
+ itasegm1\[720\] itasegm1\[721\] itasegm1\[722\] itasegm1\[723\] itasel1\[612\] itasel1\[622\]
+ itasel1\[623\] itasel1\[613\] itasel1\[614\] itasel1\[615\] itasel1\[616\] itasel1\[617\]
+ itasel1\[618\] itasel1\[619\] itasel1\[620\] itasel1\[621\] vdd vss ita52
Xita41 wb_clk_i itasegm1\[560\] itasegm1\[570\] itasegm1\[571\] itasegm1\[572\] itasegm1\[573\]
+ itasegm1\[561\] itasegm1\[562\] itasegm1\[563\] itasegm1\[564\] itasegm1\[565\]
+ itasegm1\[566\] itasegm1\[567\] itasegm1\[568\] itasegm1\[569\] itasel1\[480\] itasel1\[490\]
+ itasel1\[491\] itasel1\[481\] itasel1\[482\] itasel1\[483\] itasel1\[484\] itasel1\[485\]
+ itasel1\[486\] itasel1\[487\] itasel1\[488\] itasel1\[489\] vdd vss ita41
Xita64 wb_clk_i itasegm1\[882\] itasegm1\[892\] itasegm1\[893\] itasegm1\[894\] itasegm1\[895\]
+ itasegm1\[883\] itasegm1\[884\] itasegm1\[885\] itasegm1\[886\] itasegm1\[887\]
+ itasegm1\[888\] itasegm1\[889\] itasegm1\[890\] itasegm1\[891\] itasel1\[756\] itasel1\[766\]
+ itasel1\[767\] itasel1\[757\] itasel1\[758\] itasel1\[759\] itasel1\[760\] itasel1\[761\]
+ itasel1\[762\] itasel1\[763\] itasel1\[764\] itasel1\[765\] vdd vss ita64
Xita31 wb_clk_i itasegm1\[420\] itasegm1\[430\] itasegm1\[431\] itasegm1\[432\] itasegm1\[433\]
+ itasegm1\[421\] itasegm1\[422\] itasegm1\[423\] itasegm1\[424\] itasegm1\[425\]
+ itasegm1\[426\] itasegm1\[427\] itasegm1\[428\] itasegm1\[429\] itasel1\[360\] itasel1\[370\]
+ itasel1\[371\] itasel1\[361\] itasel1\[362\] itasel1\[363\] itasel1\[364\] itasel1\[365\]
+ itasel1\[366\] itasel1\[367\] itasel1\[368\] itasel1\[369\] vdd vss ita31
Xita6 wb_clk_i itasegm1\[70\] itasegm1\[80\] itasegm1\[81\] itasegm1\[82\] itasegm1\[83\]
+ itasegm1\[71\] itasegm1\[72\] itasegm1\[73\] itasegm1\[74\] itasegm1\[75\] itasegm1\[76\]
+ itasegm1\[77\] itasegm1\[78\] itasegm1\[79\] itasel1\[60\] itasel1\[70\] itasel1\[71\]
+ itasel1\[61\] itasel1\[62\] itasel1\[63\] itasel1\[64\] itasel1\[65\] itasel1\[66\]
+ itasel1\[67\] itasel1\[68\] itasel1\[69\] vdd vss ita6
Xita53 wb_clk_i itasegm1\[728\] itasegm1\[738\] itasegm1\[739\] itasegm1\[740\] itasegm1\[741\]
+ itasegm1\[729\] itasegm1\[730\] itasegm1\[731\] itasegm1\[732\] itasegm1\[733\]
+ itasegm1\[734\] itasegm1\[735\] itasegm1\[736\] itasegm1\[737\] itasel1\[624\] itasel1\[634\]
+ itasel1\[635\] itasel1\[625\] itasel1\[626\] itasel1\[627\] itasel1\[628\] itasel1\[629\]
+ itasel1\[630\] itasel1\[631\] itasel1\[632\] itasel1\[633\] vdd vss ita53
Xita wb_clk_i io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14] io_oeb[15]
+ io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21] io_oeb[22]
+ io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27] io_oeb[28] io_oeb[29] io_oeb[2]
+ io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34] io_oeb[35] io_oeb[36] io_oeb[37]
+ io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9] itasegm1\[0\]
+ itasegm1\[100\] itasegm1\[101\] itasegm1\[102\] itasegm1\[103\] itasegm1\[104\]
+ itasegm1\[105\] itasegm1\[106\] itasegm1\[107\] itasegm1\[108\] itasegm1\[109\]
+ itasegm1\[10\] itasegm1\[110\] itasegm1\[111\] itasegm1\[112\] itasegm1\[113\] itasegm1\[114\]
+ itasegm1\[115\] itasegm1\[116\] itasegm1\[117\] itasegm1\[118\] itasegm1\[119\]
+ itasegm1\[11\] itasegm1\[120\] itasegm1\[121\] itasegm1\[122\] itasegm1\[123\] itasegm1\[124\]
+ itasegm1\[125\] itasegm1\[126\] itasegm1\[127\] itasegm1\[128\] itasegm1\[129\]
+ itasegm1\[12\] itasegm1\[130\] itasegm1\[131\] itasegm1\[132\] itasegm1\[133\] itasegm1\[134\]
+ itasegm1\[135\] itasegm1\[136\] itasegm1\[137\] itasegm1\[138\] itasegm1\[139\]
+ itasegm1\[13\] itasegm1\[140\] itasegm1\[141\] itasegm1\[142\] itasegm1\[143\] itasegm1\[144\]
+ itasegm1\[145\] itasegm1\[146\] itasegm1\[147\] itasegm1\[148\] itasegm1\[149\]
+ itasegm1\[14\] itasegm1\[150\] itasegm1\[151\] itasegm1\[152\] itasegm1\[153\] itasegm1\[154\]
+ itasegm1\[155\] itasegm1\[156\] itasegm1\[157\] itasegm1\[158\] itasegm1\[159\]
+ itasegm1\[15\] itasegm1\[160\] itasegm1\[161\] itasegm1\[162\] itasegm1\[163\] itasegm1\[164\]
+ itasegm1\[165\] itasegm1\[166\] itasegm1\[167\] itasegm1\[168\] itasegm1\[169\]
+ itasegm1\[16\] itasegm1\[170\] itasegm1\[171\] itasegm1\[172\] itasegm1\[173\] itasegm1\[174\]
+ itasegm1\[175\] itasegm1\[176\] itasegm1\[177\] itasegm1\[178\] itasegm1\[179\]
+ itasegm1\[17\] itasegm1\[180\] itasegm1\[181\] itasegm1\[182\] itasegm1\[183\] itasegm1\[184\]
+ itasegm1\[185\] itasegm1\[186\] itasegm1\[187\] itasegm1\[188\] itasegm1\[189\]
+ itasegm1\[18\] itasegm1\[190\] itasegm1\[191\] itasegm1\[192\] itasegm1\[193\] itasegm1\[194\]
+ itasegm1\[195\] itasegm1\[196\] itasegm1\[197\] itasegm1\[198\] itasegm1\[199\]
+ itasegm1\[19\] itasegm1\[1\] itasegm1\[200\] itasegm1\[201\] itasegm1\[202\] itasegm1\[203\]
+ itasegm1\[204\] itasegm1\[205\] itasegm1\[206\] itasegm1\[207\] itasegm1\[208\]
+ itasegm1\[209\] itasegm1\[20\] itasegm1\[210\] itasegm1\[211\] itasegm1\[212\] itasegm1\[213\]
+ itasegm1\[214\] itasegm1\[215\] itasegm1\[216\] itasegm1\[217\] itasegm1\[218\]
+ itasegm1\[219\] itasegm1\[21\] itasegm1\[220\] itasegm1\[221\] itasegm1\[222\] itasegm1\[223\]
+ itasegm1\[224\] itasegm1\[225\] itasegm1\[226\] itasegm1\[227\] itasegm1\[228\]
+ itasegm1\[229\] itasegm1\[22\] itasegm1\[230\] itasegm1\[231\] itasegm1\[232\] itasegm1\[233\]
+ itasegm1\[234\] itasegm1\[235\] itasegm1\[236\] itasegm1\[237\] itasegm1\[238\]
+ itasegm1\[239\] itasegm1\[23\] itasegm1\[240\] itasegm1\[241\] itasegm1\[242\] itasegm1\[243\]
+ itasegm1\[244\] itasegm1\[245\] itasegm1\[246\] itasegm1\[247\] itasegm1\[248\]
+ itasegm1\[249\] itasegm1\[24\] itasegm1\[250\] itasegm1\[251\] itasegm1\[252\] itasegm1\[253\]
+ itasegm1\[254\] itasegm1\[255\] itasegm1\[256\] itasegm1\[257\] itasegm1\[258\]
+ itasegm1\[259\] itasegm1\[25\] itasegm1\[260\] itasegm1\[261\] itasegm1\[262\] itasegm1\[263\]
+ itasegm1\[264\] itasegm1\[265\] itasegm1\[266\] itasegm1\[267\] itasegm1\[268\]
+ itasegm1\[269\] itasegm1\[26\] itasegm1\[270\] itasegm1\[271\] itasegm1\[272\] itasegm1\[273\]
+ itasegm1\[274\] itasegm1\[275\] itasegm1\[276\] itasegm1\[277\] itasegm1\[278\]
+ itasegm1\[279\] itasegm1\[27\] itasegm1\[280\] itasegm1\[281\] itasegm1\[282\] itasegm1\[283\]
+ itasegm1\[284\] itasegm1\[285\] itasegm1\[286\] itasegm1\[287\] itasegm1\[288\]
+ itasegm1\[289\] itasegm1\[28\] itasegm1\[290\] itasegm1\[291\] itasegm1\[292\] itasegm1\[293\]
+ itasegm1\[294\] itasegm1\[295\] itasegm1\[296\] itasegm1\[297\] itasegm1\[298\]
+ itasegm1\[299\] itasegm1\[29\] itasegm1\[2\] itasegm1\[300\] itasegm1\[301\] itasegm1\[302\]
+ itasegm1\[303\] itasegm1\[304\] itasegm1\[305\] itasegm1\[306\] itasegm1\[307\]
+ itasegm1\[308\] itasegm1\[309\] itasegm1\[30\] itasegm1\[310\] itasegm1\[311\] itasegm1\[312\]
+ itasegm1\[313\] itasegm1\[314\] itasegm1\[315\] itasegm1\[316\] itasegm1\[317\]
+ itasegm1\[318\] itasegm1\[319\] itasegm1\[31\] itasegm1\[320\] itasegm1\[321\] itasegm1\[322\]
+ itasegm1\[323\] itasegm1\[324\] itasegm1\[325\] itasegm1\[326\] itasegm1\[327\]
+ itasegm1\[328\] itasegm1\[329\] itasegm1\[32\] itasegm1\[330\] itasegm1\[331\] itasegm1\[332\]
+ itasegm1\[333\] itasegm1\[334\] itasegm1\[335\] itasegm1\[336\] itasegm1\[337\]
+ itasegm1\[338\] itasegm1\[339\] itasegm1\[33\] itasegm1\[340\] itasegm1\[341\] itasegm1\[342\]
+ itasegm1\[343\] itasegm1\[344\] itasegm1\[345\] itasegm1\[346\] itasegm1\[347\]
+ itasegm1\[348\] itasegm1\[349\] itasegm1\[34\] itasegm1\[350\] itasegm1\[351\] itasegm1\[352\]
+ itasegm1\[353\] itasegm1\[354\] itasegm1\[355\] itasegm1\[356\] itasegm1\[357\]
+ itasegm1\[358\] itasegm1\[359\] itasegm1\[35\] itasegm1\[360\] itasegm1\[361\] itasegm1\[362\]
+ itasegm1\[363\] itasegm1\[364\] itasegm1\[365\] itasegm1\[366\] itasegm1\[367\]
+ itasegm1\[368\] itasegm1\[369\] itasegm1\[36\] itasegm1\[370\] itasegm1\[371\] itasegm1\[372\]
+ itasegm1\[373\] itasegm1\[374\] itasegm1\[375\] itasegm1\[376\] itasegm1\[377\]
+ itasegm1\[378\] itasegm1\[379\] itasegm1\[37\] itasegm1\[380\] itasegm1\[381\] itasegm1\[382\]
+ itasegm1\[383\] itasegm1\[384\] itasegm1\[385\] itasegm1\[386\] itasegm1\[387\]
+ itasegm1\[388\] itasegm1\[389\] itasegm1\[38\] itasegm1\[390\] itasegm1\[391\] itasegm1\[392\]
+ itasegm1\[393\] itasegm1\[394\] itasegm1\[395\] itasegm1\[396\] itasegm1\[397\]
+ itasegm1\[398\] itasegm1\[399\] itasegm1\[39\] itasegm1\[3\] itasegm1\[400\] itasegm1\[401\]
+ itasegm1\[402\] itasegm1\[403\] itasegm1\[404\] itasegm1\[405\] itasegm1\[406\]
+ itasegm1\[407\] itasegm1\[408\] itasegm1\[409\] itasegm1\[40\] itasegm1\[410\] itasegm1\[411\]
+ itasegm1\[412\] itasegm1\[413\] itasegm1\[414\] itasegm1\[415\] itasegm1\[416\]
+ itasegm1\[417\] itasegm1\[418\] itasegm1\[419\] itasegm1\[41\] itasegm1\[420\] itasegm1\[421\]
+ itasegm1\[422\] itasegm1\[423\] itasegm1\[424\] itasegm1\[425\] itasegm1\[426\]
+ itasegm1\[427\] itasegm1\[428\] itasegm1\[429\] itasegm1\[42\] itasegm1\[430\] itasegm1\[431\]
+ itasegm1\[432\] itasegm1\[433\] itasegm1\[434\] itasegm1\[435\] itasegm1\[436\]
+ itasegm1\[437\] itasegm1\[438\] itasegm1\[439\] itasegm1\[43\] itasegm1\[440\] itasegm1\[441\]
+ itasegm1\[442\] itasegm1\[443\] itasegm1\[444\] itasegm1\[445\] itasegm1\[446\]
+ itasegm1\[447\] itasegm1\[448\] itasegm1\[449\] itasegm1\[44\] itasegm1\[450\] itasegm1\[451\]
+ itasegm1\[452\] itasegm1\[453\] itasegm1\[454\] itasegm1\[455\] itasegm1\[456\]
+ itasegm1\[457\] itasegm1\[458\] itasegm1\[459\] itasegm1\[45\] itasegm1\[460\] itasegm1\[461\]
+ itasegm1\[462\] itasegm1\[463\] itasegm1\[464\] itasegm1\[465\] itasegm1\[466\]
+ itasegm1\[467\] itasegm1\[468\] itasegm1\[469\] itasegm1\[46\] itasegm1\[470\] itasegm1\[471\]
+ itasegm1\[472\] itasegm1\[473\] itasegm1\[474\] itasegm1\[475\] itasegm1\[476\]
+ itasegm1\[477\] itasegm1\[478\] itasegm1\[479\] itasegm1\[47\] itasegm1\[480\] itasegm1\[481\]
+ itasegm1\[482\] itasegm1\[483\] itasegm1\[484\] itasegm1\[485\] itasegm1\[486\]
+ itasegm1\[487\] itasegm1\[488\] itasegm1\[489\] itasegm1\[48\] itasegm1\[490\] itasegm1\[491\]
+ itasegm1\[492\] itasegm1\[493\] itasegm1\[494\] itasegm1\[495\] itasegm1\[496\]
+ itasegm1\[497\] itasegm1\[498\] itasegm1\[499\] itasegm1\[49\] itasegm1\[4\] itasegm1\[500\]
+ itasegm1\[501\] itasegm1\[502\] itasegm1\[503\] itasegm1\[504\] itasegm1\[505\]
+ itasegm1\[506\] itasegm1\[507\] itasegm1\[508\] itasegm1\[509\] itasegm1\[50\] itasegm1\[510\]
+ itasegm1\[511\] itasegm1\[512\] itasegm1\[513\] itasegm1\[514\] itasegm1\[515\]
+ itasegm1\[516\] itasegm1\[517\] itasegm1\[518\] itasegm1\[519\] itasegm1\[51\] itasegm1\[520\]
+ itasegm1\[521\] itasegm1\[522\] itasegm1\[523\] itasegm1\[524\] itasegm1\[525\]
+ itasegm1\[526\] itasegm1\[527\] itasegm1\[528\] itasegm1\[529\] itasegm1\[52\] itasegm1\[530\]
+ itasegm1\[531\] itasegm1\[532\] itasegm1\[533\] itasegm1\[534\] itasegm1\[535\]
+ itasegm1\[536\] itasegm1\[537\] itasegm1\[538\] itasegm1\[539\] itasegm1\[53\] itasegm1\[540\]
+ itasegm1\[541\] itasegm1\[542\] itasegm1\[543\] itasegm1\[544\] itasegm1\[545\]
+ itasegm1\[546\] itasegm1\[547\] itasegm1\[548\] itasegm1\[549\] itasegm1\[54\] itasegm1\[550\]
+ itasegm1\[551\] itasegm1\[552\] itasegm1\[553\] itasegm1\[554\] itasegm1\[555\]
+ itasegm1\[556\] itasegm1\[557\] itasegm1\[558\] itasegm1\[559\] itasegm1\[55\] itasegm1\[560\]
+ itasegm1\[561\] itasegm1\[562\] itasegm1\[563\] itasegm1\[564\] itasegm1\[565\]
+ itasegm1\[566\] itasegm1\[567\] itasegm1\[568\] itasegm1\[569\] itasegm1\[56\] itasegm1\[570\]
+ itasegm1\[571\] itasegm1\[572\] itasegm1\[573\] itasegm1\[574\] itasegm1\[575\]
+ itasegm1\[576\] itasegm1\[577\] itasegm1\[578\] itasegm1\[579\] itasegm1\[57\] itasegm1\[580\]
+ itasegm1\[581\] itasegm1\[582\] itasegm1\[583\] itasegm1\[584\] itasegm1\[585\]
+ itasegm1\[586\] itasegm1\[587\] itasegm1\[588\] itasegm1\[589\] itasegm1\[58\] itasegm1\[590\]
+ itasegm1\[591\] itasegm1\[592\] itasegm1\[593\] itasegm1\[594\] itasegm1\[595\]
+ itasegm1\[596\] itasegm1\[597\] itasegm1\[598\] itasegm1\[599\] itasegm1\[59\] itasegm1\[5\]
+ itasegm1\[600\] itasegm1\[601\] itasegm1\[602\] itasegm1\[603\] itasegm1\[604\]
+ itasegm1\[605\] itasegm1\[606\] itasegm1\[607\] itasegm1\[608\] itasegm1\[609\]
+ itasegm1\[60\] itasegm1\[610\] itasegm1\[611\] itasegm1\[612\] itasegm1\[613\] itasegm1\[614\]
+ itasegm1\[615\] itasegm1\[616\] itasegm1\[617\] itasegm1\[618\] itasegm1\[619\]
+ itasegm1\[61\] itasegm1\[620\] itasegm1\[621\] itasegm1\[622\] itasegm1\[623\] itasegm1\[624\]
+ itasegm1\[625\] itasegm1\[626\] itasegm1\[627\] itasegm1\[628\] itasegm1\[629\]
+ itasegm1\[62\] itasegm1\[630\] itasegm1\[631\] itasegm1\[632\] itasegm1\[633\] itasegm1\[634\]
+ itasegm1\[635\] itasegm1\[636\] itasegm1\[637\] itasegm1\[638\] itasegm1\[639\]
+ itasegm1\[63\] itasegm1\[640\] itasegm1\[641\] itasegm1\[642\] itasegm1\[643\] itasegm1\[644\]
+ itasegm1\[645\] itasegm1\[646\] itasegm1\[647\] itasegm1\[648\] itasegm1\[649\]
+ itasegm1\[64\] itasegm1\[650\] itasegm1\[651\] itasegm1\[652\] itasegm1\[653\] itasegm1\[654\]
+ itasegm1\[655\] itasegm1\[656\] itasegm1\[657\] itasegm1\[658\] itasegm1\[659\]
+ itasegm1\[65\] itasegm1\[660\] itasegm1\[661\] itasegm1\[662\] itasegm1\[663\] itasegm1\[664\]
+ itasegm1\[665\] itasegm1\[666\] itasegm1\[667\] itasegm1\[668\] itasegm1\[669\]
+ itasegm1\[66\] itasegm1\[670\] itasegm1\[671\] itasegm1\[672\] itasegm1\[673\] itasegm1\[674\]
+ itasegm1\[675\] itasegm1\[676\] itasegm1\[677\] itasegm1\[678\] itasegm1\[679\]
+ itasegm1\[67\] itasegm1\[680\] itasegm1\[681\] itasegm1\[682\] itasegm1\[683\] itasegm1\[684\]
+ itasegm1\[685\] itasegm1\[686\] itasegm1\[687\] itasegm1\[688\] itasegm1\[689\]
+ itasegm1\[68\] itasegm1\[690\] itasegm1\[691\] itasegm1\[692\] itasegm1\[693\] itasegm1\[694\]
+ itasegm1\[695\] itasegm1\[696\] itasegm1\[697\] itasegm1\[698\] itasegm1\[699\]
+ itasegm1\[69\] itasegm1\[6\] itasegm1\[700\] itasegm1\[701\] itasegm1\[702\] itasegm1\[703\]
+ itasegm1\[704\] itasegm1\[705\] itasegm1\[706\] itasegm1\[707\] itasegm1\[708\]
+ itasegm1\[709\] itasegm1\[70\] itasegm1\[710\] itasegm1\[711\] itasegm1\[712\] itasegm1\[713\]
+ itasegm1\[714\] itasegm1\[715\] itasegm1\[716\] itasegm1\[717\] itasegm1\[718\]
+ itasegm1\[719\] itasegm1\[71\] itasegm1\[720\] itasegm1\[721\] itasegm1\[722\] itasegm1\[723\]
+ itasegm1\[724\] itasegm1\[725\] itasegm1\[726\] itasegm1\[727\] itasegm1\[728\]
+ itasegm1\[729\] itasegm1\[72\] itasegm1\[730\] itasegm1\[731\] itasegm1\[732\] itasegm1\[733\]
+ itasegm1\[734\] itasegm1\[735\] itasegm1\[736\] itasegm1\[737\] itasegm1\[738\]
+ itasegm1\[739\] itasegm1\[73\] itasegm1\[740\] itasegm1\[741\] itasegm1\[742\] itasegm1\[743\]
+ itasegm1\[744\] itasegm1\[745\] itasegm1\[746\] itasegm1\[747\] itasegm1\[748\]
+ itasegm1\[749\] itasegm1\[74\] itasegm1\[750\] itasegm1\[751\] itasegm1\[752\] itasegm1\[753\]
+ itasegm1\[754\] itasegm1\[755\] itasegm1\[756\] itasegm1\[757\] itasegm1\[758\]
+ itasegm1\[759\] itasegm1\[75\] itasegm1\[760\] itasegm1\[761\] itasegm1\[762\] itasegm1\[763\]
+ itasegm1\[764\] itasegm1\[765\] itasegm1\[766\] itasegm1\[767\] itasegm1\[768\]
+ itasegm1\[769\] itasegm1\[76\] itasegm1\[770\] itasegm1\[771\] itasegm1\[772\] itasegm1\[773\]
+ itasegm1\[774\] itasegm1\[775\] itasegm1\[776\] itasegm1\[777\] itasegm1\[778\]
+ itasegm1\[779\] itasegm1\[77\] itasegm1\[780\] itasegm1\[781\] itasegm1\[782\] itasegm1\[783\]
+ itasegm1\[784\] itasegm1\[785\] itasegm1\[786\] itasegm1\[787\] itasegm1\[788\]
+ itasegm1\[789\] itasegm1\[78\] itasegm1\[790\] itasegm1\[791\] itasegm1\[792\] itasegm1\[793\]
+ itasegm1\[794\] itasegm1\[795\] itasegm1\[796\] itasegm1\[797\] itasegm1\[798\]
+ itasegm1\[799\] itasegm1\[79\] itasegm1\[7\] itasegm1\[800\] itasegm1\[801\] itasegm1\[802\]
+ itasegm1\[803\] itasegm1\[804\] itasegm1\[805\] itasegm1\[806\] itasegm1\[807\]
+ itasegm1\[808\] itasegm1\[809\] itasegm1\[80\] itasegm1\[810\] itasegm1\[811\] itasegm1\[812\]
+ itasegm1\[813\] itasegm1\[814\] itasegm1\[815\] itasegm1\[816\] itasegm1\[817\]
+ itasegm1\[818\] itasegm1\[819\] itasegm1\[81\] itasegm1\[820\] itasegm1\[821\] itasegm1\[822\]
+ itasegm1\[823\] itasegm1\[824\] itasegm1\[825\] itasegm1\[826\] itasegm1\[827\]
+ itasegm1\[828\] itasegm1\[829\] itasegm1\[82\] itasegm1\[830\] itasegm1\[831\] itasegm1\[832\]
+ itasegm1\[833\] itasegm1\[834\] itasegm1\[835\] itasegm1\[836\] itasegm1\[837\]
+ itasegm1\[838\] itasegm1\[839\] itasegm1\[83\] itasegm1\[840\] itasegm1\[841\] itasegm1\[842\]
+ itasegm1\[843\] itasegm1\[844\] itasegm1\[845\] itasegm1\[846\] itasegm1\[847\]
+ itasegm1\[848\] itasegm1\[849\] itasegm1\[84\] itasegm1\[850\] itasegm1\[851\] itasegm1\[852\]
+ itasegm1\[853\] itasegm1\[854\] itasegm1\[855\] itasegm1\[856\] itasegm1\[857\]
+ itasegm1\[858\] itasegm1\[859\] itasegm1\[85\] itasegm1\[860\] itasegm1\[861\] itasegm1\[862\]
+ itasegm1\[863\] itasegm1\[864\] itasegm1\[865\] itasegm1\[866\] itasegm1\[867\]
+ itasegm1\[868\] itasegm1\[869\] itasegm1\[86\] itasegm1\[870\] itasegm1\[871\] itasegm1\[872\]
+ itasegm1\[873\] itasegm1\[874\] itasegm1\[875\] itasegm1\[876\] itasegm1\[877\]
+ itasegm1\[878\] itasegm1\[879\] itasegm1\[87\] itasegm1\[880\] itasegm1\[881\] itasegm1\[882\]
+ itasegm1\[883\] itasegm1\[884\] itasegm1\[885\] itasegm1\[886\] itasegm1\[887\]
+ itasegm1\[888\] itasegm1\[889\] itasegm1\[88\] itasegm1\[890\] itasegm1\[891\] itasegm1\[892\]
+ itasegm1\[893\] itasegm1\[894\] itasegm1\[895\] itasegm1\[89\] itasegm1\[8\] itasegm1\[90\]
+ itasegm1\[91\] itasegm1\[92\] itasegm1\[93\] itasegm1\[94\] itasegm1\[95\] itasegm1\[96\]
+ itasegm1\[97\] itasegm1\[98\] itasegm1\[99\] itasegm1\[9\] itasel1\[0\] itasel1\[100\]
+ itasel1\[101\] itasel1\[102\] itasel1\[103\] itasel1\[104\] itasel1\[105\] itasel1\[106\]
+ itasel1\[107\] itasel1\[108\] itasel1\[109\] itasel1\[10\] itasel1\[110\] itasel1\[111\]
+ itasel1\[112\] itasel1\[113\] itasel1\[114\] itasel1\[115\] itasel1\[116\] itasel1\[117\]
+ itasel1\[118\] itasel1\[119\] itasel1\[11\] itasel1\[120\] itasel1\[121\] itasel1\[122\]
+ itasel1\[123\] itasel1\[124\] itasel1\[125\] itasel1\[126\] itasel1\[127\] itasel1\[128\]
+ itasel1\[129\] itasel1\[12\] itasel1\[130\] itasel1\[131\] itasel1\[132\] itasel1\[133\]
+ itasel1\[134\] itasel1\[135\] itasel1\[136\] itasel1\[137\] itasel1\[138\] itasel1\[139\]
+ itasel1\[13\] itasel1\[140\] itasel1\[141\] itasel1\[142\] itasel1\[143\] itasel1\[144\]
+ itasel1\[145\] itasel1\[146\] itasel1\[147\] itasel1\[148\] itasel1\[149\] itasel1\[14\]
+ itasel1\[150\] itasel1\[151\] itasel1\[152\] itasel1\[153\] itasel1\[154\] itasel1\[155\]
+ itasel1\[156\] itasel1\[157\] itasel1\[158\] itasel1\[159\] itasel1\[15\] itasel1\[160\]
+ itasel1\[161\] itasel1\[162\] itasel1\[163\] itasel1\[164\] itasel1\[165\] itasel1\[166\]
+ itasel1\[167\] itasel1\[168\] itasel1\[169\] itasel1\[16\] itasel1\[170\] itasel1\[171\]
+ itasel1\[172\] itasel1\[173\] itasel1\[174\] itasel1\[175\] itasel1\[176\] itasel1\[177\]
+ itasel1\[178\] itasel1\[179\] itasel1\[17\] itasel1\[180\] itasel1\[181\] itasel1\[182\]
+ itasel1\[183\] itasel1\[184\] itasel1\[185\] itasel1\[186\] itasel1\[187\] itasel1\[188\]
+ itasel1\[189\] itasel1\[18\] itasel1\[190\] itasel1\[191\] itasel1\[192\] itasel1\[193\]
+ itasel1\[194\] itasel1\[195\] itasel1\[196\] itasel1\[197\] itasel1\[198\] itasel1\[199\]
+ itasel1\[19\] itasel1\[1\] itasel1\[200\] itasel1\[201\] itasel1\[202\] itasel1\[203\]
+ itasel1\[204\] itasel1\[205\] itasel1\[206\] itasel1\[207\] itasel1\[208\] itasel1\[209\]
+ itasel1\[20\] itasel1\[210\] itasel1\[211\] itasel1\[212\] itasel1\[213\] itasel1\[214\]
+ itasel1\[215\] itasel1\[216\] itasel1\[217\] itasel1\[218\] itasel1\[219\] itasel1\[21\]
+ itasel1\[220\] itasel1\[221\] itasel1\[222\] itasel1\[223\] itasel1\[224\] itasel1\[225\]
+ itasel1\[226\] itasel1\[227\] itasel1\[228\] itasel1\[229\] itasel1\[22\] itasel1\[230\]
+ itasel1\[231\] itasel1\[232\] itasel1\[233\] itasel1\[234\] itasel1\[235\] itasel1\[236\]
+ itasel1\[237\] itasel1\[238\] itasel1\[239\] itasel1\[23\] itasel1\[240\] itasel1\[241\]
+ itasel1\[242\] itasel1\[243\] itasel1\[244\] itasel1\[245\] itasel1\[246\] itasel1\[247\]
+ itasel1\[248\] itasel1\[249\] itasel1\[24\] itasel1\[250\] itasel1\[251\] itasel1\[252\]
+ itasel1\[253\] itasel1\[254\] itasel1\[255\] itasel1\[256\] itasel1\[257\] itasel1\[258\]
+ itasel1\[259\] itasel1\[25\] itasel1\[260\] itasel1\[261\] itasel1\[262\] itasel1\[263\]
+ itasel1\[264\] itasel1\[265\] itasel1\[266\] itasel1\[267\] itasel1\[268\] itasel1\[269\]
+ itasel1\[26\] itasel1\[270\] itasel1\[271\] itasel1\[272\] itasel1\[273\] itasel1\[274\]
+ itasel1\[275\] itasel1\[276\] itasel1\[277\] itasel1\[278\] itasel1\[279\] itasel1\[27\]
+ itasel1\[280\] itasel1\[281\] itasel1\[282\] itasel1\[283\] itasel1\[284\] itasel1\[285\]
+ itasel1\[286\] itasel1\[287\] itasel1\[288\] itasel1\[289\] itasel1\[28\] itasel1\[290\]
+ itasel1\[291\] itasel1\[292\] itasel1\[293\] itasel1\[294\] itasel1\[295\] itasel1\[296\]
+ itasel1\[297\] itasel1\[298\] itasel1\[299\] itasel1\[29\] itasel1\[2\] itasel1\[300\]
+ itasel1\[301\] itasel1\[302\] itasel1\[303\] itasel1\[304\] itasel1\[305\] itasel1\[306\]
+ itasel1\[307\] itasel1\[308\] itasel1\[309\] itasel1\[30\] itasel1\[310\] itasel1\[311\]
+ itasel1\[312\] itasel1\[313\] itasel1\[314\] itasel1\[315\] itasel1\[316\] itasel1\[317\]
+ itasel1\[318\] itasel1\[319\] itasel1\[31\] itasel1\[320\] itasel1\[321\] itasel1\[322\]
+ itasel1\[323\] itasel1\[324\] itasel1\[325\] itasel1\[326\] itasel1\[327\] itasel1\[328\]
+ itasel1\[329\] itasel1\[32\] itasel1\[330\] itasel1\[331\] itasel1\[332\] itasel1\[333\]
+ itasel1\[334\] itasel1\[335\] itasel1\[336\] itasel1\[337\] itasel1\[338\] itasel1\[339\]
+ itasel1\[33\] itasel1\[340\] itasel1\[341\] itasel1\[342\] itasel1\[343\] itasel1\[344\]
+ itasel1\[345\] itasel1\[346\] itasel1\[347\] itasel1\[348\] itasel1\[349\] itasel1\[34\]
+ itasel1\[350\] itasel1\[351\] itasel1\[352\] itasel1\[353\] itasel1\[354\] itasel1\[355\]
+ itasel1\[356\] itasel1\[357\] itasel1\[358\] itasel1\[359\] itasel1\[35\] itasel1\[360\]
+ itasel1\[361\] itasel1\[362\] itasel1\[363\] itasel1\[364\] itasel1\[365\] itasel1\[366\]
+ itasel1\[367\] itasel1\[368\] itasel1\[369\] itasel1\[36\] itasel1\[370\] itasel1\[371\]
+ itasel1\[372\] itasel1\[373\] itasel1\[374\] itasel1\[375\] itasel1\[376\] itasel1\[377\]
+ itasel1\[378\] itasel1\[379\] itasel1\[37\] itasel1\[380\] itasel1\[381\] itasel1\[382\]
+ itasel1\[383\] itasel1\[384\] itasel1\[385\] itasel1\[386\] itasel1\[387\] itasel1\[388\]
+ itasel1\[389\] itasel1\[38\] itasel1\[390\] itasel1\[391\] itasel1\[392\] itasel1\[393\]
+ itasel1\[394\] itasel1\[395\] itasel1\[396\] itasel1\[397\] itasel1\[398\] itasel1\[399\]
+ itasel1\[39\] itasel1\[3\] itasel1\[400\] itasel1\[401\] itasel1\[402\] itasel1\[403\]
+ itasel1\[404\] itasel1\[405\] itasel1\[406\] itasel1\[407\] itasel1\[408\] itasel1\[409\]
+ itasel1\[40\] itasel1\[410\] itasel1\[411\] itasel1\[412\] itasel1\[413\] itasel1\[414\]
+ itasel1\[415\] itasel1\[416\] itasel1\[417\] itasel1\[418\] itasel1\[419\] itasel1\[41\]
+ itasel1\[420\] itasel1\[421\] itasel1\[422\] itasel1\[423\] itasel1\[424\] itasel1\[425\]
+ itasel1\[426\] itasel1\[427\] itasel1\[428\] itasel1\[429\] itasel1\[42\] itasel1\[430\]
+ itasel1\[431\] itasel1\[432\] itasel1\[433\] itasel1\[434\] itasel1\[435\] itasel1\[436\]
+ itasel1\[437\] itasel1\[438\] itasel1\[439\] itasel1\[43\] itasel1\[440\] itasel1\[441\]
+ itasel1\[442\] itasel1\[443\] itasel1\[444\] itasel1\[445\] itasel1\[446\] itasel1\[447\]
+ itasel1\[448\] itasel1\[449\] itasel1\[44\] itasel1\[450\] itasel1\[451\] itasel1\[452\]
+ itasel1\[453\] itasel1\[454\] itasel1\[455\] itasel1\[456\] itasel1\[457\] itasel1\[458\]
+ itasel1\[459\] itasel1\[45\] itasel1\[460\] itasel1\[461\] itasel1\[462\] itasel1\[463\]
+ itasel1\[464\] itasel1\[465\] itasel1\[466\] itasel1\[467\] itasel1\[468\] itasel1\[469\]
+ itasel1\[46\] itasel1\[470\] itasel1\[471\] itasel1\[472\] itasel1\[473\] itasel1\[474\]
+ itasel1\[475\] itasel1\[476\] itasel1\[477\] itasel1\[478\] itasel1\[479\] itasel1\[47\]
+ itasel1\[480\] itasel1\[481\] itasel1\[482\] itasel1\[483\] itasel1\[484\] itasel1\[485\]
+ itasel1\[486\] itasel1\[487\] itasel1\[488\] itasel1\[489\] itasel1\[48\] itasel1\[490\]
+ itasel1\[491\] itasel1\[492\] itasel1\[493\] itasel1\[494\] itasel1\[495\] itasel1\[496\]
+ itasel1\[497\] itasel1\[498\] itasel1\[499\] itasel1\[49\] itasel1\[4\] itasel1\[500\]
+ itasel1\[501\] itasel1\[502\] itasel1\[503\] itasel1\[504\] itasel1\[505\] itasel1\[506\]
+ itasel1\[507\] itasel1\[508\] itasel1\[509\] itasel1\[50\] itasel1\[510\] itasel1\[511\]
+ itasel1\[512\] itasel1\[513\] itasel1\[514\] itasel1\[515\] itasel1\[516\] itasel1\[517\]
+ itasel1\[518\] itasel1\[519\] itasel1\[51\] itasel1\[520\] itasel1\[521\] itasel1\[522\]
+ itasel1\[523\] itasel1\[524\] itasel1\[525\] itasel1\[526\] itasel1\[527\] itasel1\[528\]
+ itasel1\[529\] itasel1\[52\] itasel1\[530\] itasel1\[531\] itasel1\[532\] itasel1\[533\]
+ itasel1\[534\] itasel1\[535\] itasel1\[536\] itasel1\[537\] itasel1\[538\] itasel1\[539\]
+ itasel1\[53\] itasel1\[540\] itasel1\[541\] itasel1\[542\] itasel1\[543\] itasel1\[544\]
+ itasel1\[545\] itasel1\[546\] itasel1\[547\] itasel1\[548\] itasel1\[549\] itasel1\[54\]
+ itasel1\[550\] itasel1\[551\] itasel1\[552\] itasel1\[553\] itasel1\[554\] itasel1\[555\]
+ itasel1\[556\] itasel1\[557\] itasel1\[558\] itasel1\[559\] itasel1\[55\] itasel1\[560\]
+ itasel1\[561\] itasel1\[562\] itasel1\[563\] itasel1\[564\] itasel1\[565\] itasel1\[566\]
+ itasel1\[567\] itasel1\[568\] itasel1\[569\] itasel1\[56\] itasel1\[570\] itasel1\[571\]
+ itasel1\[572\] itasel1\[573\] itasel1\[574\] itasel1\[575\] itasel1\[576\] itasel1\[577\]
+ itasel1\[578\] itasel1\[579\] itasel1\[57\] itasel1\[580\] itasel1\[581\] itasel1\[582\]
+ itasel1\[583\] itasel1\[584\] itasel1\[585\] itasel1\[586\] itasel1\[587\] itasel1\[588\]
+ itasel1\[589\] itasel1\[58\] itasel1\[590\] itasel1\[591\] itasel1\[592\] itasel1\[593\]
+ itasel1\[594\] itasel1\[595\] itasel1\[596\] itasel1\[597\] itasel1\[598\] itasel1\[599\]
+ itasel1\[59\] itasel1\[5\] itasel1\[600\] itasel1\[601\] itasel1\[602\] itasel1\[603\]
+ itasel1\[604\] itasel1\[605\] itasel1\[606\] itasel1\[607\] itasel1\[608\] itasel1\[609\]
+ itasel1\[60\] itasel1\[610\] itasel1\[611\] itasel1\[612\] itasel1\[613\] itasel1\[614\]
+ itasel1\[615\] itasel1\[616\] itasel1\[617\] itasel1\[618\] itasel1\[619\] itasel1\[61\]
+ itasel1\[620\] itasel1\[621\] itasel1\[622\] itasel1\[623\] itasel1\[624\] itasel1\[625\]
+ itasel1\[626\] itasel1\[627\] itasel1\[628\] itasel1\[629\] itasel1\[62\] itasel1\[630\]
+ itasel1\[631\] itasel1\[632\] itasel1\[633\] itasel1\[634\] itasel1\[635\] itasel1\[636\]
+ itasel1\[637\] itasel1\[638\] itasel1\[639\] itasel1\[63\] itasel1\[640\] itasel1\[641\]
+ itasel1\[642\] itasel1\[643\] itasel1\[644\] itasel1\[645\] itasel1\[646\] itasel1\[647\]
+ itasel1\[648\] itasel1\[649\] itasel1\[64\] itasel1\[650\] itasel1\[651\] itasel1\[652\]
+ itasel1\[653\] itasel1\[654\] itasel1\[655\] itasel1\[656\] itasel1\[657\] itasel1\[658\]
+ itasel1\[659\] itasel1\[65\] itasel1\[660\] itasel1\[661\] itasel1\[662\] itasel1\[663\]
+ itasel1\[664\] itasel1\[665\] itasel1\[666\] itasel1\[667\] itasel1\[668\] itasel1\[669\]
+ itasel1\[66\] itasel1\[670\] itasel1\[671\] itasel1\[672\] itasel1\[673\] itasel1\[674\]
+ itasel1\[675\] itasel1\[676\] itasel1\[677\] itasel1\[678\] itasel1\[679\] itasel1\[67\]
+ itasel1\[680\] itasel1\[681\] itasel1\[682\] itasel1\[683\] itasel1\[684\] itasel1\[685\]
+ itasel1\[686\] itasel1\[687\] itasel1\[688\] itasel1\[689\] itasel1\[68\] itasel1\[690\]
+ itasel1\[691\] itasel1\[692\] itasel1\[693\] itasel1\[694\] itasel1\[695\] itasel1\[696\]
+ itasel1\[697\] itasel1\[698\] itasel1\[699\] itasel1\[69\] itasel1\[6\] itasel1\[700\]
+ itasel1\[701\] itasel1\[702\] itasel1\[703\] itasel1\[704\] itasel1\[705\] itasel1\[706\]
+ itasel1\[707\] itasel1\[708\] itasel1\[709\] itasel1\[70\] itasel1\[710\] itasel1\[711\]
+ itasel1\[712\] itasel1\[713\] itasel1\[714\] itasel1\[715\] itasel1\[716\] itasel1\[717\]
+ itasel1\[718\] itasel1\[719\] itasel1\[71\] itasel1\[720\] itasel1\[721\] itasel1\[722\]
+ itasel1\[723\] itasel1\[724\] itasel1\[725\] itasel1\[726\] itasel1\[727\] itasel1\[728\]
+ itasel1\[729\] itasel1\[72\] itasel1\[730\] itasel1\[731\] itasel1\[732\] itasel1\[733\]
+ itasel1\[734\] itasel1\[735\] itasel1\[736\] itasel1\[737\] itasel1\[738\] itasel1\[739\]
+ itasel1\[73\] itasel1\[740\] itasel1\[741\] itasel1\[742\] itasel1\[743\] itasel1\[744\]
+ itasel1\[745\] itasel1\[746\] itasel1\[747\] itasel1\[748\] itasel1\[749\] itasel1\[74\]
+ itasel1\[750\] itasel1\[751\] itasel1\[752\] itasel1\[753\] itasel1\[754\] itasel1\[755\]
+ itasel1\[756\] itasel1\[757\] itasel1\[758\] itasel1\[759\] itasel1\[75\] itasel1\[760\]
+ itasel1\[761\] itasel1\[762\] itasel1\[763\] itasel1\[764\] itasel1\[765\] itasel1\[766\]
+ itasel1\[767\] itasel1\[76\] itasel1\[77\] itasel1\[78\] itasel1\[79\] itasel1\[7\]
+ itasel1\[80\] itasel1\[81\] itasel1\[82\] itasel1\[83\] itasel1\[84\] itasel1\[85\]
+ itasel1\[86\] itasel1\[87\] itasel1\[88\] itasel1\[89\] itasel1\[8\] itasel1\[90\]
+ itasel1\[91\] itasel1\[92\] itasel1\[93\] itasel1\[94\] itasel1\[95\] itasel1\[96\]
+ itasel1\[97\] itasel1\[98\] itasel1\[99\] itasel1\[9\] io_in[6] io_in[7] io_in[8]
+ io_in[9] io_in[10] io_in[11] io_out[24] io_out[34] io_out[35] io_out[36] io_out[37]
+ io_out[25] io_out[26] io_out[27] io_out[28] io_out[29] io_out[30] io_out[31] io_out[32]
+ io_out[33] io_out[12] io_out[22] io_out[23] io_out[13] io_out[14] io_out[15] io_out[16]
+ io_out[17] io_out[18] io_out[19] io_out[20] io_out[21] vdd vss ita
Xita20 wb_clk_i itasegm1\[266\] itasegm1\[276\] itasegm1\[277\] itasegm1\[278\] itasegm1\[279\]
+ itasegm1\[267\] itasegm1\[268\] itasegm1\[269\] itasegm1\[270\] itasegm1\[271\]
+ itasegm1\[272\] itasegm1\[273\] itasegm1\[274\] itasegm1\[275\] itasel1\[228\] itasel1\[238\]
+ itasel1\[239\] itasel1\[229\] itasel1\[230\] itasel1\[231\] itasel1\[232\] itasel1\[233\]
+ itasel1\[234\] itasel1\[235\] itasel1\[236\] itasel1\[237\] vdd vss ita20
Xita42 wb_clk_i itasegm1\[574\] itasegm1\[584\] itasegm1\[585\] itasegm1\[586\] itasegm1\[587\]
+ itasegm1\[575\] itasegm1\[576\] itasegm1\[577\] itasegm1\[578\] itasegm1\[579\]
+ itasegm1\[580\] itasegm1\[581\] itasegm1\[582\] itasegm1\[583\] itasel1\[492\] itasel1\[502\]
+ itasel1\[503\] itasel1\[493\] itasel1\[494\] itasel1\[495\] itasel1\[496\] itasel1\[497\]
+ itasel1\[498\] itasel1\[499\] itasel1\[500\] itasel1\[501\] vdd vss ita42
Xita32 wb_clk_i itasegm1\[434\] itasegm1\[444\] itasegm1\[445\] itasegm1\[446\] itasegm1\[447\]
+ itasegm1\[435\] itasegm1\[436\] itasegm1\[437\] itasegm1\[438\] itasegm1\[439\]
+ itasegm1\[440\] itasegm1\[441\] itasegm1\[442\] itasegm1\[443\] itasel1\[372\] itasel1\[382\]
+ itasel1\[383\] itasel1\[373\] itasel1\[374\] itasel1\[375\] itasel1\[376\] itasel1\[377\]
+ itasel1\[378\] itasel1\[379\] itasel1\[380\] itasel1\[381\] vdd vss ita32
Xita7 wb_clk_i itasegm1\[84\] itasegm1\[94\] itasegm1\[95\] itasegm1\[96\] itasegm1\[97\]
+ itasegm1\[85\] itasegm1\[86\] itasegm1\[87\] itasegm1\[88\] itasegm1\[89\] itasegm1\[90\]
+ itasegm1\[91\] itasegm1\[92\] itasegm1\[93\] itasel1\[72\] itasel1\[82\] itasel1\[83\]
+ itasel1\[73\] itasel1\[74\] itasel1\[75\] itasel1\[76\] itasel1\[77\] itasel1\[78\]
+ itasel1\[79\] itasel1\[80\] itasel1\[81\] vdd vss ita7
Xita54 wb_clk_i itasegm1\[742\] itasegm1\[752\] itasegm1\[753\] itasegm1\[754\] itasegm1\[755\]
+ itasegm1\[743\] itasegm1\[744\] itasegm1\[745\] itasegm1\[746\] itasegm1\[747\]
+ itasegm1\[748\] itasegm1\[749\] itasegm1\[750\] itasegm1\[751\] itasel1\[636\] itasel1\[646\]
+ itasel1\[647\] itasel1\[637\] itasel1\[638\] itasel1\[639\] itasel1\[640\] itasel1\[641\]
+ itasel1\[642\] itasel1\[643\] itasel1\[644\] itasel1\[645\] vdd vss ita54
Xita21 wb_clk_i itasegm1\[280\] itasegm1\[290\] itasegm1\[291\] itasegm1\[292\] itasegm1\[293\]
+ itasegm1\[281\] itasegm1\[282\] itasegm1\[283\] itasegm1\[284\] itasegm1\[285\]
+ itasegm1\[286\] itasegm1\[287\] itasegm1\[288\] itasegm1\[289\] itasel1\[240\] itasel1\[250\]
+ itasel1\[251\] itasel1\[241\] itasel1\[242\] itasel1\[243\] itasel1\[244\] itasel1\[245\]
+ itasel1\[246\] itasel1\[247\] itasel1\[248\] itasel1\[249\] vdd vss ita21
Xita43 wb_clk_i itasegm1\[588\] itasegm1\[598\] itasegm1\[599\] itasegm1\[600\] itasegm1\[601\]
+ itasegm1\[589\] itasegm1\[590\] itasegm1\[591\] itasegm1\[592\] itasegm1\[593\]
+ itasegm1\[594\] itasegm1\[595\] itasegm1\[596\] itasegm1\[597\] itasel1\[504\] itasel1\[514\]
+ itasel1\[515\] itasel1\[505\] itasel1\[506\] itasel1\[507\] itasel1\[508\] itasel1\[509\]
+ itasel1\[510\] itasel1\[511\] itasel1\[512\] itasel1\[513\] vdd vss ita43
Xita10 wb_clk_i itasegm1\[126\] itasegm1\[136\] itasegm1\[137\] itasegm1\[138\] itasegm1\[139\]
+ itasegm1\[127\] itasegm1\[128\] itasegm1\[129\] itasegm1\[130\] itasegm1\[131\]
+ itasegm1\[132\] itasegm1\[133\] itasegm1\[134\] itasegm1\[135\] itasel1\[108\] itasel1\[118\]
+ itasel1\[119\] itasel1\[109\] itasel1\[110\] itasel1\[111\] itasel1\[112\] itasel1\[113\]
+ itasel1\[114\] itasel1\[115\] itasel1\[116\] itasel1\[117\] vdd vss ita10
Xita8 wb_clk_i itasegm1\[98\] itasegm1\[108\] itasegm1\[109\] itasegm1\[110\] itasegm1\[111\]
+ itasegm1\[99\] itasegm1\[100\] itasegm1\[101\] itasegm1\[102\] itasegm1\[103\] itasegm1\[104\]
+ itasegm1\[105\] itasegm1\[106\] itasegm1\[107\] itasel1\[84\] itasel1\[94\] itasel1\[95\]
+ itasel1\[85\] itasel1\[86\] itasel1\[87\] itasel1\[88\] itasel1\[89\] itasel1\[90\]
+ itasel1\[91\] itasel1\[92\] itasel1\[93\] vdd vss ita8
Xita55 wb_clk_i itasegm1\[756\] itasegm1\[766\] itasegm1\[767\] itasegm1\[768\] itasegm1\[769\]
+ itasegm1\[757\] itasegm1\[758\] itasegm1\[759\] itasegm1\[760\] itasegm1\[761\]
+ itasegm1\[762\] itasegm1\[763\] itasegm1\[764\] itasegm1\[765\] itasel1\[648\] itasel1\[658\]
+ itasel1\[659\] itasel1\[649\] itasel1\[650\] itasel1\[651\] itasel1\[652\] itasel1\[653\]
+ itasel1\[654\] itasel1\[655\] itasel1\[656\] itasel1\[657\] vdd vss ita55
Xita22 wb_clk_i itasegm1\[294\] itasegm1\[304\] itasegm1\[305\] itasegm1\[306\] itasegm1\[307\]
+ itasegm1\[295\] itasegm1\[296\] itasegm1\[297\] itasegm1\[298\] itasegm1\[299\]
+ itasegm1\[300\] itasegm1\[301\] itasegm1\[302\] itasegm1\[303\] itasel1\[252\] itasel1\[262\]
+ itasel1\[263\] itasel1\[253\] itasel1\[254\] itasel1\[255\] itasel1\[256\] itasel1\[257\]
+ itasel1\[258\] itasel1\[259\] itasel1\[260\] itasel1\[261\] vdd vss ita22
Xita44 wb_clk_i itasegm1\[602\] itasegm1\[612\] itasegm1\[613\] itasegm1\[614\] itasegm1\[615\]
+ itasegm1\[603\] itasegm1\[604\] itasegm1\[605\] itasegm1\[606\] itasegm1\[607\]
+ itasegm1\[608\] itasegm1\[609\] itasegm1\[610\] itasegm1\[611\] itasel1\[516\] itasel1\[526\]
+ itasel1\[527\] itasel1\[517\] itasel1\[518\] itasel1\[519\] itasel1\[520\] itasel1\[521\]
+ itasel1\[522\] itasel1\[523\] itasel1\[524\] itasel1\[525\] vdd vss ita44
Xita11 wb_clk_i itasegm1\[140\] itasegm1\[150\] itasegm1\[151\] itasegm1\[152\] itasegm1\[153\]
+ itasegm1\[141\] itasegm1\[142\] itasegm1\[143\] itasegm1\[144\] itasegm1\[145\]
+ itasegm1\[146\] itasegm1\[147\] itasegm1\[148\] itasegm1\[149\] itasel1\[120\] itasel1\[130\]
+ itasel1\[131\] itasel1\[121\] itasel1\[122\] itasel1\[123\] itasel1\[124\] itasel1\[125\]
+ itasel1\[126\] itasel1\[127\] itasel1\[128\] itasel1\[129\] vdd vss ita11
Xita33 wb_clk_i itasegm1\[448\] itasegm1\[458\] itasegm1\[459\] itasegm1\[460\] itasegm1\[461\]
+ itasegm1\[449\] itasegm1\[450\] itasegm1\[451\] itasegm1\[452\] itasegm1\[453\]
+ itasegm1\[454\] itasegm1\[455\] itasegm1\[456\] itasegm1\[457\] itasel1\[384\] itasel1\[394\]
+ itasel1\[395\] itasel1\[385\] itasel1\[386\] itasel1\[387\] itasel1\[388\] itasel1\[389\]
+ itasel1\[390\] itasel1\[391\] itasel1\[392\] itasel1\[393\] vdd vss ita33
Xita56 wb_clk_i itasegm1\[770\] itasegm1\[780\] itasegm1\[781\] itasegm1\[782\] itasegm1\[783\]
+ itasegm1\[771\] itasegm1\[772\] itasegm1\[773\] itasegm1\[774\] itasegm1\[775\]
+ itasegm1\[776\] itasegm1\[777\] itasegm1\[778\] itasegm1\[779\] itasel1\[660\] itasel1\[670\]
+ itasel1\[671\] itasel1\[661\] itasel1\[662\] itasel1\[663\] itasel1\[664\] itasel1\[665\]
+ itasel1\[666\] itasel1\[667\] itasel1\[668\] itasel1\[669\] vdd vss ita56
Xita23 wb_clk_i itasegm1\[308\] itasegm1\[318\] itasegm1\[319\] itasegm1\[320\] itasegm1\[321\]
+ itasegm1\[309\] itasegm1\[310\] itasegm1\[311\] itasegm1\[312\] itasegm1\[313\]
+ itasegm1\[314\] itasegm1\[315\] itasegm1\[316\] itasegm1\[317\] itasel1\[264\] itasel1\[274\]
+ itasel1\[275\] itasel1\[265\] itasel1\[266\] itasel1\[267\] itasel1\[268\] itasel1\[269\]
+ itasel1\[270\] itasel1\[271\] itasel1\[272\] itasel1\[273\] vdd vss ita23
Xita45 wb_clk_i itasegm1\[616\] itasegm1\[626\] itasegm1\[627\] itasegm1\[628\] itasegm1\[629\]
+ itasegm1\[617\] itasegm1\[618\] itasegm1\[619\] itasegm1\[620\] itasegm1\[621\]
+ itasegm1\[622\] itasegm1\[623\] itasegm1\[624\] itasegm1\[625\] itasel1\[528\] itasel1\[538\]
+ itasel1\[539\] itasel1\[529\] itasel1\[530\] itasel1\[531\] itasel1\[532\] itasel1\[533\]
+ itasel1\[534\] itasel1\[535\] itasel1\[536\] itasel1\[537\] vdd vss ita45
Xita12 wb_clk_i itasegm1\[154\] itasegm1\[164\] itasegm1\[165\] itasegm1\[166\] itasegm1\[167\]
+ itasegm1\[155\] itasegm1\[156\] itasegm1\[157\] itasegm1\[158\] itasegm1\[159\]
+ itasegm1\[160\] itasegm1\[161\] itasegm1\[162\] itasegm1\[163\] itasel1\[132\] itasel1\[142\]
+ itasel1\[143\] itasel1\[133\] itasel1\[134\] itasel1\[135\] itasel1\[136\] itasel1\[137\]
+ itasel1\[138\] itasel1\[139\] itasel1\[140\] itasel1\[141\] vdd vss ita12
Xita34 wb_clk_i itasegm1\[462\] itasegm1\[472\] itasegm1\[473\] itasegm1\[474\] itasegm1\[475\]
+ itasegm1\[463\] itasegm1\[464\] itasegm1\[465\] itasegm1\[466\] itasegm1\[467\]
+ itasegm1\[468\] itasegm1\[469\] itasegm1\[470\] itasegm1\[471\] itasel1\[396\] itasel1\[406\]
+ itasel1\[407\] itasel1\[397\] itasel1\[398\] itasel1\[399\] itasel1\[400\] itasel1\[401\]
+ itasel1\[402\] itasel1\[403\] itasel1\[404\] itasel1\[405\] vdd vss ita34
Xita9 wb_clk_i itasegm1\[112\] itasegm1\[122\] itasegm1\[123\] itasegm1\[124\] itasegm1\[125\]
+ itasegm1\[113\] itasegm1\[114\] itasegm1\[115\] itasegm1\[116\] itasegm1\[117\]
+ itasegm1\[118\] itasegm1\[119\] itasegm1\[120\] itasegm1\[121\] itasel1\[96\] itasel1\[106\]
+ itasel1\[107\] itasel1\[97\] itasel1\[98\] itasel1\[99\] itasel1\[100\] itasel1\[101\]
+ itasel1\[102\] itasel1\[103\] itasel1\[104\] itasel1\[105\] vdd vss ita9
Xita24 wb_clk_i itasegm1\[322\] itasegm1\[332\] itasegm1\[333\] itasegm1\[334\] itasegm1\[335\]
+ itasegm1\[323\] itasegm1\[324\] itasegm1\[325\] itasegm1\[326\] itasegm1\[327\]
+ itasegm1\[328\] itasegm1\[329\] itasegm1\[330\] itasegm1\[331\] itasel1\[276\] itasel1\[286\]
+ itasel1\[287\] itasel1\[277\] itasel1\[278\] itasel1\[279\] itasel1\[280\] itasel1\[281\]
+ itasel1\[282\] itasel1\[283\] itasel1\[284\] itasel1\[285\] vdd vss ita24
Xita47 wb_clk_i itasegm1\[644\] itasegm1\[654\] itasegm1\[655\] itasegm1\[656\] itasegm1\[657\]
+ itasegm1\[645\] itasegm1\[646\] itasegm1\[647\] itasegm1\[648\] itasegm1\[649\]
+ itasegm1\[650\] itasegm1\[651\] itasegm1\[652\] itasegm1\[653\] itasel1\[552\] itasel1\[562\]
+ itasel1\[563\] itasel1\[553\] itasel1\[554\] itasel1\[555\] itasel1\[556\] itasel1\[557\]
+ itasel1\[558\] itasel1\[559\] itasel1\[560\] itasel1\[561\] vdd vss ita47
Xita46 wb_clk_i itasegm1\[630\] itasegm1\[640\] itasegm1\[641\] itasegm1\[642\] itasegm1\[643\]
+ itasegm1\[631\] itasegm1\[632\] itasegm1\[633\] itasegm1\[634\] itasegm1\[635\]
+ itasegm1\[636\] itasegm1\[637\] itasegm1\[638\] itasegm1\[639\] itasel1\[540\] itasel1\[550\]
+ itasel1\[551\] itasel1\[541\] itasel1\[542\] itasel1\[543\] itasel1\[544\] itasel1\[545\]
+ itasel1\[546\] itasel1\[547\] itasel1\[548\] itasel1\[549\] vdd vss ita46
Xita14 wb_clk_i itasegm1\[182\] itasegm1\[192\] itasegm1\[193\] itasegm1\[194\] itasegm1\[195\]
+ itasegm1\[183\] itasegm1\[184\] itasegm1\[185\] itasegm1\[186\] itasegm1\[187\]
+ itasegm1\[188\] itasegm1\[189\] itasegm1\[190\] itasegm1\[191\] itasel1\[156\] itasel1\[166\]
+ itasel1\[167\] itasel1\[157\] itasel1\[158\] itasel1\[159\] itasel1\[160\] itasel1\[161\]
+ itasel1\[162\] itasel1\[163\] itasel1\[164\] itasel1\[165\] vdd vss ita14
Xita13 wb_clk_i itasegm1\[168\] itasegm1\[178\] itasegm1\[179\] itasegm1\[180\] itasegm1\[181\]
+ itasegm1\[169\] itasegm1\[170\] itasegm1\[171\] itasegm1\[172\] itasegm1\[173\]
+ itasegm1\[174\] itasegm1\[175\] itasegm1\[176\] itasegm1\[177\] itasel1\[144\] itasel1\[154\]
+ itasel1\[155\] itasel1\[145\] itasel1\[146\] itasel1\[147\] itasel1\[148\] itasel1\[149\]
+ itasel1\[150\] itasel1\[151\] itasel1\[152\] itasel1\[153\] vdd vss ita13
Xita36 wb_clk_i itasegm1\[490\] itasegm1\[500\] itasegm1\[501\] itasegm1\[502\] itasegm1\[503\]
+ itasegm1\[491\] itasegm1\[492\] itasegm1\[493\] itasegm1\[494\] itasegm1\[495\]
+ itasegm1\[496\] itasegm1\[497\] itasegm1\[498\] itasegm1\[499\] itasel1\[420\] itasel1\[430\]
+ itasel1\[431\] itasel1\[421\] itasel1\[422\] itasel1\[423\] itasel1\[424\] itasel1\[425\]
+ itasel1\[426\] itasel1\[427\] itasel1\[428\] itasel1\[429\] vdd vss ita36
Xita35 wb_clk_i itasegm1\[476\] itasegm1\[486\] itasegm1\[487\] itasegm1\[488\] itasegm1\[489\]
+ itasegm1\[477\] itasegm1\[478\] itasegm1\[479\] itasegm1\[480\] itasegm1\[481\]
+ itasegm1\[482\] itasegm1\[483\] itasegm1\[484\] itasegm1\[485\] itasel1\[408\] itasel1\[418\]
+ itasel1\[419\] itasel1\[409\] itasel1\[410\] itasel1\[411\] itasel1\[412\] itasel1\[413\]
+ itasel1\[414\] itasel1\[415\] itasel1\[416\] itasel1\[417\] vdd vss ita35
Xita57 wb_clk_i itasegm1\[784\] itasegm1\[794\] itasegm1\[795\] itasegm1\[796\] itasegm1\[797\]
+ itasegm1\[785\] itasegm1\[786\] itasegm1\[787\] itasegm1\[788\] itasegm1\[789\]
+ itasegm1\[790\] itasegm1\[791\] itasegm1\[792\] itasegm1\[793\] itasel1\[672\] itasel1\[682\]
+ itasel1\[683\] itasel1\[673\] itasel1\[674\] itasel1\[675\] itasel1\[676\] itasel1\[677\]
+ itasel1\[678\] itasel1\[679\] itasel1\[680\] itasel1\[681\] vdd vss ita57
Xita58 wb_clk_i itasegm1\[798\] itasegm1\[808\] itasegm1\[809\] itasegm1\[810\] itasegm1\[811\]
+ itasegm1\[799\] itasegm1\[800\] itasegm1\[801\] itasegm1\[802\] itasegm1\[803\]
+ itasegm1\[804\] itasegm1\[805\] itasegm1\[806\] itasegm1\[807\] itasel1\[684\] itasel1\[694\]
+ itasel1\[695\] itasel1\[685\] itasel1\[686\] itasel1\[687\] itasel1\[688\] itasel1\[689\]
+ itasel1\[690\] itasel1\[691\] itasel1\[692\] itasel1\[693\] vdd vss ita58
Xita25 wb_clk_i itasegm1\[336\] itasegm1\[346\] itasegm1\[347\] itasegm1\[348\] itasegm1\[349\]
+ itasegm1\[337\] itasegm1\[338\] itasegm1\[339\] itasegm1\[340\] itasegm1\[341\]
+ itasegm1\[342\] itasegm1\[343\] itasegm1\[344\] itasegm1\[345\] itasel1\[288\] itasel1\[298\]
+ itasel1\[299\] itasel1\[289\] itasel1\[290\] itasel1\[291\] itasel1\[292\] itasel1\[293\]
+ itasel1\[294\] itasel1\[295\] itasel1\[296\] itasel1\[297\] vdd vss ita25
Xita48 wb_clk_i itasegm1\[658\] itasegm1\[668\] itasegm1\[669\] itasegm1\[670\] itasegm1\[671\]
+ itasegm1\[659\] itasegm1\[660\] itasegm1\[661\] itasegm1\[662\] itasegm1\[663\]
+ itasegm1\[664\] itasegm1\[665\] itasegm1\[666\] itasegm1\[667\] itasel1\[564\] itasel1\[574\]
+ itasel1\[575\] itasel1\[565\] itasel1\[566\] itasel1\[567\] itasel1\[568\] itasel1\[569\]
+ itasel1\[570\] itasel1\[571\] itasel1\[572\] itasel1\[573\] vdd vss ita48
Xita15 wb_clk_i itasegm1\[196\] itasegm1\[206\] itasegm1\[207\] itasegm1\[208\] itasegm1\[209\]
+ itasegm1\[197\] itasegm1\[198\] itasegm1\[199\] itasegm1\[200\] itasegm1\[201\]
+ itasegm1\[202\] itasegm1\[203\] itasegm1\[204\] itasegm1\[205\] itasel1\[168\] itasel1\[178\]
+ itasel1\[179\] itasel1\[169\] itasel1\[170\] itasel1\[171\] itasel1\[172\] itasel1\[173\]
+ itasel1\[174\] itasel1\[175\] itasel1\[176\] itasel1\[177\] vdd vss ita15
Xita37 wb_clk_i itasegm1\[504\] itasegm1\[514\] itasegm1\[515\] itasegm1\[516\] itasegm1\[517\]
+ itasegm1\[505\] itasegm1\[506\] itasegm1\[507\] itasegm1\[508\] itasegm1\[509\]
+ itasegm1\[510\] itasegm1\[511\] itasegm1\[512\] itasegm1\[513\] itasel1\[432\] itasel1\[442\]
+ itasel1\[443\] itasel1\[433\] itasel1\[434\] itasel1\[435\] itasel1\[436\] itasel1\[437\]
+ itasel1\[438\] itasel1\[439\] itasel1\[440\] itasel1\[441\] vdd vss ita37
Xita59 wb_clk_i itasegm1\[812\] itasegm1\[822\] itasegm1\[823\] itasegm1\[824\] itasegm1\[825\]
+ itasegm1\[813\] itasegm1\[814\] itasegm1\[815\] itasegm1\[816\] itasegm1\[817\]
+ itasegm1\[818\] itasegm1\[819\] itasegm1\[820\] itasegm1\[821\] itasel1\[696\] itasel1\[706\]
+ itasel1\[707\] itasel1\[697\] itasel1\[698\] itasel1\[699\] itasel1\[700\] itasel1\[701\]
+ itasel1\[702\] itasel1\[703\] itasel1\[704\] itasel1\[705\] vdd vss ita59
Xita26 wb_clk_i itasegm1\[350\] itasegm1\[360\] itasegm1\[361\] itasegm1\[362\] itasegm1\[363\]
+ itasegm1\[351\] itasegm1\[352\] itasegm1\[353\] itasegm1\[354\] itasegm1\[355\]
+ itasegm1\[356\] itasegm1\[357\] itasegm1\[358\] itasegm1\[359\] itasel1\[300\] itasel1\[310\]
+ itasel1\[311\] itasel1\[301\] itasel1\[302\] itasel1\[303\] itasel1\[304\] itasel1\[305\]
+ itasel1\[306\] itasel1\[307\] itasel1\[308\] itasel1\[309\] vdd vss ita26
Xita16 wb_clk_i itasegm1\[210\] itasegm1\[220\] itasegm1\[221\] itasegm1\[222\] itasegm1\[223\]
+ itasegm1\[211\] itasegm1\[212\] itasegm1\[213\] itasegm1\[214\] itasegm1\[215\]
+ itasegm1\[216\] itasegm1\[217\] itasegm1\[218\] itasegm1\[219\] itasel1\[180\] itasel1\[190\]
+ itasel1\[191\] itasel1\[181\] itasel1\[182\] itasel1\[183\] itasel1\[184\] itasel1\[185\]
+ itasel1\[186\] itasel1\[187\] itasel1\[188\] itasel1\[189\] vdd vss ita16
Xita38 wb_clk_i itasegm1\[518\] itasegm1\[528\] itasegm1\[529\] itasegm1\[530\] itasegm1\[531\]
+ itasegm1\[519\] itasegm1\[520\] itasegm1\[521\] itasegm1\[522\] itasegm1\[523\]
+ itasegm1\[524\] itasegm1\[525\] itasegm1\[526\] itasegm1\[527\] itasel1\[444\] itasel1\[454\]
+ itasel1\[455\] itasel1\[445\] itasel1\[446\] itasel1\[447\] itasel1\[448\] itasel1\[449\]
+ itasel1\[450\] itasel1\[451\] itasel1\[452\] itasel1\[453\] vdd vss ita38
Xita27 wb_clk_i itasegm1\[364\] itasegm1\[374\] itasegm1\[375\] itasegm1\[376\] itasegm1\[377\]
+ itasegm1\[365\] itasegm1\[366\] itasegm1\[367\] itasegm1\[368\] itasegm1\[369\]
+ itasegm1\[370\] itasegm1\[371\] itasegm1\[372\] itasegm1\[373\] itasel1\[312\] itasel1\[322\]
+ itasel1\[323\] itasel1\[313\] itasel1\[314\] itasel1\[315\] itasel1\[316\] itasel1\[317\]
+ itasel1\[318\] itasel1\[319\] itasel1\[320\] itasel1\[321\] vdd vss ita27
Xita49 wb_clk_i itasegm1\[672\] itasegm1\[682\] itasegm1\[683\] itasegm1\[684\] itasegm1\[685\]
+ itasegm1\[673\] itasegm1\[674\] itasegm1\[675\] itasegm1\[676\] itasegm1\[677\]
+ itasegm1\[678\] itasegm1\[679\] itasegm1\[680\] itasegm1\[681\] itasel1\[576\] itasel1\[586\]
+ itasel1\[587\] itasel1\[577\] itasel1\[578\] itasel1\[579\] itasel1\[580\] itasel1\[581\]
+ itasel1\[582\] itasel1\[583\] itasel1\[584\] itasel1\[585\] vdd vss ita49
Xita39 wb_clk_i itasegm1\[532\] itasegm1\[542\] itasegm1\[543\] itasegm1\[544\] itasegm1\[545\]
+ itasegm1\[533\] itasegm1\[534\] itasegm1\[535\] itasegm1\[536\] itasegm1\[537\]
+ itasegm1\[538\] itasegm1\[539\] itasegm1\[540\] itasegm1\[541\] itasel1\[456\] itasel1\[466\]
+ itasel1\[467\] itasel1\[457\] itasel1\[458\] itasel1\[459\] itasel1\[460\] itasel1\[461\]
+ itasel1\[462\] itasel1\[463\] itasel1\[464\] itasel1\[465\] vdd vss ita39
Xita28 wb_clk_i itasegm1\[378\] itasegm1\[388\] itasegm1\[389\] itasegm1\[390\] itasegm1\[391\]
+ itasegm1\[379\] itasegm1\[380\] itasegm1\[381\] itasegm1\[382\] itasegm1\[383\]
+ itasegm1\[384\] itasegm1\[385\] itasegm1\[386\] itasegm1\[387\] itasel1\[324\] itasel1\[334\]
+ itasel1\[335\] itasel1\[325\] itasel1\[326\] itasel1\[327\] itasel1\[328\] itasel1\[329\]
+ itasel1\[330\] itasel1\[331\] itasel1\[332\] itasel1\[333\] vdd vss ita28
Xita17 wb_clk_i itasegm1\[224\] itasegm1\[234\] itasegm1\[235\] itasegm1\[236\] itasegm1\[237\]
+ itasegm1\[225\] itasegm1\[226\] itasegm1\[227\] itasegm1\[228\] itasegm1\[229\]
+ itasegm1\[230\] itasegm1\[231\] itasegm1\[232\] itasegm1\[233\] itasel1\[192\] itasel1\[202\]
+ itasel1\[203\] itasel1\[193\] itasel1\[194\] itasel1\[195\] itasel1\[196\] itasel1\[197\]
+ itasel1\[198\] itasel1\[199\] itasel1\[200\] itasel1\[201\] vdd vss ita17
Xita29 wb_clk_i itasegm1\[392\] itasegm1\[402\] itasegm1\[403\] itasegm1\[404\] itasegm1\[405\]
+ itasegm1\[393\] itasegm1\[394\] itasegm1\[395\] itasegm1\[396\] itasegm1\[397\]
+ itasegm1\[398\] itasegm1\[399\] itasegm1\[400\] itasegm1\[401\] itasel1\[336\] itasel1\[346\]
+ itasel1\[347\] itasel1\[337\] itasel1\[338\] itasel1\[339\] itasel1\[340\] itasel1\[341\]
+ itasel1\[342\] itasel1\[343\] itasel1\[344\] itasel1\[345\] vdd vss ita29
Xita18 wb_clk_i itasegm1\[238\] itasegm1\[248\] itasegm1\[249\] itasegm1\[250\] itasegm1\[251\]
+ itasegm1\[239\] itasegm1\[240\] itasegm1\[241\] itasegm1\[242\] itasegm1\[243\]
+ itasegm1\[244\] itasegm1\[245\] itasegm1\[246\] itasegm1\[247\] itasel1\[204\] itasel1\[214\]
+ itasel1\[215\] itasel1\[205\] itasel1\[206\] itasel1\[207\] itasel1\[208\] itasel1\[209\]
+ itasel1\[210\] itasel1\[211\] itasel1\[212\] itasel1\[213\] vdd vss ita18
Xita19 wb_clk_i itasegm1\[252\] itasegm1\[262\] itasegm1\[263\] itasegm1\[264\] itasegm1\[265\]
+ itasegm1\[253\] itasegm1\[254\] itasegm1\[255\] itasegm1\[256\] itasegm1\[257\]
+ itasegm1\[258\] itasegm1\[259\] itasegm1\[260\] itasegm1\[261\] itasel1\[216\] itasel1\[226\]
+ itasel1\[227\] itasel1\[217\] itasel1\[218\] itasel1\[219\] itasel1\[220\] itasel1\[221\]
+ itasel1\[222\] itasel1\[223\] itasel1\[224\] itasel1\[225\] vdd vss ita19
.ends

