magic
tech gf180mcuD
magscale 1 10
timestamp 1699641497
<< metal1 >>
rect 1344 38442 40656 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 40656 38442
rect 1344 38356 40656 38390
rect 22430 38274 22482 38286
rect 22430 38210 22482 38222
rect 25566 38274 25618 38286
rect 25566 38210 25618 38222
rect 18834 38110 18846 38162
rect 18898 38110 18910 38162
rect 19730 37998 19742 38050
rect 19794 37998 19806 38050
rect 21410 37998 21422 38050
rect 21474 37998 21486 38050
rect 24546 37998 24558 38050
rect 24610 37998 24622 38050
rect 27470 37938 27522 37950
rect 27470 37874 27522 37886
rect 1344 37658 40656 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 40656 37658
rect 1344 37572 40656 37606
rect 18398 37490 18450 37502
rect 18398 37426 18450 37438
rect 20750 37490 20802 37502
rect 20750 37426 20802 37438
rect 19730 37214 19742 37266
rect 19794 37214 19806 37266
rect 1344 36874 40656 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 40656 36874
rect 1344 36788 40656 36822
rect 18734 36706 18786 36718
rect 18734 36642 18786 36654
rect 24782 36706 24834 36718
rect 24782 36642 24834 36654
rect 17714 36430 17726 36482
rect 17778 36430 17790 36482
rect 24098 36430 24110 36482
rect 24162 36430 24174 36482
rect 1710 36370 1762 36382
rect 1710 36306 1762 36318
rect 1344 36090 40656 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 40656 36090
rect 1344 36004 40656 36038
rect 1344 35306 40656 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 40656 35306
rect 1344 35220 40656 35254
rect 1344 34522 40656 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 40656 34522
rect 1344 34436 40656 34470
rect 1344 33738 40656 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 40656 33738
rect 1344 33652 40656 33686
rect 1344 32954 40656 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 40656 32954
rect 1344 32868 40656 32902
rect 1344 32170 40656 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 40656 32170
rect 1344 32084 40656 32118
rect 1344 31386 40656 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 40656 31386
rect 1344 31300 40656 31334
rect 1344 30602 40656 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 40656 30602
rect 1344 30516 40656 30550
rect 1344 29818 40656 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 40656 29818
rect 1344 29732 40656 29766
rect 1344 29034 40656 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 40656 29034
rect 1344 28948 40656 28982
rect 18622 28642 18674 28654
rect 18622 28578 18674 28590
rect 18174 28530 18226 28542
rect 18174 28466 18226 28478
rect 18846 28530 18898 28542
rect 18846 28466 18898 28478
rect 18958 28530 19010 28542
rect 18958 28466 19010 28478
rect 19406 28530 19458 28542
rect 19406 28466 19458 28478
rect 19518 28530 19570 28542
rect 19518 28466 19570 28478
rect 17838 28418 17890 28430
rect 17838 28354 17890 28366
rect 18062 28418 18114 28430
rect 18062 28354 18114 28366
rect 19742 28418 19794 28430
rect 19742 28354 19794 28366
rect 1344 28250 40656 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 40656 28250
rect 1344 28164 40656 28198
rect 24098 28030 24110 28082
rect 24162 28030 24174 28082
rect 24446 27858 24498 27870
rect 15026 27806 15038 27858
rect 15090 27806 15102 27858
rect 17490 27806 17502 27858
rect 17554 27806 17566 27858
rect 20962 27806 20974 27858
rect 21026 27806 21038 27858
rect 24446 27794 24498 27806
rect 15598 27746 15650 27758
rect 12114 27694 12126 27746
rect 12178 27694 12190 27746
rect 14242 27694 14254 27746
rect 14306 27694 14318 27746
rect 18162 27694 18174 27746
rect 18226 27694 18238 27746
rect 20290 27694 20302 27746
rect 20354 27694 20366 27746
rect 21634 27694 21646 27746
rect 21698 27694 21710 27746
rect 23762 27694 23774 27746
rect 23826 27694 23838 27746
rect 15598 27682 15650 27694
rect 1344 27466 40656 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 40656 27466
rect 1344 27380 40656 27414
rect 14142 27298 14194 27310
rect 14142 27234 14194 27246
rect 1934 27186 1986 27198
rect 21646 27186 21698 27198
rect 17154 27134 17166 27186
rect 17218 27134 17230 27186
rect 19282 27134 19294 27186
rect 19346 27134 19358 27186
rect 1934 27122 1986 27134
rect 21646 27122 21698 27134
rect 22542 27186 22594 27198
rect 22542 27122 22594 27134
rect 19518 27074 19570 27086
rect 4274 27022 4286 27074
rect 4338 27022 4350 27074
rect 16482 27022 16494 27074
rect 16546 27022 16558 27074
rect 19518 27010 19570 27022
rect 19854 27074 19906 27086
rect 19854 27010 19906 27022
rect 21422 27074 21474 27086
rect 21970 27022 21982 27074
rect 22034 27022 22046 27074
rect 21422 27010 21474 27022
rect 14142 26962 14194 26974
rect 14142 26898 14194 26910
rect 14254 26962 14306 26974
rect 14254 26898 14306 26910
rect 21758 26962 21810 26974
rect 21758 26898 21810 26910
rect 22430 26962 22482 26974
rect 22430 26898 22482 26910
rect 19742 26850 19794 26862
rect 19742 26786 19794 26798
rect 20526 26850 20578 26862
rect 20526 26786 20578 26798
rect 21534 26850 21586 26862
rect 21534 26786 21586 26798
rect 23998 26850 24050 26862
rect 23998 26786 24050 26798
rect 1344 26682 40656 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 40656 26682
rect 1344 26596 40656 26630
rect 23550 26402 23602 26414
rect 23550 26338 23602 26350
rect 13906 26238 13918 26290
rect 13970 26238 13982 26290
rect 22978 26238 22990 26290
rect 23042 26238 23054 26290
rect 17502 26178 17554 26190
rect 14690 26126 14702 26178
rect 14754 26126 14766 26178
rect 16818 26126 16830 26178
rect 16882 26126 16894 26178
rect 17502 26114 17554 26126
rect 19518 26178 19570 26190
rect 20178 26126 20190 26178
rect 20242 26126 20254 26178
rect 22306 26126 22318 26178
rect 22370 26126 22382 26178
rect 19518 26114 19570 26126
rect 1344 25898 40656 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 40656 25898
rect 1344 25812 40656 25846
rect 15710 25730 15762 25742
rect 15710 25666 15762 25678
rect 1934 25618 1986 25630
rect 22430 25618 22482 25630
rect 16930 25566 16942 25618
rect 16994 25566 17006 25618
rect 21858 25566 21870 25618
rect 21922 25566 21934 25618
rect 1934 25554 1986 25566
rect 22430 25554 22482 25566
rect 14254 25506 14306 25518
rect 4274 25454 4286 25506
rect 4338 25454 4350 25506
rect 14254 25442 14306 25454
rect 15822 25506 15874 25518
rect 17054 25506 17106 25518
rect 16818 25454 16830 25506
rect 16882 25454 16894 25506
rect 15822 25442 15874 25454
rect 17054 25442 17106 25454
rect 12798 25394 12850 25406
rect 12798 25330 12850 25342
rect 13582 25394 13634 25406
rect 13582 25330 13634 25342
rect 13694 25394 13746 25406
rect 13694 25330 13746 25342
rect 14478 25394 14530 25406
rect 14478 25330 14530 25342
rect 14590 25394 14642 25406
rect 17502 25394 17554 25406
rect 21310 25394 21362 25406
rect 16146 25342 16158 25394
rect 16210 25342 16222 25394
rect 18610 25342 18622 25394
rect 18674 25342 18686 25394
rect 14590 25330 14642 25342
rect 17502 25330 17554 25342
rect 21310 25330 21362 25342
rect 21870 25394 21922 25406
rect 21870 25330 21922 25342
rect 12462 25282 12514 25294
rect 12462 25218 12514 25230
rect 12686 25282 12738 25294
rect 12686 25218 12738 25230
rect 13358 25282 13410 25294
rect 13358 25218 13410 25230
rect 16494 25282 16546 25294
rect 16494 25218 16546 25230
rect 17278 25282 17330 25294
rect 17278 25218 17330 25230
rect 18286 25282 18338 25294
rect 18286 25218 18338 25230
rect 21534 25282 21586 25294
rect 21534 25218 21586 25230
rect 21758 25282 21810 25294
rect 21758 25218 21810 25230
rect 22318 25282 22370 25294
rect 22318 25218 22370 25230
rect 1344 25114 40656 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 40656 25114
rect 1344 25028 40656 25062
rect 13918 24946 13970 24958
rect 13918 24882 13970 24894
rect 20190 24946 20242 24958
rect 20190 24882 20242 24894
rect 19966 24834 20018 24846
rect 19966 24770 20018 24782
rect 24110 24834 24162 24846
rect 24110 24770 24162 24782
rect 19854 24722 19906 24734
rect 4274 24670 4286 24722
rect 4338 24670 4350 24722
rect 13458 24670 13470 24722
rect 13522 24670 13534 24722
rect 19854 24658 19906 24670
rect 23998 24722 24050 24734
rect 37650 24670 37662 24722
rect 37714 24670 37726 24722
rect 23998 24658 24050 24670
rect 10546 24558 10558 24610
rect 10610 24558 10622 24610
rect 12674 24558 12686 24610
rect 12738 24558 12750 24610
rect 1934 24498 1986 24510
rect 1934 24434 1986 24446
rect 24110 24498 24162 24510
rect 24110 24434 24162 24446
rect 40014 24498 40066 24510
rect 40014 24434 40066 24446
rect 1344 24330 40656 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 40656 24330
rect 1344 24244 40656 24278
rect 1934 24050 1986 24062
rect 13582 24050 13634 24062
rect 40014 24050 40066 24062
rect 9986 23998 9998 24050
rect 10050 23998 10062 24050
rect 12114 23998 12126 24050
rect 12178 23998 12190 24050
rect 20738 23998 20750 24050
rect 20802 23998 20814 24050
rect 25666 23998 25678 24050
rect 25730 23998 25742 24050
rect 1934 23986 1986 23998
rect 13582 23986 13634 23998
rect 40014 23986 40066 23998
rect 13470 23938 13522 23950
rect 4274 23886 4286 23938
rect 4338 23886 4350 23938
rect 12898 23886 12910 23938
rect 12962 23886 12974 23938
rect 13470 23874 13522 23886
rect 13694 23938 13746 23950
rect 13694 23874 13746 23886
rect 17838 23938 17890 23950
rect 18498 23886 18510 23938
rect 18562 23886 18574 23938
rect 19618 23886 19630 23938
rect 19682 23886 19694 23938
rect 20290 23886 20302 23938
rect 20354 23886 20366 23938
rect 22866 23886 22878 23938
rect 22930 23886 22942 23938
rect 37650 23886 37662 23938
rect 37714 23886 37726 23938
rect 17838 23874 17890 23886
rect 14030 23826 14082 23838
rect 18162 23774 18174 23826
rect 18226 23774 18238 23826
rect 19954 23774 19966 23826
rect 20018 23774 20030 23826
rect 20626 23774 20638 23826
rect 20690 23774 20702 23826
rect 23538 23774 23550 23826
rect 23602 23774 23614 23826
rect 14030 23762 14082 23774
rect 26126 23714 26178 23726
rect 26126 23650 26178 23662
rect 28366 23714 28418 23726
rect 28366 23650 28418 23662
rect 1344 23546 40656 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 40656 23546
rect 1344 23460 40656 23494
rect 12462 23378 12514 23390
rect 12462 23314 12514 23326
rect 12686 23378 12738 23390
rect 19518 23378 19570 23390
rect 17714 23326 17726 23378
rect 17778 23326 17790 23378
rect 12686 23314 12738 23326
rect 19518 23314 19570 23326
rect 20414 23378 20466 23390
rect 20414 23314 20466 23326
rect 21646 23378 21698 23390
rect 21646 23314 21698 23326
rect 23662 23378 23714 23390
rect 23662 23314 23714 23326
rect 17390 23266 17442 23278
rect 19406 23266 19458 23278
rect 17602 23214 17614 23266
rect 17666 23214 17678 23266
rect 17390 23202 17442 23214
rect 19406 23202 19458 23214
rect 21198 23266 21250 23278
rect 21198 23202 21250 23214
rect 12798 23154 12850 23166
rect 18286 23154 18338 23166
rect 16818 23102 16830 23154
rect 16882 23102 16894 23154
rect 12798 23090 12850 23102
rect 18286 23090 18338 23102
rect 18846 23154 18898 23166
rect 20078 23154 20130 23166
rect 19170 23102 19182 23154
rect 19234 23102 19246 23154
rect 19730 23102 19742 23154
rect 19794 23102 19806 23154
rect 18846 23090 18898 23102
rect 20078 23090 20130 23102
rect 20190 23154 20242 23166
rect 20190 23090 20242 23102
rect 20526 23154 20578 23166
rect 21422 23154 21474 23166
rect 20962 23102 20974 23154
rect 21026 23102 21038 23154
rect 20526 23090 20578 23102
rect 21422 23090 21474 23102
rect 21758 23154 21810 23166
rect 21758 23090 21810 23102
rect 23550 23154 23602 23166
rect 23550 23090 23602 23102
rect 23774 23154 23826 23166
rect 24098 23102 24110 23154
rect 24162 23102 24174 23154
rect 25218 23102 25230 23154
rect 25282 23102 25294 23154
rect 28466 23102 28478 23154
rect 28530 23102 28542 23154
rect 37650 23102 37662 23154
rect 37714 23102 37726 23154
rect 23774 23090 23826 23102
rect 13246 23042 13298 23054
rect 18062 23042 18114 23054
rect 13906 22990 13918 23042
rect 13970 22990 13982 23042
rect 16034 22990 16046 23042
rect 16098 22990 16110 23042
rect 13246 22978 13298 22990
rect 18062 22978 18114 22990
rect 22094 23042 22146 23054
rect 26002 22990 26014 23042
rect 26066 22990 26078 23042
rect 28130 22990 28142 23042
rect 28194 22990 28206 23042
rect 29250 22990 29262 23042
rect 29314 22990 29326 23042
rect 31378 22990 31390 23042
rect 31442 22990 31454 23042
rect 22094 22978 22146 22990
rect 17838 22930 17890 22942
rect 17838 22866 17890 22878
rect 22206 22930 22258 22942
rect 22206 22866 22258 22878
rect 40014 22930 40066 22942
rect 40014 22866 40066 22878
rect 1344 22762 40656 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 40656 22762
rect 1344 22676 40656 22710
rect 16046 22594 16098 22606
rect 16046 22530 16098 22542
rect 17726 22594 17778 22606
rect 17726 22530 17778 22542
rect 20414 22594 20466 22606
rect 20414 22530 20466 22542
rect 25118 22594 25170 22606
rect 25118 22530 25170 22542
rect 15934 22482 15986 22494
rect 15934 22418 15986 22430
rect 17054 22482 17106 22494
rect 17054 22418 17106 22430
rect 23550 22482 23602 22494
rect 23550 22418 23602 22430
rect 27134 22482 27186 22494
rect 27134 22418 27186 22430
rect 28590 22482 28642 22494
rect 28590 22418 28642 22430
rect 22542 22370 22594 22382
rect 24782 22370 24834 22382
rect 19170 22318 19182 22370
rect 19234 22318 19246 22370
rect 19842 22318 19854 22370
rect 19906 22318 19918 22370
rect 20402 22318 20414 22370
rect 20466 22318 20478 22370
rect 21410 22318 21422 22370
rect 21474 22318 21486 22370
rect 24546 22318 24558 22370
rect 24610 22318 24622 22370
rect 22542 22306 22594 22318
rect 24782 22306 24834 22318
rect 25006 22370 25058 22382
rect 25006 22306 25058 22318
rect 26126 22370 26178 22382
rect 27694 22370 27746 22382
rect 27346 22318 27358 22370
rect 27410 22318 27422 22370
rect 26126 22306 26178 22318
rect 27694 22306 27746 22318
rect 18062 22258 18114 22270
rect 18062 22194 18114 22206
rect 18398 22258 18450 22270
rect 20750 22258 20802 22270
rect 20066 22206 20078 22258
rect 20130 22206 20142 22258
rect 18398 22194 18450 22206
rect 20750 22194 20802 22206
rect 26014 22258 26066 22270
rect 26014 22194 26066 22206
rect 26238 22258 26290 22270
rect 26238 22194 26290 22206
rect 27246 22258 27298 22270
rect 27246 22194 27298 22206
rect 17838 22146 17890 22158
rect 17838 22082 17890 22094
rect 18510 22146 18562 22158
rect 18510 22082 18562 22094
rect 18734 22146 18786 22158
rect 21982 22146 22034 22158
rect 22878 22146 22930 22158
rect 18946 22094 18958 22146
rect 19010 22094 19022 22146
rect 21634 22094 21646 22146
rect 21698 22094 21710 22146
rect 22306 22094 22318 22146
rect 22370 22094 22382 22146
rect 18734 22082 18786 22094
rect 21982 22082 22034 22094
rect 22878 22082 22930 22094
rect 23102 22146 23154 22158
rect 23102 22082 23154 22094
rect 23214 22146 23266 22158
rect 23214 22082 23266 22094
rect 23438 22146 23490 22158
rect 23438 22082 23490 22094
rect 23662 22146 23714 22158
rect 23662 22082 23714 22094
rect 23886 22146 23938 22158
rect 23886 22082 23938 22094
rect 27022 22146 27074 22158
rect 27022 22082 27074 22094
rect 28142 22146 28194 22158
rect 28142 22082 28194 22094
rect 28478 22146 28530 22158
rect 28478 22082 28530 22094
rect 1344 21978 40656 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 40656 21978
rect 1344 21892 40656 21926
rect 22990 21810 23042 21822
rect 22990 21746 23042 21758
rect 23102 21698 23154 21710
rect 17714 21646 17726 21698
rect 17778 21646 17790 21698
rect 23102 21634 23154 21646
rect 24222 21698 24274 21710
rect 24222 21634 24274 21646
rect 27022 21698 27074 21710
rect 27022 21634 27074 21646
rect 27246 21698 27298 21710
rect 27246 21634 27298 21646
rect 27358 21698 27410 21710
rect 27458 21646 27470 21698
rect 27522 21646 27534 21698
rect 27358 21634 27410 21646
rect 23214 21586 23266 21598
rect 24110 21586 24162 21598
rect 22642 21534 22654 21586
rect 22706 21534 22718 21586
rect 23538 21534 23550 21586
rect 23602 21534 23614 21586
rect 23214 21522 23266 21534
rect 24110 21522 24162 21534
rect 24670 21586 24722 21598
rect 37874 21534 37886 21586
rect 37938 21534 37950 21586
rect 24670 21522 24722 21534
rect 24446 21474 24498 21486
rect 27346 21422 27358 21474
rect 27410 21422 27422 21474
rect 39890 21422 39902 21474
rect 39954 21422 39966 21474
rect 24446 21410 24498 21422
rect 1344 21194 40656 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 40656 21194
rect 1344 21108 40656 21142
rect 18386 20974 18398 21026
rect 18450 20974 18462 21026
rect 18834 20974 18846 21026
rect 18898 20974 18910 21026
rect 17278 20914 17330 20926
rect 40014 20914 40066 20926
rect 20290 20862 20302 20914
rect 20354 20862 20366 20914
rect 22642 20862 22654 20914
rect 22706 20911 22718 20914
rect 23202 20911 23214 20914
rect 22706 20865 23214 20911
rect 22706 20862 22718 20865
rect 23202 20862 23214 20865
rect 23266 20862 23278 20914
rect 26338 20862 26350 20914
rect 26402 20862 26414 20914
rect 17278 20850 17330 20862
rect 40014 20850 40066 20862
rect 14814 20802 14866 20814
rect 14354 20750 14366 20802
rect 14418 20750 14430 20802
rect 14814 20738 14866 20750
rect 16942 20802 16994 20814
rect 17726 20802 17778 20814
rect 19518 20802 19570 20814
rect 17154 20750 17166 20802
rect 17218 20750 17230 20802
rect 19282 20750 19294 20802
rect 19346 20750 19358 20802
rect 16942 20738 16994 20750
rect 17726 20738 17778 20750
rect 19518 20738 19570 20750
rect 19854 20802 19906 20814
rect 19854 20738 19906 20750
rect 21198 20802 21250 20814
rect 21198 20738 21250 20750
rect 21534 20802 21586 20814
rect 21970 20750 21982 20802
rect 22034 20750 22046 20802
rect 22418 20750 22430 20802
rect 22482 20750 22494 20802
rect 23202 20750 23214 20802
rect 23266 20750 23278 20802
rect 37650 20750 37662 20802
rect 37714 20750 37726 20802
rect 21534 20738 21586 20750
rect 15486 20690 15538 20702
rect 15486 20626 15538 20638
rect 17838 20690 17890 20702
rect 17838 20626 17890 20638
rect 17950 20690 18002 20702
rect 17950 20626 18002 20638
rect 15374 20578 15426 20590
rect 15374 20514 15426 20526
rect 1344 20410 40656 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 40656 20410
rect 1344 20324 40656 20358
rect 17950 20242 18002 20254
rect 17950 20178 18002 20190
rect 16270 20130 16322 20142
rect 25678 20130 25730 20142
rect 11666 20078 11678 20130
rect 11730 20078 11742 20130
rect 23202 20078 23214 20130
rect 23266 20078 23278 20130
rect 27570 20078 27582 20130
rect 27634 20078 27646 20130
rect 16270 20066 16322 20078
rect 25678 20066 25730 20078
rect 19070 20018 19122 20030
rect 10994 19966 11006 20018
rect 11058 19966 11070 20018
rect 14354 19966 14366 20018
rect 14418 19966 14430 20018
rect 14802 19966 14814 20018
rect 14866 19966 14878 20018
rect 19506 19966 19518 20018
rect 19570 19966 19582 20018
rect 25218 19966 25230 20018
rect 25282 19966 25294 20018
rect 25442 19966 25454 20018
rect 25506 19966 25518 20018
rect 26898 19966 26910 20018
rect 26962 19966 26974 20018
rect 19070 19954 19122 19966
rect 14142 19906 14194 19918
rect 18510 19906 18562 19918
rect 13794 19854 13806 19906
rect 13858 19854 13870 19906
rect 16706 19854 16718 19906
rect 16770 19854 16782 19906
rect 14142 19842 14194 19854
rect 18510 19842 18562 19854
rect 25342 19906 25394 19918
rect 30158 19906 30210 19918
rect 29698 19854 29710 19906
rect 29762 19854 29774 19906
rect 25342 19842 25394 19854
rect 30158 19842 30210 19854
rect 1344 19626 40656 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 40656 19626
rect 1344 19540 40656 19574
rect 17726 19458 17778 19470
rect 17726 19394 17778 19406
rect 21198 19458 21250 19470
rect 21198 19394 21250 19406
rect 29150 19458 29202 19470
rect 29150 19394 29202 19406
rect 19854 19346 19906 19358
rect 29262 19346 29314 19358
rect 12898 19294 12910 19346
rect 12962 19294 12974 19346
rect 24546 19294 24558 19346
rect 24610 19294 24622 19346
rect 26674 19294 26686 19346
rect 26738 19294 26750 19346
rect 19854 19282 19906 19294
rect 29262 19282 29314 19294
rect 13806 19234 13858 19246
rect 15486 19234 15538 19246
rect 10098 19182 10110 19234
rect 10162 19182 10174 19234
rect 14802 19182 14814 19234
rect 14866 19182 14878 19234
rect 13806 19170 13858 19182
rect 15486 19170 15538 19182
rect 16046 19234 16098 19246
rect 20078 19234 20130 19246
rect 19282 19182 19294 19234
rect 19346 19182 19358 19234
rect 16046 19170 16098 19182
rect 20078 19170 20130 19182
rect 21310 19234 21362 19246
rect 23102 19234 23154 19246
rect 21858 19182 21870 19234
rect 21922 19182 21934 19234
rect 22530 19182 22542 19234
rect 22594 19182 22606 19234
rect 23874 19182 23886 19234
rect 23938 19182 23950 19234
rect 21310 19170 21362 19182
rect 23102 19170 23154 19182
rect 13470 19122 13522 19134
rect 17838 19122 17890 19134
rect 10770 19070 10782 19122
rect 10834 19070 10846 19122
rect 17042 19070 17054 19122
rect 17106 19070 17118 19122
rect 21522 19070 21534 19122
rect 21586 19070 21598 19122
rect 13470 19058 13522 19070
rect 17838 19058 17890 19070
rect 14254 19010 14306 19022
rect 16718 19010 16770 19022
rect 27134 19010 27186 19022
rect 15026 18958 15038 19010
rect 15090 18958 15102 19010
rect 19506 18958 19518 19010
rect 19570 18958 19582 19010
rect 20402 18958 20414 19010
rect 20466 18958 20478 19010
rect 23426 18958 23438 19010
rect 23490 18958 23502 19010
rect 14254 18946 14306 18958
rect 16718 18946 16770 18958
rect 27134 18946 27186 18958
rect 1344 18842 40656 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 40656 18842
rect 1344 18756 40656 18790
rect 16270 18674 16322 18686
rect 25902 18674 25954 18686
rect 23314 18622 23326 18674
rect 23378 18622 23390 18674
rect 16270 18610 16322 18622
rect 25902 18610 25954 18622
rect 27022 18674 27074 18686
rect 27022 18610 27074 18622
rect 16382 18562 16434 18574
rect 25790 18562 25842 18574
rect 19618 18510 19630 18562
rect 19682 18510 19694 18562
rect 20402 18510 20414 18562
rect 20466 18510 20478 18562
rect 22754 18510 22766 18562
rect 22818 18510 22830 18562
rect 22978 18510 22990 18562
rect 23042 18510 23054 18562
rect 16382 18498 16434 18510
rect 25790 18498 25842 18510
rect 17614 18450 17666 18462
rect 17614 18386 17666 18398
rect 17950 18450 18002 18462
rect 17950 18386 18002 18398
rect 18510 18450 18562 18462
rect 23438 18450 23490 18462
rect 26014 18450 26066 18462
rect 18834 18398 18846 18450
rect 18898 18398 18910 18450
rect 20514 18398 20526 18450
rect 20578 18398 20590 18450
rect 25218 18398 25230 18450
rect 25282 18398 25294 18450
rect 25554 18398 25566 18450
rect 25618 18398 25630 18450
rect 18510 18386 18562 18398
rect 23438 18386 23490 18398
rect 26014 18386 26066 18398
rect 26574 18450 26626 18462
rect 26574 18386 26626 18398
rect 26798 18450 26850 18462
rect 26798 18386 26850 18398
rect 27246 18450 27298 18462
rect 37650 18398 37662 18450
rect 37714 18398 37726 18450
rect 27246 18386 27298 18398
rect 13134 18338 13186 18350
rect 13134 18274 13186 18286
rect 17502 18338 17554 18350
rect 21410 18286 21422 18338
rect 21474 18286 21486 18338
rect 27122 18286 27134 18338
rect 27186 18286 27198 18338
rect 17502 18274 17554 18286
rect 16270 18226 16322 18238
rect 16270 18162 16322 18174
rect 26350 18226 26402 18238
rect 26350 18162 26402 18174
rect 40014 18226 40066 18238
rect 40014 18162 40066 18174
rect 1344 18058 40656 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 40656 18058
rect 1344 17972 40656 18006
rect 21310 17890 21362 17902
rect 21310 17826 21362 17838
rect 21870 17890 21922 17902
rect 21870 17826 21922 17838
rect 29150 17890 29202 17902
rect 29150 17826 29202 17838
rect 24446 17778 24498 17790
rect 16146 17726 16158 17778
rect 16210 17726 16222 17778
rect 21634 17726 21646 17778
rect 21698 17726 21710 17778
rect 24446 17714 24498 17726
rect 17054 17666 17106 17678
rect 17054 17602 17106 17614
rect 18846 17666 18898 17678
rect 18846 17602 18898 17614
rect 19854 17666 19906 17678
rect 19854 17602 19906 17614
rect 20526 17666 20578 17678
rect 20526 17602 20578 17614
rect 21534 17666 21586 17678
rect 21534 17602 21586 17614
rect 22094 17666 22146 17678
rect 22094 17602 22146 17614
rect 22542 17666 22594 17678
rect 26014 17666 26066 17678
rect 24546 17614 24558 17666
rect 24610 17614 24622 17666
rect 22542 17602 22594 17614
rect 26014 17602 26066 17614
rect 26350 17666 26402 17678
rect 26350 17602 26402 17614
rect 14814 17554 14866 17566
rect 14814 17490 14866 17502
rect 14926 17554 14978 17566
rect 14926 17490 14978 17502
rect 16270 17554 16322 17566
rect 16270 17490 16322 17502
rect 16494 17554 16546 17566
rect 16494 17490 16546 17502
rect 16718 17554 16770 17566
rect 22654 17554 22706 17566
rect 18498 17502 18510 17554
rect 18562 17502 18574 17554
rect 20178 17502 20190 17554
rect 20242 17502 20254 17554
rect 16718 17490 16770 17502
rect 22654 17490 22706 17502
rect 24110 17554 24162 17566
rect 24110 17490 24162 17502
rect 24334 17554 24386 17566
rect 24334 17490 24386 17502
rect 29262 17554 29314 17566
rect 29262 17490 29314 17502
rect 14590 17442 14642 17454
rect 14590 17378 14642 17390
rect 16942 17442 16994 17454
rect 16942 17378 16994 17390
rect 18174 17442 18226 17454
rect 22878 17442 22930 17454
rect 19170 17390 19182 17442
rect 19234 17390 19246 17442
rect 19506 17390 19518 17442
rect 19570 17390 19582 17442
rect 18174 17378 18226 17390
rect 22878 17378 22930 17390
rect 23102 17442 23154 17454
rect 26126 17442 26178 17454
rect 23426 17390 23438 17442
rect 23490 17390 23502 17442
rect 23102 17378 23154 17390
rect 26126 17378 26178 17390
rect 1344 17274 40656 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 40656 17274
rect 1344 17188 40656 17222
rect 21646 17106 21698 17118
rect 17378 17054 17390 17106
rect 17442 17054 17454 17106
rect 21646 17042 21698 17054
rect 25790 17106 25842 17118
rect 25790 17042 25842 17054
rect 26014 17106 26066 17118
rect 26014 17042 26066 17054
rect 21534 16994 21586 17006
rect 21534 16930 21586 16942
rect 24110 16994 24162 17006
rect 24110 16930 24162 16942
rect 25566 16994 25618 17006
rect 27570 16942 27582 16994
rect 27634 16942 27646 16994
rect 25566 16930 25618 16942
rect 24334 16882 24386 16894
rect 4274 16830 4286 16882
rect 4338 16830 4350 16882
rect 12898 16830 12910 16882
rect 12962 16830 12974 16882
rect 13570 16830 13582 16882
rect 13634 16830 13646 16882
rect 24334 16818 24386 16830
rect 24782 16882 24834 16894
rect 30158 16882 30210 16894
rect 26226 16830 26238 16882
rect 26290 16830 26302 16882
rect 26898 16830 26910 16882
rect 26962 16830 26974 16882
rect 37650 16830 37662 16882
rect 37714 16830 37726 16882
rect 24782 16818 24834 16830
rect 30158 16818 30210 16830
rect 16158 16770 16210 16782
rect 15698 16718 15710 16770
rect 15762 16718 15774 16770
rect 16158 16706 16210 16718
rect 17726 16770 17778 16782
rect 17726 16706 17778 16718
rect 17950 16770 18002 16782
rect 17950 16706 18002 16718
rect 19966 16770 20018 16782
rect 19966 16706 20018 16718
rect 24558 16770 24610 16782
rect 24558 16706 24610 16718
rect 25902 16770 25954 16782
rect 29698 16718 29710 16770
rect 29762 16718 29774 16770
rect 25902 16706 25954 16718
rect 1934 16658 1986 16670
rect 1934 16594 1986 16606
rect 19854 16658 19906 16670
rect 19854 16594 19906 16606
rect 20190 16658 20242 16670
rect 20190 16594 20242 16606
rect 20302 16658 20354 16670
rect 20302 16594 20354 16606
rect 21646 16658 21698 16670
rect 21646 16594 21698 16606
rect 40014 16658 40066 16670
rect 40014 16594 40066 16606
rect 1344 16490 40656 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 40656 16490
rect 1344 16404 40656 16438
rect 15934 16322 15986 16334
rect 15934 16258 15986 16270
rect 18174 16322 18226 16334
rect 18174 16258 18226 16270
rect 29262 16210 29314 16222
rect 26450 16158 26462 16210
rect 26514 16158 26526 16210
rect 28578 16158 28590 16210
rect 28642 16158 28654 16210
rect 29262 16146 29314 16158
rect 15822 16098 15874 16110
rect 18062 16098 18114 16110
rect 16482 16046 16494 16098
rect 16546 16046 16558 16098
rect 16818 16046 16830 16098
rect 16882 16046 16894 16098
rect 15822 16034 15874 16046
rect 18062 16034 18114 16046
rect 20190 16098 20242 16110
rect 20190 16034 20242 16046
rect 24894 16098 24946 16110
rect 24894 16034 24946 16046
rect 25230 16098 25282 16110
rect 25778 16046 25790 16098
rect 25842 16046 25854 16098
rect 25230 16034 25282 16046
rect 14478 15986 14530 15998
rect 14478 15922 14530 15934
rect 16270 15986 16322 15998
rect 16270 15922 16322 15934
rect 16606 15986 16658 15998
rect 16606 15922 16658 15934
rect 14254 15874 14306 15886
rect 14254 15810 14306 15822
rect 14366 15874 14418 15886
rect 14366 15810 14418 15822
rect 17390 15874 17442 15886
rect 18174 15874 18226 15886
rect 17714 15822 17726 15874
rect 17778 15822 17790 15874
rect 17390 15810 17442 15822
rect 18174 15810 18226 15822
rect 19854 15874 19906 15886
rect 19854 15810 19906 15822
rect 20078 15874 20130 15886
rect 20078 15810 20130 15822
rect 25118 15874 25170 15886
rect 25118 15810 25170 15822
rect 1344 15706 40656 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 40656 15706
rect 1344 15620 40656 15654
rect 17502 15538 17554 15550
rect 17502 15474 17554 15486
rect 19182 15538 19234 15550
rect 19182 15474 19234 15486
rect 22990 15538 23042 15550
rect 22990 15474 23042 15486
rect 17614 15426 17666 15438
rect 23438 15426 23490 15438
rect 14354 15374 14366 15426
rect 14418 15374 14430 15426
rect 22642 15374 22654 15426
rect 22706 15374 22718 15426
rect 17614 15362 17666 15374
rect 23438 15362 23490 15374
rect 17278 15314 17330 15326
rect 15138 15262 15150 15314
rect 15202 15262 15214 15314
rect 17278 15250 17330 15262
rect 19406 15314 19458 15326
rect 20078 15314 20130 15326
rect 19506 15262 19518 15314
rect 19570 15262 19582 15314
rect 19406 15250 19458 15262
rect 20078 15250 20130 15262
rect 23662 15314 23714 15326
rect 23662 15250 23714 15262
rect 24110 15314 24162 15326
rect 24110 15250 24162 15262
rect 15598 15202 15650 15214
rect 19854 15202 19906 15214
rect 12226 15150 12238 15202
rect 12290 15150 12302 15202
rect 19282 15150 19294 15202
rect 19346 15150 19358 15202
rect 15598 15138 15650 15150
rect 19854 15138 19906 15150
rect 23886 15202 23938 15214
rect 23886 15138 23938 15150
rect 1344 14922 40656 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 40656 14922
rect 1344 14836 40656 14870
rect 19966 14754 20018 14766
rect 19966 14690 20018 14702
rect 21646 14754 21698 14766
rect 21646 14690 21698 14702
rect 19406 14642 19458 14654
rect 15474 14590 15486 14642
rect 15538 14590 15550 14642
rect 17602 14590 17614 14642
rect 17666 14590 17678 14642
rect 21298 14590 21310 14642
rect 21362 14590 21374 14642
rect 24210 14590 24222 14642
rect 24274 14590 24286 14642
rect 26338 14590 26350 14642
rect 26402 14590 26414 14642
rect 19406 14578 19458 14590
rect 20638 14530 20690 14542
rect 14802 14478 14814 14530
rect 14866 14478 14878 14530
rect 20290 14478 20302 14530
rect 20354 14478 20366 14530
rect 20638 14466 20690 14478
rect 22878 14530 22930 14542
rect 22878 14466 22930 14478
rect 23214 14530 23266 14542
rect 23426 14478 23438 14530
rect 23490 14478 23502 14530
rect 23214 14466 23266 14478
rect 19294 14418 19346 14430
rect 19294 14354 19346 14366
rect 18062 14306 18114 14318
rect 18062 14242 18114 14254
rect 19518 14306 19570 14318
rect 19518 14242 19570 14254
rect 20414 14306 20466 14318
rect 20414 14242 20466 14254
rect 20526 14306 20578 14318
rect 20526 14242 20578 14254
rect 21422 14306 21474 14318
rect 21422 14242 21474 14254
rect 22990 14306 23042 14318
rect 22990 14242 23042 14254
rect 26798 14306 26850 14318
rect 26798 14242 26850 14254
rect 1344 14138 40656 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 40656 14138
rect 1344 14052 40656 14086
rect 19282 13806 19294 13858
rect 19346 13806 19358 13858
rect 22530 13806 22542 13858
rect 22594 13806 22606 13858
rect 25342 13746 25394 13758
rect 18610 13694 18622 13746
rect 18674 13694 18686 13746
rect 21858 13694 21870 13746
rect 21922 13694 21934 13746
rect 25342 13682 25394 13694
rect 21410 13582 21422 13634
rect 21474 13582 21486 13634
rect 24658 13582 24670 13634
rect 24722 13582 24734 13634
rect 1344 13354 40656 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 40656 13354
rect 1344 13268 40656 13302
rect 21646 13074 21698 13086
rect 18610 13022 18622 13074
rect 18674 13022 18686 13074
rect 20738 13022 20750 13074
rect 20802 13022 20814 13074
rect 21646 13010 21698 13022
rect 17938 12910 17950 12962
rect 18002 12910 18014 12962
rect 1344 12570 40656 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 40656 12570
rect 1344 12484 40656 12518
rect 21086 12402 21138 12414
rect 21086 12338 21138 12350
rect 1344 11786 40656 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 40656 11786
rect 1344 11700 40656 11734
rect 1344 11002 40656 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 40656 11002
rect 1344 10916 40656 10950
rect 1344 10218 40656 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 40656 10218
rect 1344 10132 40656 10166
rect 1344 9434 40656 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 40656 9434
rect 1344 9348 40656 9382
rect 1344 8650 40656 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 40656 8650
rect 1344 8564 40656 8598
rect 1344 7866 40656 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 40656 7866
rect 1344 7780 40656 7814
rect 1344 7082 40656 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 40656 7082
rect 1344 6996 40656 7030
rect 1344 6298 40656 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 40656 6298
rect 1344 6212 40656 6246
rect 1344 5514 40656 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 40656 5514
rect 1344 5428 40656 5462
rect 1344 4730 40656 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 40656 4730
rect 1344 4644 40656 4678
rect 21074 4286 21086 4338
rect 21138 4286 21150 4338
rect 25778 4286 25790 4338
rect 25842 4286 25854 4338
rect 22094 4114 22146 4126
rect 22094 4050 22146 4062
rect 26798 4114 26850 4126
rect 26798 4050 26850 4062
rect 1344 3946 40656 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 40656 3946
rect 1344 3860 40656 3894
rect 22430 3666 22482 3678
rect 22430 3602 22482 3614
rect 25566 3666 25618 3678
rect 25566 3602 25618 3614
rect 21410 3502 21422 3554
rect 21474 3502 21486 3554
rect 24546 3502 24558 3554
rect 24610 3502 24622 3554
rect 16942 3330 16994 3342
rect 16942 3266 16994 3278
rect 1344 3162 40656 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 40656 3162
rect 1344 3076 40656 3110
<< via1 >>
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 22430 38222 22482 38274
rect 25566 38222 25618 38274
rect 18846 38110 18898 38162
rect 19742 37998 19794 38050
rect 21422 37998 21474 38050
rect 24558 37998 24610 38050
rect 27470 37886 27522 37938
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 18398 37438 18450 37490
rect 20750 37438 20802 37490
rect 19742 37214 19794 37266
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 18734 36654 18786 36706
rect 24782 36654 24834 36706
rect 17726 36430 17778 36482
rect 24110 36430 24162 36482
rect 1710 36318 1762 36370
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 18622 28590 18674 28642
rect 18174 28478 18226 28530
rect 18846 28478 18898 28530
rect 18958 28478 19010 28530
rect 19406 28478 19458 28530
rect 19518 28478 19570 28530
rect 17838 28366 17890 28418
rect 18062 28366 18114 28418
rect 19742 28366 19794 28418
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 24110 28030 24162 28082
rect 15038 27806 15090 27858
rect 17502 27806 17554 27858
rect 20974 27806 21026 27858
rect 24446 27806 24498 27858
rect 12126 27694 12178 27746
rect 14254 27694 14306 27746
rect 15598 27694 15650 27746
rect 18174 27694 18226 27746
rect 20302 27694 20354 27746
rect 21646 27694 21698 27746
rect 23774 27694 23826 27746
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 14142 27246 14194 27298
rect 1934 27134 1986 27186
rect 17166 27134 17218 27186
rect 19294 27134 19346 27186
rect 21646 27134 21698 27186
rect 22542 27134 22594 27186
rect 4286 27022 4338 27074
rect 16494 27022 16546 27074
rect 19518 27022 19570 27074
rect 19854 27022 19906 27074
rect 21422 27022 21474 27074
rect 21982 27022 22034 27074
rect 14142 26910 14194 26962
rect 14254 26910 14306 26962
rect 21758 26910 21810 26962
rect 22430 26910 22482 26962
rect 19742 26798 19794 26850
rect 20526 26798 20578 26850
rect 21534 26798 21586 26850
rect 23998 26798 24050 26850
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 23550 26350 23602 26402
rect 13918 26238 13970 26290
rect 22990 26238 23042 26290
rect 14702 26126 14754 26178
rect 16830 26126 16882 26178
rect 17502 26126 17554 26178
rect 19518 26126 19570 26178
rect 20190 26126 20242 26178
rect 22318 26126 22370 26178
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 15710 25678 15762 25730
rect 1934 25566 1986 25618
rect 16942 25566 16994 25618
rect 21870 25566 21922 25618
rect 22430 25566 22482 25618
rect 4286 25454 4338 25506
rect 14254 25454 14306 25506
rect 15822 25454 15874 25506
rect 16830 25454 16882 25506
rect 17054 25454 17106 25506
rect 12798 25342 12850 25394
rect 13582 25342 13634 25394
rect 13694 25342 13746 25394
rect 14478 25342 14530 25394
rect 14590 25342 14642 25394
rect 16158 25342 16210 25394
rect 17502 25342 17554 25394
rect 18622 25342 18674 25394
rect 21310 25342 21362 25394
rect 21870 25342 21922 25394
rect 12462 25230 12514 25282
rect 12686 25230 12738 25282
rect 13358 25230 13410 25282
rect 16494 25230 16546 25282
rect 17278 25230 17330 25282
rect 18286 25230 18338 25282
rect 21534 25230 21586 25282
rect 21758 25230 21810 25282
rect 22318 25230 22370 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 13918 24894 13970 24946
rect 20190 24894 20242 24946
rect 19966 24782 20018 24834
rect 24110 24782 24162 24834
rect 4286 24670 4338 24722
rect 13470 24670 13522 24722
rect 19854 24670 19906 24722
rect 23998 24670 24050 24722
rect 37662 24670 37714 24722
rect 10558 24558 10610 24610
rect 12686 24558 12738 24610
rect 1934 24446 1986 24498
rect 24110 24446 24162 24498
rect 40014 24446 40066 24498
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 1934 23998 1986 24050
rect 9998 23998 10050 24050
rect 12126 23998 12178 24050
rect 13582 23998 13634 24050
rect 20750 23998 20802 24050
rect 25678 23998 25730 24050
rect 40014 23998 40066 24050
rect 4286 23886 4338 23938
rect 12910 23886 12962 23938
rect 13470 23886 13522 23938
rect 13694 23886 13746 23938
rect 17838 23886 17890 23938
rect 18510 23886 18562 23938
rect 19630 23886 19682 23938
rect 20302 23886 20354 23938
rect 22878 23886 22930 23938
rect 37662 23886 37714 23938
rect 14030 23774 14082 23826
rect 18174 23774 18226 23826
rect 19966 23774 20018 23826
rect 20638 23774 20690 23826
rect 23550 23774 23602 23826
rect 26126 23662 26178 23714
rect 28366 23662 28418 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 12462 23326 12514 23378
rect 12686 23326 12738 23378
rect 17726 23326 17778 23378
rect 19518 23326 19570 23378
rect 20414 23326 20466 23378
rect 21646 23326 21698 23378
rect 23662 23326 23714 23378
rect 17390 23214 17442 23266
rect 17614 23214 17666 23266
rect 19406 23214 19458 23266
rect 21198 23214 21250 23266
rect 12798 23102 12850 23154
rect 16830 23102 16882 23154
rect 18286 23102 18338 23154
rect 18846 23102 18898 23154
rect 19182 23102 19234 23154
rect 19742 23102 19794 23154
rect 20078 23102 20130 23154
rect 20190 23102 20242 23154
rect 20526 23102 20578 23154
rect 20974 23102 21026 23154
rect 21422 23102 21474 23154
rect 21758 23102 21810 23154
rect 23550 23102 23602 23154
rect 23774 23102 23826 23154
rect 24110 23102 24162 23154
rect 25230 23102 25282 23154
rect 28478 23102 28530 23154
rect 37662 23102 37714 23154
rect 13246 22990 13298 23042
rect 13918 22990 13970 23042
rect 16046 22990 16098 23042
rect 18062 22990 18114 23042
rect 22094 22990 22146 23042
rect 26014 22990 26066 23042
rect 28142 22990 28194 23042
rect 29262 22990 29314 23042
rect 31390 22990 31442 23042
rect 17838 22878 17890 22930
rect 22206 22878 22258 22930
rect 40014 22878 40066 22930
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 16046 22542 16098 22594
rect 17726 22542 17778 22594
rect 20414 22542 20466 22594
rect 25118 22542 25170 22594
rect 15934 22430 15986 22482
rect 17054 22430 17106 22482
rect 23550 22430 23602 22482
rect 27134 22430 27186 22482
rect 28590 22430 28642 22482
rect 19182 22318 19234 22370
rect 19854 22318 19906 22370
rect 20414 22318 20466 22370
rect 21422 22318 21474 22370
rect 22542 22318 22594 22370
rect 24558 22318 24610 22370
rect 24782 22318 24834 22370
rect 25006 22318 25058 22370
rect 26126 22318 26178 22370
rect 27358 22318 27410 22370
rect 27694 22318 27746 22370
rect 18062 22206 18114 22258
rect 18398 22206 18450 22258
rect 20078 22206 20130 22258
rect 20750 22206 20802 22258
rect 26014 22206 26066 22258
rect 26238 22206 26290 22258
rect 27246 22206 27298 22258
rect 17838 22094 17890 22146
rect 18510 22094 18562 22146
rect 18734 22094 18786 22146
rect 18958 22094 19010 22146
rect 21646 22094 21698 22146
rect 21982 22094 22034 22146
rect 22318 22094 22370 22146
rect 22878 22094 22930 22146
rect 23102 22094 23154 22146
rect 23214 22094 23266 22146
rect 23438 22094 23490 22146
rect 23662 22094 23714 22146
rect 23886 22094 23938 22146
rect 27022 22094 27074 22146
rect 28142 22094 28194 22146
rect 28478 22094 28530 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 22990 21758 23042 21810
rect 17726 21646 17778 21698
rect 23102 21646 23154 21698
rect 24222 21646 24274 21698
rect 27022 21646 27074 21698
rect 27246 21646 27298 21698
rect 27358 21646 27410 21698
rect 27470 21646 27522 21698
rect 22654 21534 22706 21586
rect 23214 21534 23266 21586
rect 23550 21534 23602 21586
rect 24110 21534 24162 21586
rect 24670 21534 24722 21586
rect 37886 21534 37938 21586
rect 24446 21422 24498 21474
rect 27358 21422 27410 21474
rect 39902 21422 39954 21474
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 18398 20974 18450 21026
rect 18846 20974 18898 21026
rect 17278 20862 17330 20914
rect 20302 20862 20354 20914
rect 22654 20862 22706 20914
rect 23214 20862 23266 20914
rect 26350 20862 26402 20914
rect 40014 20862 40066 20914
rect 14366 20750 14418 20802
rect 14814 20750 14866 20802
rect 16942 20750 16994 20802
rect 17166 20750 17218 20802
rect 17726 20750 17778 20802
rect 19294 20750 19346 20802
rect 19518 20750 19570 20802
rect 19854 20750 19906 20802
rect 21198 20750 21250 20802
rect 21534 20750 21586 20802
rect 21982 20750 22034 20802
rect 22430 20750 22482 20802
rect 23214 20750 23266 20802
rect 37662 20750 37714 20802
rect 15486 20638 15538 20690
rect 17838 20638 17890 20690
rect 17950 20638 18002 20690
rect 15374 20526 15426 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 17950 20190 18002 20242
rect 11678 20078 11730 20130
rect 16270 20078 16322 20130
rect 23214 20078 23266 20130
rect 25678 20078 25730 20130
rect 27582 20078 27634 20130
rect 11006 19966 11058 20018
rect 14366 19966 14418 20018
rect 14814 19966 14866 20018
rect 19070 19966 19122 20018
rect 19518 19966 19570 20018
rect 25230 19966 25282 20018
rect 25454 19966 25506 20018
rect 26910 19966 26962 20018
rect 13806 19854 13858 19906
rect 14142 19854 14194 19906
rect 16718 19854 16770 19906
rect 18510 19854 18562 19906
rect 25342 19854 25394 19906
rect 29710 19854 29762 19906
rect 30158 19854 30210 19906
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 17726 19406 17778 19458
rect 21198 19406 21250 19458
rect 29150 19406 29202 19458
rect 12910 19294 12962 19346
rect 19854 19294 19906 19346
rect 24558 19294 24610 19346
rect 26686 19294 26738 19346
rect 29262 19294 29314 19346
rect 10110 19182 10162 19234
rect 13806 19182 13858 19234
rect 14814 19182 14866 19234
rect 15486 19182 15538 19234
rect 16046 19182 16098 19234
rect 19294 19182 19346 19234
rect 20078 19182 20130 19234
rect 21310 19182 21362 19234
rect 21870 19182 21922 19234
rect 22542 19182 22594 19234
rect 23102 19182 23154 19234
rect 23886 19182 23938 19234
rect 10782 19070 10834 19122
rect 13470 19070 13522 19122
rect 17054 19070 17106 19122
rect 17838 19070 17890 19122
rect 21534 19070 21586 19122
rect 14254 18958 14306 19010
rect 15038 18958 15090 19010
rect 16718 18958 16770 19010
rect 19518 18958 19570 19010
rect 20414 18958 20466 19010
rect 23438 18958 23490 19010
rect 27134 18958 27186 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 16270 18622 16322 18674
rect 23326 18622 23378 18674
rect 25902 18622 25954 18674
rect 27022 18622 27074 18674
rect 16382 18510 16434 18562
rect 19630 18510 19682 18562
rect 20414 18510 20466 18562
rect 22766 18510 22818 18562
rect 22990 18510 23042 18562
rect 25790 18510 25842 18562
rect 17614 18398 17666 18450
rect 17950 18398 18002 18450
rect 18510 18398 18562 18450
rect 18846 18398 18898 18450
rect 20526 18398 20578 18450
rect 23438 18398 23490 18450
rect 25230 18398 25282 18450
rect 25566 18398 25618 18450
rect 26014 18398 26066 18450
rect 26574 18398 26626 18450
rect 26798 18398 26850 18450
rect 27246 18398 27298 18450
rect 37662 18398 37714 18450
rect 13134 18286 13186 18338
rect 17502 18286 17554 18338
rect 21422 18286 21474 18338
rect 27134 18286 27186 18338
rect 16270 18174 16322 18226
rect 26350 18174 26402 18226
rect 40014 18174 40066 18226
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 21310 17838 21362 17890
rect 21870 17838 21922 17890
rect 29150 17838 29202 17890
rect 16158 17726 16210 17778
rect 21646 17726 21698 17778
rect 24446 17726 24498 17778
rect 17054 17614 17106 17666
rect 18846 17614 18898 17666
rect 19854 17614 19906 17666
rect 20526 17614 20578 17666
rect 21534 17614 21586 17666
rect 22094 17614 22146 17666
rect 22542 17614 22594 17666
rect 24558 17614 24610 17666
rect 26014 17614 26066 17666
rect 26350 17614 26402 17666
rect 14814 17502 14866 17554
rect 14926 17502 14978 17554
rect 16270 17502 16322 17554
rect 16494 17502 16546 17554
rect 16718 17502 16770 17554
rect 18510 17502 18562 17554
rect 20190 17502 20242 17554
rect 22654 17502 22706 17554
rect 24110 17502 24162 17554
rect 24334 17502 24386 17554
rect 29262 17502 29314 17554
rect 14590 17390 14642 17442
rect 16942 17390 16994 17442
rect 18174 17390 18226 17442
rect 19182 17390 19234 17442
rect 19518 17390 19570 17442
rect 22878 17390 22930 17442
rect 23102 17390 23154 17442
rect 23438 17390 23490 17442
rect 26126 17390 26178 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 17390 17054 17442 17106
rect 21646 17054 21698 17106
rect 25790 17054 25842 17106
rect 26014 17054 26066 17106
rect 21534 16942 21586 16994
rect 24110 16942 24162 16994
rect 25566 16942 25618 16994
rect 27582 16942 27634 16994
rect 4286 16830 4338 16882
rect 12910 16830 12962 16882
rect 13582 16830 13634 16882
rect 24334 16830 24386 16882
rect 24782 16830 24834 16882
rect 26238 16830 26290 16882
rect 26910 16830 26962 16882
rect 30158 16830 30210 16882
rect 37662 16830 37714 16882
rect 15710 16718 15762 16770
rect 16158 16718 16210 16770
rect 17726 16718 17778 16770
rect 17950 16718 18002 16770
rect 19966 16718 20018 16770
rect 24558 16718 24610 16770
rect 25902 16718 25954 16770
rect 29710 16718 29762 16770
rect 1934 16606 1986 16658
rect 19854 16606 19906 16658
rect 20190 16606 20242 16658
rect 20302 16606 20354 16658
rect 21646 16606 21698 16658
rect 40014 16606 40066 16658
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 15934 16270 15986 16322
rect 18174 16270 18226 16322
rect 26462 16158 26514 16210
rect 28590 16158 28642 16210
rect 29262 16158 29314 16210
rect 15822 16046 15874 16098
rect 16494 16046 16546 16098
rect 16830 16046 16882 16098
rect 18062 16046 18114 16098
rect 20190 16046 20242 16098
rect 24894 16046 24946 16098
rect 25230 16046 25282 16098
rect 25790 16046 25842 16098
rect 14478 15934 14530 15986
rect 16270 15934 16322 15986
rect 16606 15934 16658 15986
rect 14254 15822 14306 15874
rect 14366 15822 14418 15874
rect 17390 15822 17442 15874
rect 17726 15822 17778 15874
rect 18174 15822 18226 15874
rect 19854 15822 19906 15874
rect 20078 15822 20130 15874
rect 25118 15822 25170 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 17502 15486 17554 15538
rect 19182 15486 19234 15538
rect 22990 15486 23042 15538
rect 14366 15374 14418 15426
rect 17614 15374 17666 15426
rect 22654 15374 22706 15426
rect 23438 15374 23490 15426
rect 15150 15262 15202 15314
rect 17278 15262 17330 15314
rect 19406 15262 19458 15314
rect 19518 15262 19570 15314
rect 20078 15262 20130 15314
rect 23662 15262 23714 15314
rect 24110 15262 24162 15314
rect 12238 15150 12290 15202
rect 15598 15150 15650 15202
rect 19294 15150 19346 15202
rect 19854 15150 19906 15202
rect 23886 15150 23938 15202
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 19966 14702 20018 14754
rect 21646 14702 21698 14754
rect 15486 14590 15538 14642
rect 17614 14590 17666 14642
rect 19406 14590 19458 14642
rect 21310 14590 21362 14642
rect 24222 14590 24274 14642
rect 26350 14590 26402 14642
rect 14814 14478 14866 14530
rect 20302 14478 20354 14530
rect 20638 14478 20690 14530
rect 22878 14478 22930 14530
rect 23214 14478 23266 14530
rect 23438 14478 23490 14530
rect 19294 14366 19346 14418
rect 18062 14254 18114 14306
rect 19518 14254 19570 14306
rect 20414 14254 20466 14306
rect 20526 14254 20578 14306
rect 21422 14254 21474 14306
rect 22990 14254 23042 14306
rect 26798 14254 26850 14306
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 19294 13806 19346 13858
rect 22542 13806 22594 13858
rect 18622 13694 18674 13746
rect 21870 13694 21922 13746
rect 25342 13694 25394 13746
rect 21422 13582 21474 13634
rect 24670 13582 24722 13634
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 18622 13022 18674 13074
rect 20750 13022 20802 13074
rect 21646 13022 21698 13074
rect 17950 12910 18002 12962
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 21086 12350 21138 12402
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 21086 4286 21138 4338
rect 25790 4286 25842 4338
rect 22094 4062 22146 4114
rect 26798 4062 26850 4114
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 22430 3614 22482 3666
rect 25566 3614 25618 3666
rect 21422 3502 21474 3554
rect 24558 3502 24610 3554
rect 16942 3278 16994 3330
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
<< metal2 >>
rect 17472 41200 17584 42000
rect 18144 41200 18256 42000
rect 18816 41200 18928 42000
rect 19488 41200 19600 42000
rect 22176 41200 22288 42000
rect 22848 41200 22960 42000
rect 23520 41200 23632 42000
rect 26208 41200 26320 42000
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 17500 36708 17556 41200
rect 18172 37492 18228 41200
rect 18844 38162 18900 41200
rect 19516 38612 19572 41200
rect 19516 38546 19572 38556
rect 20748 38612 20804 38622
rect 18844 38110 18846 38162
rect 18898 38110 18900 38162
rect 18844 38098 18900 38110
rect 19740 38052 19796 38062
rect 19068 38050 19796 38052
rect 19068 37998 19742 38050
rect 19794 37998 19796 38050
rect 19068 37996 19796 37998
rect 18396 37492 18452 37502
rect 18172 37490 18452 37492
rect 18172 37438 18398 37490
rect 18450 37438 18452 37490
rect 18172 37436 18452 37438
rect 18396 37426 18452 37436
rect 17500 36642 17556 36652
rect 18732 36708 18788 36718
rect 18732 36614 18788 36652
rect 17724 36482 17780 36494
rect 17724 36430 17726 36482
rect 17778 36430 17780 36482
rect 1708 36372 1764 36382
rect 1708 36278 1764 36316
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 16828 28868 16884 28878
rect 15036 27858 15092 27870
rect 15036 27806 15038 27858
rect 15090 27806 15092 27858
rect 12124 27746 12180 27758
rect 14252 27748 14308 27758
rect 12124 27694 12126 27746
rect 12178 27694 12180 27746
rect 4172 27636 4228 27646
rect 1932 27188 1988 27198
rect 1932 27094 1988 27132
rect 1932 25618 1988 25630
rect 1932 25566 1934 25618
rect 1986 25566 1988 25618
rect 1932 24948 1988 25566
rect 1932 24882 1988 24892
rect 1932 24500 1988 24510
rect 1932 24406 1988 24444
rect 1932 24050 1988 24062
rect 1932 23998 1934 24050
rect 1986 23998 1988 24050
rect 1932 23604 1988 23998
rect 1932 23538 1988 23548
rect 4172 20020 4228 27580
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 12124 27188 12180 27694
rect 14140 27746 14308 27748
rect 14140 27694 14254 27746
rect 14306 27694 14308 27746
rect 14140 27692 14308 27694
rect 14140 27298 14196 27692
rect 14252 27682 14308 27692
rect 15036 27748 15092 27806
rect 15036 27682 15092 27692
rect 15596 27748 15652 27758
rect 15596 27654 15652 27692
rect 16492 27748 16548 27758
rect 14140 27246 14142 27298
rect 14194 27246 14196 27298
rect 14140 27234 14196 27246
rect 12124 27122 12180 27132
rect 14476 27188 14532 27198
rect 4284 27076 4340 27086
rect 4284 26982 4340 27020
rect 14140 27076 14196 27086
rect 14140 26962 14196 27020
rect 14140 26910 14142 26962
rect 14194 26910 14196 26962
rect 14140 26898 14196 26910
rect 14252 26962 14308 26974
rect 14252 26910 14254 26962
rect 14306 26910 14308 26962
rect 13916 26290 13972 26302
rect 13916 26238 13918 26290
rect 13970 26238 13972 26290
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 4284 25508 4340 25518
rect 4284 25414 4340 25452
rect 10556 25508 10612 25518
rect 4284 24724 4340 24734
rect 4284 24630 4340 24668
rect 9996 24724 10052 24734
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 9996 24052 10052 24668
rect 10556 24610 10612 25452
rect 13580 25508 13636 25518
rect 12796 25394 12852 25406
rect 12796 25342 12798 25394
rect 12850 25342 12852 25394
rect 12460 25284 12516 25294
rect 10556 24558 10558 24610
rect 10610 24558 10612 24610
rect 10556 24546 10612 24558
rect 12124 25282 12516 25284
rect 12124 25230 12462 25282
rect 12514 25230 12516 25282
rect 12124 25228 12516 25230
rect 9996 23958 10052 23996
rect 12124 24050 12180 25228
rect 12460 25218 12516 25228
rect 12684 25282 12740 25294
rect 12684 25230 12686 25282
rect 12738 25230 12740 25282
rect 12684 24836 12740 25230
rect 12124 23998 12126 24050
rect 12178 23998 12180 24050
rect 12124 23986 12180 23998
rect 12348 24780 12740 24836
rect 4284 23940 4340 23950
rect 4284 23846 4340 23884
rect 12348 23156 12404 24780
rect 12684 24612 12740 24622
rect 12460 24610 12740 24612
rect 12460 24558 12686 24610
rect 12738 24558 12740 24610
rect 12460 24556 12740 24558
rect 12460 23378 12516 24556
rect 12684 24546 12740 24556
rect 12796 24388 12852 25342
rect 13580 25394 13636 25452
rect 13580 25342 13582 25394
rect 13634 25342 13636 25394
rect 13580 25330 13636 25342
rect 13692 25396 13748 25406
rect 13356 25282 13412 25294
rect 13356 25230 13358 25282
rect 13410 25230 13412 25282
rect 13356 24948 13412 25230
rect 13692 25060 13748 25340
rect 13580 25004 13748 25060
rect 12796 24322 12852 24332
rect 13132 24892 13412 24948
rect 13468 24948 13524 24958
rect 13132 24164 13188 24892
rect 13468 24724 13524 24892
rect 12460 23326 12462 23378
rect 12514 23326 12516 23378
rect 12460 23314 12516 23326
rect 12684 24108 13188 24164
rect 13356 24722 13524 24724
rect 13356 24670 13470 24722
rect 13522 24670 13524 24722
rect 13356 24668 13524 24670
rect 12684 23378 12740 24108
rect 12684 23326 12686 23378
rect 12738 23326 12740 23378
rect 12684 23314 12740 23326
rect 12908 23938 12964 23950
rect 12908 23886 12910 23938
rect 12962 23886 12964 23938
rect 12796 23156 12852 23166
rect 12348 23154 12852 23156
rect 12348 23102 12798 23154
rect 12850 23102 12852 23154
rect 12348 23100 12852 23102
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 12796 22596 12852 23100
rect 12908 23044 12964 23886
rect 13244 23044 13300 23054
rect 13356 23044 13412 24668
rect 13468 24658 13524 24668
rect 13580 24500 13636 25004
rect 13916 24948 13972 26238
rect 14252 25506 14308 26910
rect 14252 25454 14254 25506
rect 14306 25454 14308 25506
rect 14252 25442 14308 25454
rect 14476 25394 14532 27132
rect 16492 27074 16548 27692
rect 16492 27022 16494 27074
rect 16546 27022 16548 27074
rect 14700 26180 14756 26190
rect 14700 26086 14756 26124
rect 15708 26180 15764 26190
rect 15708 25730 15764 26124
rect 16492 26180 16548 27022
rect 16492 26114 16548 26124
rect 16828 26180 16884 28812
rect 17724 28868 17780 36430
rect 19068 31948 19124 37996
rect 19740 37986 19796 37996
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 20748 37490 20804 38556
rect 22204 38276 22260 41200
rect 22428 38276 22484 38286
rect 22204 38274 22484 38276
rect 22204 38222 22430 38274
rect 22482 38222 22484 38274
rect 22204 38220 22484 38222
rect 22428 38210 22484 38220
rect 22876 38276 22932 41200
rect 22876 38210 22932 38220
rect 20748 37438 20750 37490
rect 20802 37438 20804 37490
rect 20748 37426 20804 37438
rect 21420 38050 21476 38062
rect 21420 37998 21422 38050
rect 21474 37998 21476 38050
rect 19740 37268 19796 37278
rect 17724 28802 17780 28812
rect 18844 31892 19124 31948
rect 19516 37266 19796 37268
rect 19516 37214 19742 37266
rect 19794 37214 19796 37266
rect 19516 37212 19796 37214
rect 18620 28644 18676 28654
rect 18172 28642 18676 28644
rect 18172 28590 18622 28642
rect 18674 28590 18676 28642
rect 18172 28588 18676 28590
rect 18172 28530 18228 28588
rect 18620 28578 18676 28588
rect 18172 28478 18174 28530
rect 18226 28478 18228 28530
rect 18172 28466 18228 28478
rect 18844 28530 18900 31892
rect 18844 28478 18846 28530
rect 18898 28478 18900 28530
rect 17836 28420 17892 28430
rect 18060 28420 18116 28430
rect 17164 28418 17892 28420
rect 17164 28366 17838 28418
rect 17890 28366 17892 28418
rect 17164 28364 17892 28366
rect 17164 27186 17220 28364
rect 17836 28354 17892 28364
rect 17948 28418 18116 28420
rect 17948 28366 18062 28418
rect 18114 28366 18116 28418
rect 17948 28364 18116 28366
rect 17948 28084 18004 28364
rect 18060 28354 18116 28364
rect 18844 28308 18900 28478
rect 18956 28532 19012 28542
rect 19404 28532 19460 28542
rect 18956 28530 19460 28532
rect 18956 28478 18958 28530
rect 19010 28478 19406 28530
rect 19458 28478 19460 28530
rect 18956 28476 19460 28478
rect 18956 28466 19012 28476
rect 18844 28252 19348 28308
rect 17164 27134 17166 27186
rect 17218 27134 17220 27186
rect 17164 27122 17220 27134
rect 17388 28028 18004 28084
rect 16828 26178 17108 26180
rect 16828 26126 16830 26178
rect 16882 26126 17108 26178
rect 16828 26124 17108 26126
rect 16828 26114 16884 26124
rect 15708 25678 15710 25730
rect 15762 25678 15764 25730
rect 15708 25666 15764 25678
rect 16940 25618 16996 25630
rect 16940 25566 16942 25618
rect 16994 25566 16996 25618
rect 15820 25508 15876 25518
rect 15820 25414 15876 25452
rect 16828 25506 16884 25518
rect 16828 25454 16830 25506
rect 16882 25454 16884 25506
rect 14476 25342 14478 25394
rect 14530 25342 14532 25394
rect 14476 25330 14532 25342
rect 14588 25396 14644 25406
rect 14588 25302 14644 25340
rect 16156 25396 16212 25406
rect 16156 25302 16212 25340
rect 16828 25396 16884 25454
rect 16940 25508 16996 25566
rect 16940 25442 16996 25452
rect 17052 25506 17108 26124
rect 17052 25454 17054 25506
rect 17106 25454 17108 25506
rect 17052 25442 17108 25454
rect 16828 25330 16884 25340
rect 16492 25284 16548 25294
rect 17276 25284 17332 25294
rect 16492 25190 16548 25228
rect 17164 25282 17332 25284
rect 17164 25230 17278 25282
rect 17330 25230 17332 25282
rect 17164 25228 17332 25230
rect 13916 24854 13972 24892
rect 17052 25172 17108 25182
rect 13468 24444 13636 24500
rect 13468 23938 13524 24444
rect 13580 24276 13636 24286
rect 13580 24050 13636 24220
rect 13580 23998 13582 24050
rect 13634 23998 13636 24050
rect 13580 23986 13636 23998
rect 13692 24052 13748 24062
rect 13468 23886 13470 23938
rect 13522 23886 13524 23938
rect 13468 23874 13524 23886
rect 13692 23938 13748 23996
rect 13692 23886 13694 23938
rect 13746 23886 13748 23938
rect 13692 23874 13748 23886
rect 13916 23940 13972 23950
rect 12908 22988 13244 23044
rect 13300 22988 13412 23044
rect 13916 23268 13972 23884
rect 13916 23042 13972 23212
rect 13916 22990 13918 23042
rect 13970 22990 13972 23042
rect 13244 22950 13300 22988
rect 13916 22978 13972 22990
rect 14028 23826 14084 23838
rect 14028 23774 14030 23826
rect 14082 23774 14084 23826
rect 14028 22932 14084 23774
rect 15932 23380 15988 23390
rect 15372 23156 15428 23166
rect 14028 22866 14084 22876
rect 15260 23044 15316 23054
rect 12796 22530 12852 22540
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 14364 20802 14420 20814
rect 14364 20750 14366 20802
rect 14418 20750 14420 20802
rect 11676 20580 11732 20590
rect 4172 19954 4228 19964
rect 10108 20132 10164 20142
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 10108 19234 10164 20076
rect 11004 20132 11060 20142
rect 11004 20018 11060 20076
rect 11676 20130 11732 20524
rect 11676 20078 11678 20130
rect 11730 20078 11732 20130
rect 11676 20066 11732 20078
rect 14252 20132 14308 20142
rect 11004 19966 11006 20018
rect 11058 19966 11060 20018
rect 11004 19954 11060 19966
rect 13804 19908 13860 19918
rect 14140 19908 14196 19918
rect 13804 19814 13860 19852
rect 13916 19906 14196 19908
rect 13916 19854 14142 19906
rect 14194 19854 14196 19906
rect 13916 19852 14196 19854
rect 12908 19348 12964 19358
rect 12908 19254 12964 19292
rect 10108 19182 10110 19234
rect 10162 19182 10164 19234
rect 10108 19170 10164 19182
rect 13804 19236 13860 19246
rect 13916 19236 13972 19852
rect 14140 19842 14196 19852
rect 13804 19234 13972 19236
rect 13804 19182 13806 19234
rect 13858 19182 13972 19234
rect 13804 19180 13972 19182
rect 13804 19170 13860 19180
rect 10780 19124 10836 19134
rect 10780 19030 10836 19068
rect 13468 19124 13524 19134
rect 13468 19030 13524 19068
rect 14252 19010 14308 20076
rect 14364 20018 14420 20750
rect 14812 20804 14868 20814
rect 14812 20710 14868 20748
rect 15036 20132 15204 20188
rect 14364 19966 14366 20018
rect 14418 19966 14420 20018
rect 14364 19348 14420 19966
rect 14364 19282 14420 19292
rect 14812 20018 14868 20030
rect 14812 19966 14814 20018
rect 14866 19966 14868 20018
rect 14812 19908 14868 19966
rect 14812 19236 14868 19852
rect 14812 19142 14868 19180
rect 14252 18958 14254 19010
rect 14306 18958 14308 19010
rect 13132 18338 13188 18350
rect 13132 18286 13134 18338
rect 13186 18286 13188 18338
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 4284 16884 4340 16894
rect 4284 16790 4340 16828
rect 12236 16884 12292 16894
rect 1932 16658 1988 16670
rect 1932 16606 1934 16658
rect 1986 16606 1988 16658
rect 1932 16212 1988 16606
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 1932 16146 1988 16156
rect 12236 16100 12292 16828
rect 12908 16884 12964 16894
rect 13132 16884 13188 18286
rect 13692 16996 13748 17006
rect 12964 16828 13188 16884
rect 13580 16940 13692 16996
rect 13580 16882 13636 16940
rect 13692 16930 13748 16940
rect 13580 16830 13582 16882
rect 13634 16830 13636 16882
rect 12908 16790 12964 16828
rect 13580 16818 13636 16830
rect 14252 16884 14308 18958
rect 15036 19010 15092 20132
rect 15148 19908 15204 20132
rect 15260 20132 15316 22988
rect 15372 20580 15428 23100
rect 15932 22482 15988 23324
rect 16828 23154 16884 23166
rect 16828 23102 16830 23154
rect 16882 23102 16884 23154
rect 16044 23042 16100 23054
rect 16044 22990 16046 23042
rect 16098 22990 16100 23042
rect 16044 22594 16100 22990
rect 16828 23044 16884 23102
rect 17052 23044 17108 25116
rect 17164 23940 17220 25228
rect 17276 25218 17332 25228
rect 17164 23874 17220 23884
rect 17388 23492 17444 28028
rect 17500 27858 17556 27870
rect 17500 27806 17502 27858
rect 17554 27806 17556 27858
rect 17500 26180 17556 27806
rect 18172 27748 18228 27758
rect 18172 27654 18228 27692
rect 19292 27186 19348 28252
rect 19292 27134 19294 27186
rect 19346 27134 19348 27186
rect 19292 27122 19348 27134
rect 19404 26964 19460 28476
rect 19516 28532 19572 37212
rect 19740 37202 19796 37212
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 21420 31948 21476 37998
rect 23548 36708 23604 41200
rect 25564 38276 25620 38286
rect 25564 38182 25620 38220
rect 24556 38052 24612 38062
rect 23548 36642 23604 36652
rect 23772 38050 24612 38052
rect 23772 37998 24558 38050
rect 24610 37998 24612 38050
rect 23772 37996 24612 37998
rect 20188 31892 21476 31948
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 19516 28438 19572 28476
rect 19740 28420 19796 28430
rect 19628 28418 19796 28420
rect 19628 28366 19742 28418
rect 19794 28366 19796 28418
rect 19628 28364 19796 28366
rect 19516 27748 19572 27758
rect 19516 27074 19572 27692
rect 19516 27022 19518 27074
rect 19570 27022 19572 27074
rect 19516 27010 19572 27022
rect 19628 27076 19684 28364
rect 19740 28354 19796 28364
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 19852 27076 19908 27086
rect 19628 27074 19908 27076
rect 19628 27022 19854 27074
rect 19906 27022 19908 27074
rect 19628 27020 19908 27022
rect 19852 27010 19908 27020
rect 19292 26908 19460 26964
rect 19628 26908 19796 26964
rect 18620 26852 19348 26908
rect 17556 26124 17668 26180
rect 17500 26086 17556 26124
rect 17500 25394 17556 25406
rect 17500 25342 17502 25394
rect 17554 25342 17556 25394
rect 17500 23604 17556 25342
rect 17612 25172 17668 26124
rect 18620 25396 18676 26852
rect 19516 26180 19572 26190
rect 19516 26086 19572 26124
rect 18620 25302 18676 25340
rect 17612 25106 17668 25116
rect 17836 25284 17892 25294
rect 17836 23938 17892 25228
rect 18284 25284 18340 25294
rect 18284 25190 18340 25228
rect 19628 24948 19684 26908
rect 19740 26850 19796 26908
rect 19740 26798 19742 26850
rect 19794 26798 19796 26850
rect 19740 26786 19796 26798
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 20188 26178 20244 31892
rect 20300 28532 20356 28542
rect 20300 27746 20356 28476
rect 20300 27694 20302 27746
rect 20354 27694 20356 27746
rect 20300 27682 20356 27694
rect 20972 27858 21028 27870
rect 20972 27806 20974 27858
rect 21026 27806 21028 27858
rect 20188 26126 20190 26178
rect 20242 26126 20244 26178
rect 20188 25620 20244 26126
rect 20524 26850 20580 26862
rect 20524 26798 20526 26850
rect 20578 26798 20580 26850
rect 20524 26180 20580 26798
rect 20524 26114 20580 26124
rect 20748 26852 20804 26862
rect 20188 25554 20244 25564
rect 20188 25284 20244 25294
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 19404 24892 19684 24948
rect 20188 24946 20244 25228
rect 20188 24894 20190 24946
rect 20242 24894 20244 24946
rect 17836 23886 17838 23938
rect 17890 23886 17892 23938
rect 17724 23828 17780 23838
rect 17500 23538 17556 23548
rect 17612 23772 17724 23828
rect 16884 22988 17108 23044
rect 16828 22978 16884 22988
rect 16044 22542 16046 22594
rect 16098 22542 16100 22594
rect 16044 22530 16100 22542
rect 15932 22430 15934 22482
rect 15986 22430 15988 22482
rect 15932 22418 15988 22430
rect 17052 22482 17108 22988
rect 17052 22430 17054 22482
rect 17106 22430 17108 22482
rect 16380 22148 16436 22158
rect 16380 20804 16436 22092
rect 17052 21700 17108 22430
rect 17276 23436 17444 23492
rect 17276 22484 17332 23436
rect 17388 23268 17444 23278
rect 17388 23174 17444 23212
rect 17612 23266 17668 23772
rect 17724 23762 17780 23772
rect 17724 23380 17780 23390
rect 17724 23286 17780 23324
rect 17612 23214 17614 23266
rect 17666 23214 17668 23266
rect 17612 23202 17668 23214
rect 17836 23156 17892 23886
rect 18284 24836 18340 24846
rect 18172 23828 18228 23838
rect 18172 23734 18228 23772
rect 17724 23100 17892 23156
rect 18284 23154 18340 24780
rect 18508 23940 18564 23950
rect 18564 23884 18900 23940
rect 18508 23846 18564 23884
rect 18284 23102 18286 23154
rect 18338 23102 18340 23154
rect 17724 22594 17780 23100
rect 18060 23044 18116 23054
rect 18060 22950 18116 22988
rect 17836 22932 17892 22942
rect 17836 22838 17892 22876
rect 17724 22542 17726 22594
rect 17778 22542 17780 22594
rect 17724 22530 17780 22542
rect 17276 22428 17444 22484
rect 17052 21634 17108 21644
rect 17276 22260 17332 22270
rect 15372 20486 15428 20524
rect 15484 20690 15540 20702
rect 15484 20638 15486 20690
rect 15538 20638 15540 20690
rect 15260 20066 15316 20076
rect 15484 19908 15540 20638
rect 16268 20132 16324 20142
rect 16380 20132 16436 20748
rect 16268 20130 16436 20132
rect 16268 20078 16270 20130
rect 16322 20078 16436 20130
rect 16268 20076 16436 20078
rect 16604 21028 16660 21038
rect 16268 20066 16324 20076
rect 16604 19908 16660 20972
rect 17164 21028 17220 21038
rect 16940 20802 16996 20814
rect 16940 20750 16942 20802
rect 16994 20750 16996 20802
rect 16716 19908 16772 19918
rect 15148 19852 15540 19908
rect 16380 19906 16772 19908
rect 16380 19854 16718 19906
rect 16770 19854 16772 19906
rect 16380 19852 16772 19854
rect 15484 19236 15540 19246
rect 15484 19142 15540 19180
rect 16044 19234 16100 19246
rect 16044 19182 16046 19234
rect 16098 19182 16100 19234
rect 15036 18958 15038 19010
rect 15090 18958 15092 19010
rect 15036 18676 15092 18958
rect 16044 19012 16100 19182
rect 16044 18946 16100 18956
rect 16268 18676 16324 18686
rect 15036 18610 15092 18620
rect 16156 18620 16268 18676
rect 14812 18004 14868 18014
rect 16156 18004 16212 18620
rect 16268 18582 16324 18620
rect 16380 18562 16436 19852
rect 16716 19842 16772 19852
rect 16716 19010 16772 19022
rect 16716 18958 16718 19010
rect 16770 18958 16772 19010
rect 16716 18676 16772 18958
rect 16940 19012 16996 20750
rect 17164 20802 17220 20972
rect 17276 20914 17332 22204
rect 17276 20862 17278 20914
rect 17330 20862 17332 20914
rect 17276 20850 17332 20862
rect 17164 20750 17166 20802
rect 17218 20750 17220 20802
rect 17164 20738 17220 20750
rect 17388 19460 17444 22428
rect 18060 22258 18116 22270
rect 18060 22206 18062 22258
rect 18114 22206 18116 22258
rect 17836 22146 17892 22158
rect 17836 22094 17838 22146
rect 17890 22094 17892 22146
rect 17724 21700 17780 21710
rect 17724 21606 17780 21644
rect 17276 19404 17388 19460
rect 17052 19236 17108 19246
rect 17052 19122 17108 19180
rect 17052 19070 17054 19122
rect 17106 19070 17108 19122
rect 17052 19058 17108 19070
rect 16940 18946 16996 18956
rect 16716 18610 16772 18620
rect 16380 18510 16382 18562
rect 16434 18510 16436 18562
rect 16380 18498 16436 18510
rect 16268 18228 16324 18238
rect 17052 18228 17108 18238
rect 16324 18172 16436 18228
rect 16268 18134 16324 18172
rect 16156 17948 16324 18004
rect 14812 17554 14868 17948
rect 16156 17780 16212 17790
rect 15932 17778 16212 17780
rect 15932 17726 16158 17778
rect 16210 17726 16212 17778
rect 15932 17724 16212 17726
rect 14812 17502 14814 17554
rect 14866 17502 14868 17554
rect 14812 17490 14868 17502
rect 14924 17556 14980 17566
rect 14924 17462 14980 17500
rect 14588 17442 14644 17454
rect 14588 17390 14590 17442
rect 14642 17390 14644 17442
rect 14588 16996 14644 17390
rect 14588 16930 14644 16940
rect 14252 16818 14308 16828
rect 15708 16772 15764 16782
rect 15708 16678 15764 16716
rect 15932 16322 15988 17724
rect 16156 17714 16212 17724
rect 16268 17554 16324 17948
rect 16268 17502 16270 17554
rect 16322 17502 16324 17554
rect 16268 17490 16324 17502
rect 15932 16270 15934 16322
rect 15986 16270 15988 16322
rect 15932 16258 15988 16270
rect 16156 16884 16212 16894
rect 16156 16770 16212 16828
rect 16156 16718 16158 16770
rect 16210 16718 16212 16770
rect 12236 15202 12292 16044
rect 15820 16100 15876 16110
rect 15820 16006 15876 16044
rect 14476 15988 14532 15998
rect 14476 15894 14532 15932
rect 14252 15874 14308 15886
rect 14252 15822 14254 15874
rect 14306 15822 14308 15874
rect 14252 15428 14308 15822
rect 14252 15362 14308 15372
rect 14364 15874 14420 15886
rect 14364 15822 14366 15874
rect 14418 15822 14420 15874
rect 14364 15426 14420 15822
rect 14364 15374 14366 15426
rect 14418 15374 14420 15426
rect 14364 15362 14420 15374
rect 12236 15150 12238 15202
rect 12290 15150 12292 15202
rect 12236 15138 12292 15150
rect 15148 15314 15204 15326
rect 15148 15262 15150 15314
rect 15202 15262 15204 15314
rect 15148 15204 15204 15262
rect 15596 15204 15652 15214
rect 15148 15202 15652 15204
rect 15148 15150 15598 15202
rect 15650 15150 15652 15202
rect 15148 15148 15652 15150
rect 16156 15148 16212 16718
rect 16380 16884 16436 18172
rect 17052 17666 17108 18172
rect 17052 17614 17054 17666
rect 17106 17614 17108 17666
rect 17052 17602 17108 17614
rect 16492 17554 16548 17566
rect 16492 17502 16494 17554
rect 16546 17502 16548 17554
rect 16492 17108 16548 17502
rect 16716 17556 16772 17566
rect 16716 17462 16772 17500
rect 16940 17444 16996 17454
rect 16940 17350 16996 17388
rect 16492 17042 16548 17052
rect 16268 16660 16324 16670
rect 16268 15986 16324 16604
rect 16380 16100 16436 16828
rect 16492 16100 16548 16110
rect 16380 16098 16548 16100
rect 16380 16046 16494 16098
rect 16546 16046 16548 16098
rect 16380 16044 16548 16046
rect 16492 16034 16548 16044
rect 16828 16098 16884 16110
rect 16828 16046 16830 16098
rect 16882 16046 16884 16098
rect 16268 15934 16270 15986
rect 16322 15934 16324 15986
rect 16268 15922 16324 15934
rect 16604 15988 16660 15998
rect 16604 15894 16660 15932
rect 16828 15876 16884 16046
rect 16828 15810 16884 15820
rect 17276 15652 17332 19404
rect 17388 19394 17444 19404
rect 17612 20916 17668 20926
rect 17836 20916 17892 22094
rect 17612 18450 17668 20860
rect 17724 20860 17892 20916
rect 18060 20916 18116 22206
rect 17724 20802 17780 20860
rect 18060 20850 18116 20860
rect 17724 20750 17726 20802
rect 17778 20750 17780 20802
rect 17724 20468 17780 20750
rect 17836 20692 17892 20702
rect 17836 20598 17892 20636
rect 17948 20692 18004 20702
rect 17948 20690 18116 20692
rect 17948 20638 17950 20690
rect 18002 20638 18116 20690
rect 17948 20636 18116 20638
rect 17948 20626 18004 20636
rect 17724 20412 18004 20468
rect 17724 19458 17780 20412
rect 17948 20242 18004 20412
rect 17948 20190 17950 20242
rect 18002 20190 18004 20242
rect 17948 20178 18004 20190
rect 17724 19406 17726 19458
rect 17778 19406 17780 19458
rect 17724 19394 17780 19406
rect 17612 18398 17614 18450
rect 17666 18398 17668 18450
rect 17500 18338 17556 18350
rect 17500 18286 17502 18338
rect 17554 18286 17556 18338
rect 17388 17108 17444 17118
rect 17388 17014 17444 17052
rect 17500 16772 17556 18286
rect 17612 17668 17668 18398
rect 17836 19122 17892 19134
rect 17836 19070 17838 19122
rect 17890 19070 17892 19122
rect 17836 18452 17892 19070
rect 17948 19124 18004 19134
rect 18060 19124 18116 20636
rect 18284 19236 18340 23102
rect 18396 23604 18452 23614
rect 18396 22260 18452 23548
rect 18396 22166 18452 22204
rect 18844 23154 18900 23884
rect 19404 23716 19460 24892
rect 20188 24882 20244 24894
rect 19964 24836 20020 24846
rect 19964 24742 20020 24780
rect 19852 24722 19908 24734
rect 19852 24670 19854 24722
rect 19906 24670 19908 24722
rect 19628 23938 19684 23950
rect 19628 23886 19630 23938
rect 19682 23886 19684 23938
rect 19404 23660 19572 23716
rect 19516 23378 19572 23660
rect 19628 23604 19684 23886
rect 19852 23940 19908 24670
rect 20748 24050 20804 26796
rect 20972 26404 21028 27806
rect 22540 27860 22596 27870
rect 21644 27746 21700 27758
rect 21644 27694 21646 27746
rect 21698 27694 21700 27746
rect 21644 27186 21700 27694
rect 21644 27134 21646 27186
rect 21698 27134 21700 27186
rect 21644 27122 21700 27134
rect 22540 27186 22596 27804
rect 23772 27860 23828 37996
rect 24556 37986 24612 37996
rect 26236 37940 26292 41200
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 26236 37874 26292 37884
rect 27468 37940 27524 37950
rect 27468 37846 27524 37884
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 24780 36708 24836 36718
rect 24780 36614 24836 36652
rect 24108 36482 24164 36494
rect 24108 36430 24110 36482
rect 24162 36430 24164 36482
rect 24108 28082 24164 36430
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 24108 28030 24110 28082
rect 24162 28030 24164 28082
rect 24108 28018 24164 28030
rect 23772 27746 23828 27804
rect 24444 27860 24500 27870
rect 24444 27766 24500 27804
rect 23772 27694 23774 27746
rect 23826 27694 23828 27746
rect 23772 27682 23828 27694
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 22540 27134 22542 27186
rect 22594 27134 22596 27186
rect 22540 27122 22596 27134
rect 20972 26338 21028 26348
rect 21420 27076 21476 27086
rect 20748 23998 20750 24050
rect 20802 23998 20804 24050
rect 20748 23986 20804 23998
rect 21308 25394 21364 25406
rect 21308 25342 21310 25394
rect 21362 25342 21364 25394
rect 19852 23874 19908 23884
rect 20300 23938 20356 23950
rect 20300 23886 20302 23938
rect 20354 23886 20356 23938
rect 19964 23828 20020 23838
rect 20020 23772 20132 23828
rect 19964 23734 20020 23772
rect 20076 23716 20132 23772
rect 20076 23660 20244 23716
rect 19628 23538 19684 23548
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 20188 23380 20244 23660
rect 19516 23326 19518 23378
rect 19570 23326 19572 23378
rect 19516 23314 19572 23326
rect 19628 23324 20020 23380
rect 19404 23268 19460 23278
rect 19404 23174 19460 23212
rect 18844 23102 18846 23154
rect 18898 23102 18900 23154
rect 18508 22146 18564 22158
rect 18508 22094 18510 22146
rect 18562 22094 18564 22146
rect 18396 21924 18452 21934
rect 18396 21026 18452 21868
rect 18396 20974 18398 21026
rect 18450 20974 18452 21026
rect 18396 20962 18452 20974
rect 18508 20804 18564 22094
rect 18508 20738 18564 20748
rect 18732 22146 18788 22158
rect 18732 22094 18734 22146
rect 18786 22094 18788 22146
rect 18508 19908 18564 19918
rect 18508 19814 18564 19852
rect 18284 19170 18340 19180
rect 18004 19068 18116 19124
rect 17948 19058 18004 19068
rect 17948 18452 18004 18462
rect 17836 18450 18004 18452
rect 17836 18398 17950 18450
rect 18002 18398 18004 18450
rect 17836 18396 18004 18398
rect 17612 17602 17668 17612
rect 17724 16772 17780 16782
rect 17500 16716 17724 16772
rect 17724 16678 17780 16716
rect 17948 16770 18004 18396
rect 18508 18452 18564 18462
rect 18508 18358 18564 18396
rect 18508 17780 18564 17790
rect 18508 17554 18564 17724
rect 18508 17502 18510 17554
rect 18562 17502 18564 17554
rect 18508 17490 18564 17502
rect 17948 16718 17950 16770
rect 18002 16718 18004 16770
rect 17948 16548 18004 16718
rect 18172 17442 18228 17454
rect 18172 17390 18174 17442
rect 18226 17390 18228 17442
rect 18172 16772 18228 17390
rect 18732 16996 18788 22094
rect 18844 21026 18900 23102
rect 19180 23156 19236 23166
rect 19180 23154 19348 23156
rect 19180 23102 19182 23154
rect 19234 23102 19348 23154
rect 19180 23100 19348 23102
rect 19180 23090 19236 23100
rect 19292 23044 19348 23100
rect 19628 23044 19684 23324
rect 19292 22988 19684 23044
rect 19740 23154 19796 23166
rect 19740 23102 19742 23154
rect 19794 23102 19796 23154
rect 18844 20974 18846 21026
rect 18898 20974 18900 21026
rect 18844 20962 18900 20974
rect 18956 22932 19012 22942
rect 18956 22146 19012 22876
rect 18956 22094 18958 22146
rect 19010 22094 19012 22146
rect 18844 20692 18900 20702
rect 18844 19908 18900 20636
rect 18844 18450 18900 19852
rect 18844 18398 18846 18450
rect 18898 18398 18900 18450
rect 18844 18386 18900 18398
rect 18844 17668 18900 17678
rect 18844 17574 18900 17612
rect 18732 16930 18788 16940
rect 18172 16706 18228 16716
rect 18284 16884 18340 16894
rect 17500 16492 18004 16548
rect 17276 15586 17332 15596
rect 17388 15876 17444 15886
rect 17500 15876 17556 16492
rect 17388 15874 17556 15876
rect 17388 15822 17390 15874
rect 17442 15822 17556 15874
rect 17388 15820 17556 15822
rect 17612 16380 18228 16436
rect 15148 15092 15204 15148
rect 14812 15036 15204 15092
rect 15596 15092 16212 15148
rect 17276 15314 17332 15326
rect 17276 15262 17278 15314
rect 17330 15262 17332 15314
rect 17276 15204 17332 15262
rect 17276 15138 17332 15148
rect 17388 15148 17444 15820
rect 17500 15540 17556 15578
rect 17500 15474 17556 15484
rect 17612 15426 17668 16380
rect 18172 16322 18228 16380
rect 18172 16270 18174 16322
rect 18226 16270 18228 16322
rect 18172 16258 18228 16270
rect 18060 16100 18116 16110
rect 18284 16100 18340 16828
rect 18060 16098 18340 16100
rect 18060 16046 18062 16098
rect 18114 16046 18340 16098
rect 18060 16044 18340 16046
rect 18060 16034 18116 16044
rect 17724 15876 17780 15886
rect 17724 15782 17780 15820
rect 18172 15874 18228 15886
rect 18172 15822 18174 15874
rect 18226 15822 18228 15874
rect 17612 15374 17614 15426
rect 17666 15374 17668 15426
rect 17612 15362 17668 15374
rect 18172 15316 18228 15822
rect 18172 15250 18228 15260
rect 18956 15204 19012 22094
rect 19180 22372 19236 22382
rect 19740 22372 19796 23102
rect 19180 22370 19796 22372
rect 19180 22318 19182 22370
rect 19234 22318 19796 22370
rect 19180 22316 19796 22318
rect 19852 22370 19908 22382
rect 19852 22318 19854 22370
rect 19906 22318 19908 22370
rect 19180 21924 19236 22316
rect 19852 22148 19908 22318
rect 19964 22260 20020 23324
rect 20076 23324 20244 23380
rect 20076 23154 20132 23324
rect 20076 23102 20078 23154
rect 20130 23102 20132 23154
rect 20076 23090 20132 23102
rect 20188 23156 20244 23166
rect 20300 23156 20356 23886
rect 20636 23826 20692 23838
rect 20636 23774 20638 23826
rect 20690 23774 20692 23826
rect 20412 23716 20468 23726
rect 20412 23378 20468 23660
rect 20412 23326 20414 23378
rect 20466 23326 20468 23378
rect 20412 23314 20468 23326
rect 20244 23100 20356 23156
rect 20524 23156 20580 23166
rect 20636 23156 20692 23774
rect 21308 23716 21364 25342
rect 21308 23650 21364 23660
rect 21420 23380 21476 27020
rect 21980 27074 22036 27086
rect 21980 27022 21982 27074
rect 22034 27022 22036 27074
rect 21756 26964 21812 26974
rect 21756 26870 21812 26908
rect 21532 26852 21588 26862
rect 21532 26758 21588 26796
rect 21868 26180 21924 26190
rect 21868 25618 21924 26124
rect 21868 25566 21870 25618
rect 21922 25566 21924 25618
rect 21868 25554 21924 25566
rect 21868 25396 21924 25406
rect 21980 25396 22036 27022
rect 22428 26964 22484 26974
rect 22428 26870 22484 26908
rect 23996 26850 24052 26862
rect 23996 26798 23998 26850
rect 24050 26798 24052 26850
rect 22988 26404 23044 26414
rect 22988 26290 23044 26348
rect 23548 26404 23604 26414
rect 23548 26310 23604 26348
rect 23996 26404 24052 26798
rect 23996 26338 24052 26348
rect 25228 26404 25284 26414
rect 22988 26238 22990 26290
rect 23042 26238 23044 26290
rect 22316 26180 22372 26190
rect 22316 26086 22372 26124
rect 22428 25620 22484 25630
rect 22428 25526 22484 25564
rect 21924 25340 22036 25396
rect 21868 25302 21924 25340
rect 21532 25284 21588 25294
rect 21532 25190 21588 25228
rect 21756 25284 21812 25294
rect 21756 25190 21812 25228
rect 22316 25284 22372 25294
rect 22316 25190 22372 25228
rect 22876 23940 22932 23950
rect 22988 23940 23044 26238
rect 24108 24836 24164 24846
rect 24108 24742 24164 24780
rect 22876 23938 23044 23940
rect 22876 23886 22878 23938
rect 22930 23886 23044 23938
rect 22876 23884 23044 23886
rect 23996 24722 24052 24734
rect 23996 24670 23998 24722
rect 24050 24670 24052 24722
rect 22876 23874 22932 23884
rect 23548 23828 23604 23838
rect 23996 23828 24052 24670
rect 23548 23826 23716 23828
rect 23548 23774 23550 23826
rect 23602 23774 23716 23826
rect 23548 23772 23716 23774
rect 23548 23762 23604 23772
rect 21308 23324 21476 23380
rect 21644 23380 21700 23390
rect 21196 23266 21252 23278
rect 21196 23214 21198 23266
rect 21250 23214 21252 23266
rect 20972 23156 21028 23166
rect 20636 23154 21028 23156
rect 20636 23102 20974 23154
rect 21026 23102 21028 23154
rect 20636 23100 21028 23102
rect 20188 23062 20244 23100
rect 20524 23062 20580 23100
rect 20412 23044 20468 23054
rect 20412 22594 20468 22988
rect 20412 22542 20414 22594
rect 20466 22542 20468 22594
rect 20412 22530 20468 22542
rect 20412 22370 20468 22382
rect 20412 22318 20414 22370
rect 20466 22318 20468 22370
rect 20076 22260 20132 22270
rect 19964 22258 20132 22260
rect 19964 22206 20078 22258
rect 20130 22206 20132 22258
rect 19964 22204 20132 22206
rect 20076 22148 20132 22204
rect 20076 22092 20244 22148
rect 19852 22082 19908 22092
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 19180 21858 19236 21868
rect 20188 21812 20244 22092
rect 20076 21756 20244 21812
rect 19852 20916 19908 20926
rect 19292 20804 19348 20814
rect 19516 20804 19572 20814
rect 19628 20804 19684 20814
rect 19292 20802 19460 20804
rect 19292 20750 19294 20802
rect 19346 20750 19460 20802
rect 19292 20748 19460 20750
rect 19292 20738 19348 20748
rect 19068 20020 19124 20030
rect 19068 19926 19124 19964
rect 19292 19234 19348 19246
rect 19292 19182 19294 19234
rect 19346 19182 19348 19234
rect 19292 19012 19348 19182
rect 19292 18946 19348 18956
rect 19404 18452 19460 20748
rect 19516 20802 19628 20804
rect 19516 20750 19518 20802
rect 19570 20750 19628 20802
rect 19516 20748 19628 20750
rect 19516 20738 19572 20748
rect 19516 20020 19572 20030
rect 19516 19926 19572 19964
rect 19404 18386 19460 18396
rect 19516 19010 19572 19022
rect 19516 18958 19518 19010
rect 19570 18958 19572 19010
rect 19516 17668 19572 18958
rect 19628 18562 19684 20748
rect 19852 20802 19908 20860
rect 19852 20750 19854 20802
rect 19906 20750 19908 20802
rect 19852 20738 19908 20750
rect 20076 20580 20132 21756
rect 20300 20914 20356 20926
rect 20300 20862 20302 20914
rect 20354 20862 20356 20914
rect 20300 20804 20356 20862
rect 20300 20738 20356 20748
rect 20412 20692 20468 22318
rect 20748 22258 20804 22270
rect 20748 22206 20750 22258
rect 20802 22206 20804 22258
rect 20412 20626 20468 20636
rect 20524 22148 20580 22158
rect 20076 20524 20244 20580
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 20188 20020 20244 20524
rect 20188 19954 20244 19964
rect 19852 19348 19908 19358
rect 19852 19254 19908 19292
rect 20188 19348 20244 19358
rect 20076 19234 20132 19246
rect 20076 19182 20078 19234
rect 20130 19182 20132 19234
rect 20076 19124 20132 19182
rect 20076 19058 20132 19068
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 19628 18510 19630 18562
rect 19682 18510 19684 18562
rect 19628 18498 19684 18510
rect 19516 17602 19572 17612
rect 19852 17780 19908 17790
rect 19852 17666 19908 17724
rect 19852 17614 19854 17666
rect 19906 17614 19908 17666
rect 19852 17602 19908 17614
rect 20188 17554 20244 19292
rect 20524 19236 20580 22092
rect 20748 21812 20804 22206
rect 20748 21746 20804 21756
rect 20972 20804 21028 23100
rect 21196 23156 21252 23214
rect 21196 23090 21252 23100
rect 21308 22036 21364 23324
rect 21644 23286 21700 23324
rect 22316 23380 22372 23390
rect 21420 23154 21476 23166
rect 21420 23102 21422 23154
rect 21474 23102 21476 23154
rect 21420 22596 21476 23102
rect 21420 22530 21476 22540
rect 21756 23156 21812 23166
rect 21420 22372 21476 22382
rect 21420 22370 21588 22372
rect 21420 22318 21422 22370
rect 21474 22318 21588 22370
rect 21420 22316 21588 22318
rect 21420 22306 21476 22316
rect 21308 21980 21476 22036
rect 21308 21812 21364 21822
rect 21196 20804 21252 20814
rect 20972 20802 21252 20804
rect 20972 20750 21198 20802
rect 21250 20750 21252 20802
rect 20972 20748 21252 20750
rect 21196 20738 21252 20748
rect 21196 19460 21252 19470
rect 21196 19366 21252 19404
rect 20300 19180 20580 19236
rect 21308 19348 21364 21756
rect 21308 19234 21364 19292
rect 21308 19182 21310 19234
rect 21362 19182 21364 19234
rect 20300 18340 20356 19180
rect 21308 19170 21364 19182
rect 20412 19012 20468 19022
rect 20412 19010 20692 19012
rect 20412 18958 20414 19010
rect 20466 18958 20692 19010
rect 20412 18956 20692 18958
rect 20412 18946 20468 18956
rect 20524 18788 20580 18798
rect 20412 18732 20524 18788
rect 20412 18562 20468 18732
rect 20524 18722 20580 18732
rect 20412 18510 20414 18562
rect 20466 18510 20468 18562
rect 20412 18498 20468 18510
rect 20524 18450 20580 18462
rect 20524 18398 20526 18450
rect 20578 18398 20580 18450
rect 20524 18340 20580 18398
rect 20300 18284 20580 18340
rect 20412 17892 20468 17902
rect 20188 17502 20190 17554
rect 20242 17502 20244 17554
rect 20188 17490 20244 17502
rect 20300 17668 20356 17678
rect 19180 17444 19236 17454
rect 17388 15092 17556 15148
rect 18956 15138 19012 15148
rect 19068 17442 19236 17444
rect 19068 17390 19182 17442
rect 19234 17390 19236 17442
rect 19068 17388 19236 17390
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 14812 14530 14868 15036
rect 15484 14980 15540 14990
rect 15484 14642 15540 14924
rect 15484 14590 15486 14642
rect 15538 14590 15540 14642
rect 15484 14578 15540 14590
rect 14812 14478 14814 14530
rect 14866 14478 14868 14530
rect 14812 14466 14868 14478
rect 15596 14308 15652 15092
rect 17500 14644 17556 15092
rect 19068 14868 19124 17388
rect 19180 17378 19236 17388
rect 19516 17444 19572 17454
rect 19516 17350 19572 17388
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 20300 16884 20356 17612
rect 19964 16828 20356 16884
rect 19964 16770 20020 16828
rect 19964 16718 19966 16770
rect 20018 16718 20020 16770
rect 19964 16706 20020 16718
rect 19852 16658 19908 16670
rect 19852 16606 19854 16658
rect 19906 16606 19908 16658
rect 19852 16100 19908 16606
rect 20188 16658 20244 16670
rect 20188 16606 20190 16658
rect 20242 16606 20244 16658
rect 20188 16436 20244 16606
rect 20300 16660 20356 16670
rect 20300 16566 20356 16604
rect 20412 16436 20468 17836
rect 20524 17780 20580 17790
rect 20524 17666 20580 17724
rect 20524 17614 20526 17666
rect 20578 17614 20580 17666
rect 20524 17602 20580 17614
rect 20188 16380 20468 16436
rect 20524 16996 20580 17006
rect 20524 16324 20580 16940
rect 19852 16034 19908 16044
rect 20188 16268 20580 16324
rect 20188 16098 20244 16268
rect 20188 16046 20190 16098
rect 20242 16046 20244 16098
rect 20188 16034 20244 16046
rect 20300 16100 20356 16110
rect 19852 15876 19908 15886
rect 19180 15874 19908 15876
rect 19180 15822 19854 15874
rect 19906 15822 19908 15874
rect 19180 15820 19908 15822
rect 19180 15538 19236 15820
rect 19180 15486 19182 15538
rect 19234 15486 19236 15538
rect 19180 15474 19236 15486
rect 19628 15428 19684 15820
rect 19852 15810 19908 15820
rect 20076 15876 20132 15914
rect 20076 15810 20132 15820
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 19628 15372 20020 15428
rect 19404 15314 19460 15326
rect 19404 15262 19406 15314
rect 19458 15262 19460 15314
rect 19068 14802 19124 14812
rect 19292 15202 19348 15214
rect 19292 15150 19294 15202
rect 19346 15150 19348 15202
rect 17612 14644 17668 14654
rect 19292 14644 19348 15150
rect 17500 14642 17668 14644
rect 17500 14590 17614 14642
rect 17666 14590 17668 14642
rect 17500 14588 17668 14590
rect 17612 14578 17668 14588
rect 18732 14588 19348 14644
rect 19404 14642 19460 15262
rect 19516 15316 19572 15326
rect 19516 15222 19572 15260
rect 19852 15204 19908 15242
rect 19852 15138 19908 15148
rect 19964 14754 20020 15372
rect 20076 15316 20132 15326
rect 20300 15316 20356 16044
rect 20076 15314 20356 15316
rect 20076 15262 20078 15314
rect 20130 15262 20356 15314
rect 20076 15260 20356 15262
rect 20076 15250 20132 15260
rect 19964 14702 19966 14754
rect 20018 14702 20020 14754
rect 19964 14690 20020 14702
rect 20188 15092 20244 15102
rect 19404 14590 19406 14642
rect 19458 14590 19460 14642
rect 15596 14242 15652 14252
rect 18060 14308 18116 14318
rect 18060 13748 18116 14252
rect 18620 13748 18676 13758
rect 17948 13746 18676 13748
rect 17948 13694 18622 13746
rect 18674 13694 18676 13746
rect 17948 13692 18676 13694
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 17948 12962 18004 13692
rect 18620 13524 18676 13692
rect 18620 13458 18676 13468
rect 18620 13076 18676 13086
rect 18732 13076 18788 14588
rect 19404 14578 19460 14590
rect 19292 14420 19348 14430
rect 19292 14326 19348 14364
rect 19516 14306 19572 14318
rect 19516 14254 19518 14306
rect 19570 14254 19572 14306
rect 19292 13860 19348 13870
rect 19292 13766 19348 13804
rect 18620 13074 18788 13076
rect 18620 13022 18622 13074
rect 18674 13022 18788 13074
rect 18620 13020 18788 13022
rect 19516 13076 19572 14254
rect 20188 14308 20244 15036
rect 20300 14532 20356 14542
rect 20300 14438 20356 14476
rect 20636 14530 20692 18956
rect 21420 18340 21476 21980
rect 21532 20802 21588 22316
rect 21756 22260 21812 23100
rect 21756 22194 21812 22204
rect 22092 23042 22148 23054
rect 22092 22990 22094 23042
rect 22146 22990 22148 23042
rect 21532 20750 21534 20802
rect 21586 20750 21588 20802
rect 21532 20692 21588 20750
rect 21532 20626 21588 20636
rect 21644 22146 21700 22158
rect 21980 22148 22036 22158
rect 21644 22094 21646 22146
rect 21698 22094 21700 22146
rect 21644 20356 21700 22094
rect 21532 20300 21700 20356
rect 21868 22146 22036 22148
rect 21868 22094 21982 22146
rect 22034 22094 22036 22146
rect 21868 22092 22036 22094
rect 21532 19124 21588 20300
rect 21868 20188 21924 22092
rect 21980 22082 22036 22092
rect 22092 22148 22148 22990
rect 22092 22082 22148 22092
rect 22204 22930 22260 22942
rect 22204 22878 22206 22930
rect 22258 22878 22260 22930
rect 21980 20804 22036 20814
rect 22204 20804 22260 22878
rect 22316 22148 22372 23324
rect 23660 23378 23716 23772
rect 23996 23762 24052 23772
rect 24108 24498 24164 24510
rect 24108 24446 24110 24498
rect 24162 24446 24164 24498
rect 23660 23326 23662 23378
rect 23714 23326 23716 23378
rect 23660 23314 23716 23326
rect 23548 23154 23604 23166
rect 23548 23102 23550 23154
rect 23602 23102 23604 23154
rect 22540 23044 22596 23054
rect 22540 22370 22596 22988
rect 23548 22482 23604 23102
rect 23548 22430 23550 22482
rect 23602 22430 23604 22482
rect 23548 22418 23604 22430
rect 23772 23154 23828 23166
rect 23772 23102 23774 23154
rect 23826 23102 23828 23154
rect 23772 22484 23828 23102
rect 24108 23154 24164 24446
rect 24108 23102 24110 23154
rect 24162 23102 24164 23154
rect 24108 23090 24164 23102
rect 25228 23492 25284 26348
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 25676 24836 25732 24846
rect 25676 24052 25732 24780
rect 37660 24722 37716 24734
rect 37660 24670 37662 24722
rect 37714 24670 37716 24722
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 37660 24164 37716 24670
rect 40012 24498 40068 24510
rect 40012 24446 40014 24498
rect 40066 24446 40068 24498
rect 40012 24276 40068 24446
rect 40012 24210 40068 24220
rect 37660 24098 37716 24108
rect 25676 23958 25732 23996
rect 40012 24050 40068 24062
rect 40012 23998 40014 24050
rect 40066 23998 40068 24050
rect 37660 23938 37716 23950
rect 37660 23886 37662 23938
rect 37714 23886 37716 23938
rect 25228 23154 25284 23436
rect 26124 23714 26180 23726
rect 26124 23662 26126 23714
rect 26178 23662 26180 23714
rect 26124 23492 26180 23662
rect 28364 23714 28420 23726
rect 28364 23662 28366 23714
rect 28418 23662 28420 23714
rect 26180 23436 26404 23492
rect 26124 23426 26180 23436
rect 25228 23102 25230 23154
rect 25282 23102 25284 23154
rect 25228 23090 25284 23102
rect 26236 23268 26292 23278
rect 25116 23044 25172 23054
rect 25116 22594 25172 22988
rect 26012 23044 26068 23054
rect 26012 22950 26068 22988
rect 25116 22542 25118 22594
rect 25170 22542 25172 22594
rect 25116 22530 25172 22542
rect 23772 22428 24612 22484
rect 22540 22318 22542 22370
rect 22594 22318 22596 22370
rect 22540 22306 22596 22318
rect 22540 22148 22596 22158
rect 22316 22146 22540 22148
rect 22316 22094 22318 22146
rect 22370 22094 22540 22146
rect 22316 22092 22540 22094
rect 22316 22082 22372 22092
rect 21980 20802 22204 20804
rect 21980 20750 21982 20802
rect 22034 20750 22204 20802
rect 21980 20748 22204 20750
rect 21980 20738 22036 20748
rect 22204 20710 22260 20748
rect 22428 20802 22484 20814
rect 22428 20750 22430 20802
rect 22482 20750 22484 20802
rect 21532 19030 21588 19068
rect 21644 20132 21700 20142
rect 21308 18338 21476 18340
rect 21308 18286 21422 18338
rect 21474 18286 21476 18338
rect 21308 18284 21476 18286
rect 21308 18004 21364 18284
rect 21420 18274 21476 18284
rect 21308 17890 21364 17948
rect 21308 17838 21310 17890
rect 21362 17838 21364 17890
rect 21308 17826 21364 17838
rect 21644 17778 21700 20076
rect 21756 20132 21924 20188
rect 21756 18788 21812 20132
rect 21756 18722 21812 18732
rect 21868 20020 21924 20030
rect 21868 19234 21924 19964
rect 21868 19182 21870 19234
rect 21922 19182 21924 19234
rect 21868 17892 21924 19182
rect 21868 17798 21924 17836
rect 21644 17726 21646 17778
rect 21698 17726 21700 17778
rect 21644 17714 21700 17726
rect 22428 17780 22484 20750
rect 22540 19234 22596 22092
rect 22876 22146 22932 22158
rect 22876 22094 22878 22146
rect 22930 22094 22932 22146
rect 22652 21586 22708 21598
rect 22652 21534 22654 21586
rect 22706 21534 22708 21586
rect 22652 20914 22708 21534
rect 22652 20862 22654 20914
rect 22706 20862 22708 20914
rect 22652 20850 22708 20862
rect 22540 19182 22542 19234
rect 22594 19182 22596 19234
rect 22540 19170 22596 19182
rect 22764 19348 22820 19358
rect 22764 18564 22820 19292
rect 22876 19012 22932 22094
rect 23100 22148 23156 22158
rect 23100 22054 23156 22092
rect 23212 22146 23268 22158
rect 23436 22148 23492 22158
rect 23212 22094 23214 22146
rect 23266 22094 23268 22146
rect 22988 21812 23044 21822
rect 22988 21718 23044 21756
rect 23212 21812 23268 22094
rect 23212 21746 23268 21756
rect 23324 22146 23492 22148
rect 23324 22094 23438 22146
rect 23490 22094 23492 22146
rect 23324 22092 23492 22094
rect 23324 22036 23380 22092
rect 23436 22082 23492 22092
rect 23660 22148 23716 22158
rect 23660 22054 23716 22092
rect 23100 21700 23156 21710
rect 23100 21606 23156 21644
rect 23212 21586 23268 21598
rect 23212 21534 23214 21586
rect 23266 21534 23268 21586
rect 23212 21140 23268 21534
rect 22876 18946 22932 18956
rect 22988 21084 23268 21140
rect 22988 21028 23044 21084
rect 21532 17668 21588 17678
rect 21532 17574 21588 17612
rect 22092 17666 22148 17678
rect 22092 17614 22094 17666
rect 22146 17614 22148 17666
rect 21532 17220 21588 17230
rect 21532 16994 21588 17164
rect 21644 17108 21700 17118
rect 21644 17014 21700 17052
rect 21532 16942 21534 16994
rect 21586 16942 21588 16994
rect 21532 16930 21588 16942
rect 21868 16884 21924 16894
rect 21644 16660 21700 16670
rect 21644 16566 21700 16604
rect 21868 15092 21924 16828
rect 22092 16660 22148 17614
rect 22428 17668 22484 17724
rect 22652 18562 22820 18564
rect 22652 18510 22766 18562
rect 22818 18510 22820 18562
rect 22652 18508 22820 18510
rect 22652 18452 22708 18508
rect 22764 18498 22820 18508
rect 22988 18562 23044 20972
rect 23212 20914 23268 20926
rect 23212 20862 23214 20914
rect 23266 20862 23268 20914
rect 23100 20804 23156 20814
rect 23100 19234 23156 20748
rect 23212 20802 23268 20862
rect 23212 20750 23214 20802
rect 23266 20750 23268 20802
rect 23212 20130 23268 20750
rect 23212 20078 23214 20130
rect 23266 20078 23268 20130
rect 23212 20066 23268 20078
rect 23100 19182 23102 19234
rect 23154 19182 23156 19234
rect 23100 19170 23156 19182
rect 23324 18674 23380 21980
rect 23548 21586 23604 21598
rect 23548 21534 23550 21586
rect 23602 21534 23604 21586
rect 23548 19348 23604 21534
rect 23772 20132 23828 22428
rect 24556 22370 24612 22428
rect 24556 22318 24558 22370
rect 24610 22318 24612 22370
rect 24556 22306 24612 22318
rect 24780 22372 24836 22382
rect 24780 22278 24836 22316
rect 25004 22370 25060 22382
rect 25004 22318 25006 22370
rect 25058 22318 25060 22370
rect 24108 22260 24164 22270
rect 23884 22148 23940 22158
rect 23884 22054 23940 22092
rect 24108 21586 24164 22204
rect 25004 22260 25060 22318
rect 26124 22372 26180 22382
rect 26124 22278 26180 22316
rect 25004 22194 25060 22204
rect 26012 22258 26068 22270
rect 26012 22206 26014 22258
rect 26066 22206 26068 22258
rect 24220 21812 24276 21822
rect 24220 21698 24276 21756
rect 24220 21646 24222 21698
rect 24274 21646 24276 21698
rect 24220 21634 24276 21646
rect 26012 21700 26068 22206
rect 26236 22258 26292 23212
rect 26236 22206 26238 22258
rect 26290 22206 26292 22258
rect 26236 22194 26292 22206
rect 26012 21634 26068 21644
rect 26348 21924 26404 23436
rect 28140 23268 28196 23278
rect 27132 23044 27188 23054
rect 27132 22482 27188 22988
rect 28140 23042 28196 23212
rect 28140 22990 28142 23042
rect 28194 22990 28196 23042
rect 28140 22978 28196 22990
rect 28364 23156 28420 23662
rect 37660 23492 37716 23886
rect 40012 23604 40068 23998
rect 40012 23538 40068 23548
rect 37660 23426 37716 23436
rect 28476 23156 28532 23166
rect 28364 23154 28532 23156
rect 28364 23102 28478 23154
rect 28530 23102 28532 23154
rect 28364 23100 28532 23102
rect 27132 22430 27134 22482
rect 27186 22430 27188 22482
rect 27132 22418 27188 22430
rect 27356 22372 27412 22382
rect 27356 22278 27412 22316
rect 27692 22370 27748 22382
rect 27692 22318 27694 22370
rect 27746 22318 27748 22370
rect 27244 22258 27300 22270
rect 27244 22206 27246 22258
rect 27298 22206 27300 22258
rect 27020 22146 27076 22158
rect 27020 22094 27022 22146
rect 27074 22094 27076 22146
rect 27020 22036 27076 22094
rect 27244 22148 27300 22206
rect 27692 22148 27748 22318
rect 27244 22092 27636 22148
rect 27076 21980 27524 22036
rect 27020 21970 27076 21980
rect 24108 21534 24110 21586
rect 24162 21534 24164 21586
rect 24108 21522 24164 21534
rect 24668 21586 24724 21598
rect 24668 21534 24670 21586
rect 24722 21534 24724 21586
rect 23772 20066 23828 20076
rect 24444 21474 24500 21486
rect 24444 21422 24446 21474
rect 24498 21422 24500 21474
rect 24444 19348 24500 21422
rect 24668 19908 24724 21534
rect 26348 20916 26404 21868
rect 27132 21868 27412 21924
rect 27020 21700 27076 21710
rect 27020 21606 27076 21644
rect 26348 20914 26852 20916
rect 26348 20862 26350 20914
rect 26402 20862 26852 20914
rect 26348 20860 26852 20862
rect 26348 20850 26404 20860
rect 26796 20188 26852 20860
rect 25676 20132 25732 20142
rect 25676 20038 25732 20076
rect 26684 20132 26740 20142
rect 26796 20132 26964 20188
rect 24668 19842 24724 19852
rect 25228 20018 25284 20030
rect 25228 19966 25230 20018
rect 25282 19966 25284 20018
rect 24556 19348 24612 19358
rect 24444 19346 24612 19348
rect 24444 19294 24558 19346
rect 24610 19294 24612 19346
rect 24444 19292 24612 19294
rect 23548 19282 23604 19292
rect 24556 19282 24612 19292
rect 23884 19234 23940 19246
rect 23884 19182 23886 19234
rect 23938 19182 23940 19234
rect 23324 18622 23326 18674
rect 23378 18622 23380 18674
rect 23324 18610 23380 18622
rect 23436 19012 23492 19022
rect 23436 18676 23492 18956
rect 23884 18900 23940 19182
rect 23884 18834 23940 18844
rect 24556 19124 24612 19134
rect 23436 18620 23604 18676
rect 22988 18510 22990 18562
rect 23042 18510 23044 18562
rect 22988 18498 23044 18510
rect 23436 18452 23492 18462
rect 22540 17668 22596 17678
rect 22428 17666 22596 17668
rect 22428 17614 22542 17666
rect 22594 17614 22596 17666
rect 22428 17612 22596 17614
rect 22540 17602 22596 17612
rect 22652 17554 22708 18396
rect 22652 17502 22654 17554
rect 22706 17502 22708 17554
rect 22652 17490 22708 17502
rect 23324 18450 23492 18452
rect 23324 18398 23438 18450
rect 23490 18398 23492 18450
rect 23324 18396 23492 18398
rect 22876 17444 22932 17454
rect 23100 17444 23156 17454
rect 22876 17442 23156 17444
rect 22876 17390 22878 17442
rect 22930 17390 23102 17442
rect 23154 17390 23156 17442
rect 22876 17388 23156 17390
rect 22876 17108 22932 17388
rect 23100 17378 23156 17388
rect 22876 17042 22932 17052
rect 22092 16594 22148 16604
rect 23324 16884 23380 18396
rect 23436 18386 23492 18396
rect 23548 17556 23604 18620
rect 23548 17490 23604 17500
rect 24108 18452 24164 18462
rect 24108 17668 24164 18396
rect 24556 18340 24612 19068
rect 25228 18676 25284 19966
rect 25452 20018 25508 20030
rect 25452 19966 25454 20018
rect 25506 19966 25508 20018
rect 25340 19908 25396 19918
rect 25340 19814 25396 19852
rect 24444 17780 24500 17790
rect 24108 17554 24164 17612
rect 24108 17502 24110 17554
rect 24162 17502 24164 17554
rect 24108 17490 24164 17502
rect 24220 17724 24444 17780
rect 23436 17444 23492 17454
rect 23436 17350 23492 17388
rect 24108 16996 24164 17006
rect 24108 16902 24164 16940
rect 22988 15876 23044 15886
rect 22988 15540 23044 15820
rect 22988 15446 23044 15484
rect 22652 15426 22708 15438
rect 22652 15374 22654 15426
rect 22706 15374 22708 15426
rect 22652 15316 22708 15374
rect 23324 15428 23380 16828
rect 23436 15428 23492 15438
rect 23324 15426 23492 15428
rect 23324 15374 23438 15426
rect 23490 15374 23492 15426
rect 23324 15372 23492 15374
rect 23436 15362 23492 15372
rect 22708 15260 22932 15316
rect 22652 15250 22708 15260
rect 21644 15036 21924 15092
rect 22540 15204 22596 15214
rect 21644 14754 21700 15036
rect 21644 14702 21646 14754
rect 21698 14702 21700 14754
rect 21308 14644 21364 14654
rect 20636 14478 20638 14530
rect 20690 14478 20692 14530
rect 20636 14466 20692 14478
rect 21196 14642 21364 14644
rect 21196 14590 21310 14642
rect 21362 14590 21364 14642
rect 21196 14588 21364 14590
rect 21196 14532 21252 14588
rect 21308 14578 21364 14588
rect 21196 14466 21252 14476
rect 21644 14420 21700 14702
rect 21644 14354 21700 14364
rect 20412 14308 20468 14318
rect 20188 14306 20468 14308
rect 20188 14254 20414 14306
rect 20466 14254 20468 14306
rect 20188 14252 20468 14254
rect 20412 14242 20468 14252
rect 20524 14306 20580 14318
rect 20524 14254 20526 14306
rect 20578 14254 20580 14306
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 20524 13860 20580 14254
rect 20524 13794 20580 13804
rect 21420 14306 21476 14318
rect 21420 14254 21422 14306
rect 21474 14254 21476 14306
rect 21420 13634 21476 14254
rect 22540 13858 22596 15148
rect 22876 14530 22932 15260
rect 23660 15314 23716 15326
rect 23660 15262 23662 15314
rect 23714 15262 23716 15314
rect 23660 15148 23716 15262
rect 24108 15316 24164 15326
rect 24220 15316 24276 17724
rect 24444 17686 24500 17724
rect 24556 17666 24612 18284
rect 24556 17614 24558 17666
rect 24610 17614 24612 17666
rect 24332 17556 24388 17566
rect 24332 17462 24388 17500
rect 24556 16996 24612 17614
rect 24556 16930 24612 16940
rect 25116 18620 25284 18676
rect 24332 16884 24388 16894
rect 24332 16790 24388 16828
rect 24780 16884 24836 16894
rect 25116 16884 25172 18620
rect 25228 18452 25284 18462
rect 25228 18358 25284 18396
rect 24780 16882 24948 16884
rect 24780 16830 24782 16882
rect 24834 16830 24948 16882
rect 24780 16828 24948 16830
rect 24780 16818 24836 16828
rect 24108 15314 24276 15316
rect 24108 15262 24110 15314
rect 24162 15262 24276 15314
rect 24108 15260 24276 15262
rect 24556 16770 24612 16782
rect 24556 16718 24558 16770
rect 24610 16718 24612 16770
rect 24108 15250 24164 15260
rect 23548 15092 23716 15148
rect 23884 15204 23940 15242
rect 24556 15148 24612 16718
rect 24892 16098 24948 16828
rect 25116 16818 25172 16828
rect 25228 17892 25284 17902
rect 25228 17332 25284 17836
rect 24892 16046 24894 16098
rect 24946 16046 24948 16098
rect 24892 16034 24948 16046
rect 25228 16098 25284 17276
rect 25228 16046 25230 16098
rect 25282 16046 25284 16098
rect 25228 16034 25284 16046
rect 25116 15876 25172 15886
rect 25116 15782 25172 15820
rect 25452 15540 25508 19966
rect 26684 19346 26740 20076
rect 26684 19294 26686 19346
rect 26738 19294 26740 19346
rect 26684 19282 26740 19294
rect 26908 20018 26964 20132
rect 26908 19966 26910 20018
rect 26962 19966 26964 20018
rect 25900 19236 25956 19246
rect 25900 18674 25956 19180
rect 25900 18622 25902 18674
rect 25954 18622 25956 18674
rect 25900 18610 25956 18622
rect 26796 19124 26852 19134
rect 25788 18562 25844 18574
rect 25788 18510 25790 18562
rect 25842 18510 25844 18562
rect 25564 18450 25620 18462
rect 25564 18398 25566 18450
rect 25618 18398 25620 18450
rect 25564 18340 25620 18398
rect 25788 18452 25844 18510
rect 25788 18340 25844 18396
rect 25564 18274 25620 18284
rect 25676 18284 25844 18340
rect 26012 18450 26068 18462
rect 26012 18398 26014 18450
rect 26066 18398 26068 18450
rect 25564 17780 25620 17790
rect 25564 16994 25620 17724
rect 25676 17556 25732 18284
rect 26012 18004 26068 18398
rect 26572 18452 26628 18462
rect 26572 18358 26628 18396
rect 26796 18450 26852 19068
rect 26796 18398 26798 18450
rect 26850 18398 26852 18450
rect 26796 18386 26852 18398
rect 26908 19012 26964 19966
rect 27132 19236 27188 21868
rect 27244 21698 27300 21710
rect 27244 21646 27246 21698
rect 27298 21646 27300 21698
rect 27244 19460 27300 21646
rect 27356 21698 27412 21868
rect 27356 21646 27358 21698
rect 27410 21646 27412 21698
rect 27356 21634 27412 21646
rect 27468 21698 27524 21980
rect 27468 21646 27470 21698
rect 27522 21646 27524 21698
rect 27468 21634 27524 21646
rect 27356 21474 27412 21486
rect 27356 21422 27358 21474
rect 27410 21422 27412 21474
rect 27356 20188 27412 21422
rect 27580 21140 27636 22092
rect 27692 22082 27748 22092
rect 27804 22260 27860 22270
rect 27580 21084 27748 21140
rect 27356 20132 27636 20188
rect 27580 20130 27636 20132
rect 27580 20078 27582 20130
rect 27634 20078 27636 20130
rect 27580 20066 27636 20078
rect 27244 19394 27300 19404
rect 27132 19170 27188 19180
rect 27692 19124 27748 21084
rect 27692 19058 27748 19068
rect 27132 19012 27188 19022
rect 26964 19010 27188 19012
rect 26964 18958 27134 19010
rect 27186 18958 27188 19010
rect 26964 18956 27188 18958
rect 26348 18228 26404 18238
rect 26012 17938 26068 17948
rect 26236 18226 26404 18228
rect 26236 18174 26350 18226
rect 26402 18174 26404 18226
rect 26236 18172 26404 18174
rect 26012 17780 26068 17790
rect 25676 17490 25732 17500
rect 25788 17668 25844 17678
rect 25788 17106 25844 17612
rect 26012 17666 26068 17724
rect 26012 17614 26014 17666
rect 26066 17614 26068 17666
rect 26012 17602 26068 17614
rect 25788 17054 25790 17106
rect 25842 17054 25844 17106
rect 25788 17042 25844 17054
rect 25900 17444 25956 17454
rect 25900 17108 25956 17388
rect 26124 17442 26180 17454
rect 26124 17390 26126 17442
rect 26178 17390 26180 17442
rect 26012 17108 26068 17118
rect 25900 17106 26068 17108
rect 25900 17054 26014 17106
rect 26066 17054 26068 17106
rect 25900 17052 26068 17054
rect 26012 17042 26068 17052
rect 26124 17108 26180 17390
rect 26124 17042 26180 17052
rect 26236 17220 26292 18172
rect 26348 18162 26404 18172
rect 26348 17668 26404 17678
rect 26348 17574 26404 17612
rect 25564 16942 25566 16994
rect 25618 16942 25620 16994
rect 25564 16930 25620 16942
rect 26236 16882 26292 17164
rect 26908 16884 26964 18956
rect 27132 18946 27188 18956
rect 27804 18788 27860 22204
rect 28140 22148 28196 22158
rect 28364 22148 28420 23100
rect 28476 23090 28532 23100
rect 37660 23156 37716 23166
rect 37660 23062 37716 23100
rect 29260 23044 29316 23054
rect 29260 22950 29316 22988
rect 31388 23044 31444 23054
rect 28588 22484 28644 22494
rect 28588 22390 28644 22428
rect 31388 22484 31444 22988
rect 40012 22932 40068 22942
rect 40012 22838 40068 22876
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 31388 22418 31444 22428
rect 28140 22146 28420 22148
rect 28140 22094 28142 22146
rect 28194 22094 28420 22146
rect 28140 22092 28420 22094
rect 28476 22148 28532 22158
rect 28140 21924 28196 22092
rect 28476 22054 28532 22092
rect 28140 21858 28196 21868
rect 37884 21586 37940 21598
rect 37884 21534 37886 21586
rect 37938 21534 37940 21586
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 37660 20802 37716 20814
rect 37660 20750 37662 20802
rect 37714 20750 37716 20802
rect 29708 19908 29764 19918
rect 29260 19852 29708 19908
rect 29148 19460 29204 19470
rect 29148 19366 29204 19404
rect 29260 19346 29316 19852
rect 29708 19814 29764 19852
rect 30156 19906 30212 19918
rect 30156 19854 30158 19906
rect 30210 19854 30212 19906
rect 29260 19294 29262 19346
rect 29314 19294 29316 19346
rect 29260 19282 29316 19294
rect 27020 18732 27860 18788
rect 27020 18674 27076 18732
rect 27020 18622 27022 18674
rect 27074 18622 27076 18674
rect 27020 17108 27076 18622
rect 27244 18452 27300 18462
rect 27244 18358 27300 18396
rect 29148 18452 29204 18462
rect 27132 18338 27188 18350
rect 27132 18286 27134 18338
rect 27186 18286 27188 18338
rect 27132 17556 27188 18286
rect 29148 17890 29204 18396
rect 29148 17838 29150 17890
rect 29202 17838 29204 17890
rect 29148 17826 29204 17838
rect 29260 17556 29316 17566
rect 27132 17500 27636 17556
rect 27020 17042 27076 17052
rect 27580 16994 27636 17500
rect 29260 17462 29316 17500
rect 29708 17556 29764 17566
rect 27580 16942 27582 16994
rect 27634 16942 27636 16994
rect 27580 16930 27636 16942
rect 28588 16996 28644 17006
rect 26236 16830 26238 16882
rect 26290 16830 26292 16882
rect 26236 16818 26292 16830
rect 26796 16828 26908 16884
rect 25900 16770 25956 16782
rect 25900 16718 25902 16770
rect 25954 16718 25956 16770
rect 25900 16436 25956 16718
rect 25900 16380 26516 16436
rect 26460 16210 26516 16380
rect 26460 16158 26462 16210
rect 26514 16158 26516 16210
rect 26460 16146 26516 16158
rect 25452 15474 25508 15484
rect 25788 16098 25844 16110
rect 25788 16046 25790 16098
rect 25842 16046 25844 16098
rect 23884 15138 23940 15148
rect 24220 15092 24612 15148
rect 22876 14478 22878 14530
rect 22930 14478 22932 14530
rect 22876 14466 22932 14478
rect 23212 15036 23604 15092
rect 23212 14530 23268 15036
rect 24220 14642 24276 15092
rect 24220 14590 24222 14642
rect 24274 14590 24276 14642
rect 24220 14578 24276 14590
rect 23212 14478 23214 14530
rect 23266 14478 23268 14530
rect 23212 14466 23268 14478
rect 23436 14530 23492 14542
rect 23436 14478 23438 14530
rect 23490 14478 23492 14530
rect 22540 13806 22542 13858
rect 22594 13806 22596 13858
rect 22540 13794 22596 13806
rect 22988 14306 23044 14318
rect 22988 14254 22990 14306
rect 23042 14254 23044 14306
rect 21868 13748 21924 13758
rect 21868 13654 21924 13692
rect 21420 13582 21422 13634
rect 21474 13582 21476 13634
rect 21084 13524 21140 13534
rect 18620 13010 18676 13020
rect 19516 13010 19572 13020
rect 20748 13076 20804 13086
rect 17948 12910 17950 12962
rect 18002 12910 18004 12962
rect 17948 12898 18004 12910
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 20748 8428 20804 13020
rect 21084 12402 21140 13468
rect 21084 12350 21086 12402
rect 21138 12350 21140 12402
rect 21084 12338 21140 12350
rect 20748 8372 21140 8428
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 21084 4338 21140 8372
rect 21084 4286 21086 4338
rect 21138 4286 21140 4338
rect 21084 4274 21140 4286
rect 20860 4116 20916 4126
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 16156 3332 16212 3342
rect 16156 800 16212 3276
rect 16940 3332 16996 3342
rect 16940 3238 16996 3276
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 20860 800 20916 4060
rect 21420 3554 21476 13582
rect 22988 13636 23044 14254
rect 23436 13748 23492 14478
rect 23436 13682 23492 13692
rect 25340 13748 25396 13758
rect 25340 13654 25396 13692
rect 25788 13748 25844 16046
rect 25788 13682 25844 13692
rect 26348 15876 26404 15886
rect 26348 14642 26404 15820
rect 26348 14590 26350 14642
rect 26402 14590 26404 14642
rect 22988 13570 23044 13580
rect 24668 13636 24724 13646
rect 21644 13524 21700 13534
rect 21644 13074 21700 13468
rect 21644 13022 21646 13074
rect 21698 13022 21700 13074
rect 21644 13010 21700 13022
rect 24668 8428 24724 13580
rect 26348 8428 26404 14590
rect 26796 14306 26852 16828
rect 26908 16790 26964 16828
rect 28588 16210 28644 16940
rect 28588 16158 28590 16210
rect 28642 16158 28644 16210
rect 28588 16146 28644 16158
rect 29260 16884 29316 16894
rect 29260 16210 29316 16828
rect 29708 16770 29764 17500
rect 30156 16884 30212 19854
rect 37660 19908 37716 20750
rect 37884 20132 37940 21534
rect 39900 21474 39956 21486
rect 39900 21422 39902 21474
rect 39954 21422 39956 21474
rect 39900 20916 39956 21422
rect 39900 20850 39956 20860
rect 40012 20914 40068 20926
rect 40012 20862 40014 20914
rect 40066 20862 40068 20914
rect 40012 20244 40068 20862
rect 40012 20178 40068 20188
rect 37884 20066 37940 20076
rect 37660 19842 37716 19852
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 37660 18450 37716 18462
rect 37660 18398 37662 18450
rect 37714 18398 37716 18450
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 37660 17556 37716 18398
rect 40012 18228 40068 18238
rect 40012 18134 40068 18172
rect 37660 17490 37716 17500
rect 30156 16790 30212 16828
rect 37660 16884 37716 16894
rect 37660 16790 37716 16828
rect 29708 16718 29710 16770
rect 29762 16718 29764 16770
rect 29708 16706 29764 16718
rect 40012 16658 40068 16670
rect 40012 16606 40014 16658
rect 40066 16606 40068 16658
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 29260 16158 29262 16210
rect 29314 16158 29316 16210
rect 29260 16146 29316 16158
rect 40012 16212 40068 16606
rect 40012 16146 40068 16156
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 26796 14254 26798 14306
rect 26850 14254 26852 14306
rect 26796 13748 26852 14254
rect 26796 13682 26852 13692
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 24556 8372 24724 8428
rect 25788 8372 26404 8428
rect 22092 4116 22148 4126
rect 22092 4022 22148 4060
rect 21420 3502 21422 3554
rect 21474 3502 21476 3554
rect 21420 3490 21476 3502
rect 21532 3668 21588 3678
rect 21532 800 21588 3612
rect 22428 3668 22484 3678
rect 22428 3574 22484 3612
rect 24220 3668 24276 3678
rect 24220 800 24276 3612
rect 24556 3554 24612 8372
rect 25788 4338 25844 8372
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 25788 4286 25790 4338
rect 25842 4286 25844 4338
rect 25788 4274 25844 4286
rect 26796 4114 26852 4126
rect 26796 4062 26798 4114
rect 26850 4062 26852 4114
rect 25564 3668 25620 3678
rect 25564 3574 25620 3612
rect 24556 3502 24558 3554
rect 24610 3502 24612 3554
rect 24556 3490 24612 3502
rect 25564 3444 25620 3454
rect 25564 800 25620 3388
rect 26796 3444 26852 4062
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 26796 3378 26852 3388
rect 16128 0 16240 800
rect 20832 0 20944 800
rect 21504 0 21616 800
rect 24192 0 24304 800
rect 25536 0 25648 800
<< via2 >>
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 19516 38556 19572 38612
rect 20748 38556 20804 38612
rect 17500 36652 17556 36708
rect 18732 36706 18788 36708
rect 18732 36654 18734 36706
rect 18734 36654 18786 36706
rect 18786 36654 18788 36706
rect 18732 36652 18788 36654
rect 1708 36370 1764 36372
rect 1708 36318 1710 36370
rect 1710 36318 1762 36370
rect 1762 36318 1764 36370
rect 1708 36316 1764 36318
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 16828 28812 16884 28868
rect 4172 27580 4228 27636
rect 1932 27186 1988 27188
rect 1932 27134 1934 27186
rect 1934 27134 1986 27186
rect 1986 27134 1988 27186
rect 1932 27132 1988 27134
rect 1932 24892 1988 24948
rect 1932 24498 1988 24500
rect 1932 24446 1934 24498
rect 1934 24446 1986 24498
rect 1986 24446 1988 24498
rect 1932 24444 1988 24446
rect 1932 23548 1988 23604
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 15036 27692 15092 27748
rect 15596 27746 15652 27748
rect 15596 27694 15598 27746
rect 15598 27694 15650 27746
rect 15650 27694 15652 27746
rect 15596 27692 15652 27694
rect 16492 27692 16548 27748
rect 12124 27132 12180 27188
rect 14476 27132 14532 27188
rect 4284 27074 4340 27076
rect 4284 27022 4286 27074
rect 4286 27022 4338 27074
rect 4338 27022 4340 27074
rect 4284 27020 4340 27022
rect 14140 27020 14196 27076
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 4284 25506 4340 25508
rect 4284 25454 4286 25506
rect 4286 25454 4338 25506
rect 4338 25454 4340 25506
rect 4284 25452 4340 25454
rect 10556 25452 10612 25508
rect 4284 24722 4340 24724
rect 4284 24670 4286 24722
rect 4286 24670 4338 24722
rect 4338 24670 4340 24722
rect 4284 24668 4340 24670
rect 9996 24668 10052 24724
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 13580 25452 13636 25508
rect 9996 24050 10052 24052
rect 9996 23998 9998 24050
rect 9998 23998 10050 24050
rect 10050 23998 10052 24050
rect 9996 23996 10052 23998
rect 4284 23938 4340 23940
rect 4284 23886 4286 23938
rect 4286 23886 4338 23938
rect 4338 23886 4340 23938
rect 4284 23884 4340 23886
rect 13692 25394 13748 25396
rect 13692 25342 13694 25394
rect 13694 25342 13746 25394
rect 13746 25342 13748 25394
rect 13692 25340 13748 25342
rect 12796 24332 12852 24388
rect 13468 24892 13524 24948
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 14700 26178 14756 26180
rect 14700 26126 14702 26178
rect 14702 26126 14754 26178
rect 14754 26126 14756 26178
rect 14700 26124 14756 26126
rect 15708 26124 15764 26180
rect 16492 26124 16548 26180
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 22876 38220 22932 38276
rect 17724 28812 17780 28868
rect 15820 25506 15876 25508
rect 15820 25454 15822 25506
rect 15822 25454 15874 25506
rect 15874 25454 15876 25506
rect 15820 25452 15876 25454
rect 14588 25394 14644 25396
rect 14588 25342 14590 25394
rect 14590 25342 14642 25394
rect 14642 25342 14644 25394
rect 14588 25340 14644 25342
rect 16156 25394 16212 25396
rect 16156 25342 16158 25394
rect 16158 25342 16210 25394
rect 16210 25342 16212 25394
rect 16156 25340 16212 25342
rect 16940 25452 16996 25508
rect 16828 25340 16884 25396
rect 16492 25282 16548 25284
rect 16492 25230 16494 25282
rect 16494 25230 16546 25282
rect 16546 25230 16548 25282
rect 16492 25228 16548 25230
rect 13916 24946 13972 24948
rect 13916 24894 13918 24946
rect 13918 24894 13970 24946
rect 13970 24894 13972 24946
rect 13916 24892 13972 24894
rect 17052 25116 17108 25172
rect 13580 24220 13636 24276
rect 13692 23996 13748 24052
rect 13916 23884 13972 23940
rect 13244 23042 13300 23044
rect 13244 22990 13246 23042
rect 13246 22990 13298 23042
rect 13298 22990 13300 23042
rect 13244 22988 13300 22990
rect 13916 23212 13972 23268
rect 15932 23324 15988 23380
rect 15372 23100 15428 23156
rect 14028 22876 14084 22932
rect 15260 22988 15316 23044
rect 12796 22540 12852 22596
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 11676 20524 11732 20580
rect 4172 19964 4228 20020
rect 10108 20076 10164 20132
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 11004 20076 11060 20132
rect 14252 20076 14308 20132
rect 13804 19906 13860 19908
rect 13804 19854 13806 19906
rect 13806 19854 13858 19906
rect 13858 19854 13860 19906
rect 13804 19852 13860 19854
rect 12908 19346 12964 19348
rect 12908 19294 12910 19346
rect 12910 19294 12962 19346
rect 12962 19294 12964 19346
rect 12908 19292 12964 19294
rect 10780 19122 10836 19124
rect 10780 19070 10782 19122
rect 10782 19070 10834 19122
rect 10834 19070 10836 19122
rect 10780 19068 10836 19070
rect 13468 19122 13524 19124
rect 13468 19070 13470 19122
rect 13470 19070 13522 19122
rect 13522 19070 13524 19122
rect 13468 19068 13524 19070
rect 14812 20802 14868 20804
rect 14812 20750 14814 20802
rect 14814 20750 14866 20802
rect 14866 20750 14868 20802
rect 14812 20748 14868 20750
rect 14364 19292 14420 19348
rect 14812 19852 14868 19908
rect 14812 19234 14868 19236
rect 14812 19182 14814 19234
rect 14814 19182 14866 19234
rect 14866 19182 14868 19234
rect 14812 19180 14868 19182
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 4284 16882 4340 16884
rect 4284 16830 4286 16882
rect 4286 16830 4338 16882
rect 4338 16830 4340 16882
rect 4284 16828 4340 16830
rect 12236 16828 12292 16884
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 1932 16156 1988 16212
rect 12908 16882 12964 16884
rect 12908 16830 12910 16882
rect 12910 16830 12962 16882
rect 12962 16830 12964 16882
rect 12908 16828 12964 16830
rect 13692 16940 13748 16996
rect 17164 23884 17220 23940
rect 18172 27746 18228 27748
rect 18172 27694 18174 27746
rect 18174 27694 18226 27746
rect 18226 27694 18228 27746
rect 18172 27692 18228 27694
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 25564 38274 25620 38276
rect 25564 38222 25566 38274
rect 25566 38222 25618 38274
rect 25618 38222 25620 38274
rect 25564 38220 25620 38222
rect 23548 36652 23604 36708
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 19516 28530 19572 28532
rect 19516 28478 19518 28530
rect 19518 28478 19570 28530
rect 19570 28478 19572 28530
rect 19516 28476 19572 28478
rect 19516 27692 19572 27748
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 17500 26178 17556 26180
rect 17500 26126 17502 26178
rect 17502 26126 17554 26178
rect 17554 26126 17556 26178
rect 17500 26124 17556 26126
rect 19516 26178 19572 26180
rect 19516 26126 19518 26178
rect 19518 26126 19570 26178
rect 19570 26126 19572 26178
rect 19516 26124 19572 26126
rect 18620 25394 18676 25396
rect 18620 25342 18622 25394
rect 18622 25342 18674 25394
rect 18674 25342 18676 25394
rect 18620 25340 18676 25342
rect 17612 25116 17668 25172
rect 17836 25228 17892 25284
rect 18284 25282 18340 25284
rect 18284 25230 18286 25282
rect 18286 25230 18338 25282
rect 18338 25230 18340 25282
rect 18284 25228 18340 25230
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 20300 28476 20356 28532
rect 20524 26124 20580 26180
rect 20748 26796 20804 26852
rect 20188 25564 20244 25620
rect 20188 25228 20244 25284
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 17500 23548 17556 23604
rect 17724 23772 17780 23828
rect 16828 22988 16884 23044
rect 16380 22092 16436 22148
rect 17388 23266 17444 23268
rect 17388 23214 17390 23266
rect 17390 23214 17442 23266
rect 17442 23214 17444 23266
rect 17388 23212 17444 23214
rect 17724 23378 17780 23380
rect 17724 23326 17726 23378
rect 17726 23326 17778 23378
rect 17778 23326 17780 23378
rect 17724 23324 17780 23326
rect 18284 24780 18340 24836
rect 18172 23826 18228 23828
rect 18172 23774 18174 23826
rect 18174 23774 18226 23826
rect 18226 23774 18228 23826
rect 18172 23772 18228 23774
rect 18508 23938 18564 23940
rect 18508 23886 18510 23938
rect 18510 23886 18562 23938
rect 18562 23886 18564 23938
rect 18508 23884 18564 23886
rect 18060 23042 18116 23044
rect 18060 22990 18062 23042
rect 18062 22990 18114 23042
rect 18114 22990 18116 23042
rect 18060 22988 18116 22990
rect 17836 22930 17892 22932
rect 17836 22878 17838 22930
rect 17838 22878 17890 22930
rect 17890 22878 17892 22930
rect 17836 22876 17892 22878
rect 17052 21644 17108 21700
rect 17276 22204 17332 22260
rect 16380 20748 16436 20804
rect 15372 20578 15428 20580
rect 15372 20526 15374 20578
rect 15374 20526 15426 20578
rect 15426 20526 15428 20578
rect 15372 20524 15428 20526
rect 15260 20076 15316 20132
rect 16604 20972 16660 21028
rect 17164 20972 17220 21028
rect 15484 19234 15540 19236
rect 15484 19182 15486 19234
rect 15486 19182 15538 19234
rect 15538 19182 15540 19234
rect 15484 19180 15540 19182
rect 16044 18956 16100 19012
rect 15036 18620 15092 18676
rect 16268 18674 16324 18676
rect 16268 18622 16270 18674
rect 16270 18622 16322 18674
rect 16322 18622 16324 18674
rect 16268 18620 16324 18622
rect 14812 17948 14868 18004
rect 17724 21698 17780 21700
rect 17724 21646 17726 21698
rect 17726 21646 17778 21698
rect 17778 21646 17780 21698
rect 17724 21644 17780 21646
rect 17388 19404 17444 19460
rect 17052 19180 17108 19236
rect 16940 18956 16996 19012
rect 16716 18620 16772 18676
rect 16268 18226 16324 18228
rect 16268 18174 16270 18226
rect 16270 18174 16322 18226
rect 16322 18174 16324 18226
rect 16268 18172 16324 18174
rect 14924 17554 14980 17556
rect 14924 17502 14926 17554
rect 14926 17502 14978 17554
rect 14978 17502 14980 17554
rect 14924 17500 14980 17502
rect 14588 16940 14644 16996
rect 14252 16828 14308 16884
rect 15708 16770 15764 16772
rect 15708 16718 15710 16770
rect 15710 16718 15762 16770
rect 15762 16718 15764 16770
rect 15708 16716 15764 16718
rect 16156 16828 16212 16884
rect 12236 16044 12292 16100
rect 15820 16098 15876 16100
rect 15820 16046 15822 16098
rect 15822 16046 15874 16098
rect 15874 16046 15876 16098
rect 15820 16044 15876 16046
rect 14476 15986 14532 15988
rect 14476 15934 14478 15986
rect 14478 15934 14530 15986
rect 14530 15934 14532 15986
rect 14476 15932 14532 15934
rect 14252 15372 14308 15428
rect 17052 18172 17108 18228
rect 16716 17554 16772 17556
rect 16716 17502 16718 17554
rect 16718 17502 16770 17554
rect 16770 17502 16772 17554
rect 16716 17500 16772 17502
rect 16940 17442 16996 17444
rect 16940 17390 16942 17442
rect 16942 17390 16994 17442
rect 16994 17390 16996 17442
rect 16940 17388 16996 17390
rect 16492 17052 16548 17108
rect 16380 16828 16436 16884
rect 16268 16604 16324 16660
rect 16604 15986 16660 15988
rect 16604 15934 16606 15986
rect 16606 15934 16658 15986
rect 16658 15934 16660 15986
rect 16604 15932 16660 15934
rect 16828 15820 16884 15876
rect 17612 20860 17668 20916
rect 18060 20860 18116 20916
rect 17836 20690 17892 20692
rect 17836 20638 17838 20690
rect 17838 20638 17890 20690
rect 17890 20638 17892 20690
rect 17836 20636 17892 20638
rect 17388 17106 17444 17108
rect 17388 17054 17390 17106
rect 17390 17054 17442 17106
rect 17442 17054 17444 17106
rect 17388 17052 17444 17054
rect 18396 23548 18452 23604
rect 18396 22258 18452 22260
rect 18396 22206 18398 22258
rect 18398 22206 18450 22258
rect 18450 22206 18452 22258
rect 18396 22204 18452 22206
rect 19964 24834 20020 24836
rect 19964 24782 19966 24834
rect 19966 24782 20018 24834
rect 20018 24782 20020 24834
rect 19964 24780 20020 24782
rect 22540 27804 22596 27860
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 26236 37884 26292 37940
rect 27468 37938 27524 37940
rect 27468 37886 27470 37938
rect 27470 37886 27522 37938
rect 27522 37886 27524 37938
rect 27468 37884 27524 37886
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 24780 36706 24836 36708
rect 24780 36654 24782 36706
rect 24782 36654 24834 36706
rect 24834 36654 24836 36706
rect 24780 36652 24836 36654
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 23772 27804 23828 27860
rect 24444 27858 24500 27860
rect 24444 27806 24446 27858
rect 24446 27806 24498 27858
rect 24498 27806 24500 27858
rect 24444 27804 24500 27806
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 20972 26348 21028 26404
rect 21420 27074 21476 27076
rect 21420 27022 21422 27074
rect 21422 27022 21474 27074
rect 21474 27022 21476 27074
rect 21420 27020 21476 27022
rect 19852 23884 19908 23940
rect 19964 23826 20020 23828
rect 19964 23774 19966 23826
rect 19966 23774 20018 23826
rect 20018 23774 20020 23826
rect 19964 23772 20020 23774
rect 19628 23548 19684 23604
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 19404 23266 19460 23268
rect 19404 23214 19406 23266
rect 19406 23214 19458 23266
rect 19458 23214 19460 23266
rect 19404 23212 19460 23214
rect 18396 21868 18452 21924
rect 18508 20748 18564 20804
rect 18508 19906 18564 19908
rect 18508 19854 18510 19906
rect 18510 19854 18562 19906
rect 18562 19854 18564 19906
rect 18508 19852 18564 19854
rect 18284 19180 18340 19236
rect 17948 19068 18004 19124
rect 17612 17612 17668 17668
rect 17724 16770 17780 16772
rect 17724 16718 17726 16770
rect 17726 16718 17778 16770
rect 17778 16718 17780 16770
rect 17724 16716 17780 16718
rect 18508 18450 18564 18452
rect 18508 18398 18510 18450
rect 18510 18398 18562 18450
rect 18562 18398 18564 18450
rect 18508 18396 18564 18398
rect 18508 17724 18564 17780
rect 18956 22876 19012 22932
rect 18844 20636 18900 20692
rect 18844 19852 18900 19908
rect 18844 17666 18900 17668
rect 18844 17614 18846 17666
rect 18846 17614 18898 17666
rect 18898 17614 18900 17666
rect 18844 17612 18900 17614
rect 18732 16940 18788 16996
rect 18172 16716 18228 16772
rect 18284 16828 18340 16884
rect 17276 15596 17332 15652
rect 17276 15148 17332 15204
rect 17500 15538 17556 15540
rect 17500 15486 17502 15538
rect 17502 15486 17554 15538
rect 17554 15486 17556 15538
rect 17500 15484 17556 15486
rect 17724 15874 17780 15876
rect 17724 15822 17726 15874
rect 17726 15822 17778 15874
rect 17778 15822 17780 15874
rect 17724 15820 17780 15822
rect 18172 15260 18228 15316
rect 20412 23660 20468 23716
rect 20188 23154 20244 23156
rect 20188 23102 20190 23154
rect 20190 23102 20242 23154
rect 20242 23102 20244 23154
rect 20188 23100 20244 23102
rect 20524 23154 20580 23156
rect 20524 23102 20526 23154
rect 20526 23102 20578 23154
rect 20578 23102 20580 23154
rect 20524 23100 20580 23102
rect 21308 23660 21364 23716
rect 21756 26962 21812 26964
rect 21756 26910 21758 26962
rect 21758 26910 21810 26962
rect 21810 26910 21812 26962
rect 21756 26908 21812 26910
rect 21532 26850 21588 26852
rect 21532 26798 21534 26850
rect 21534 26798 21586 26850
rect 21586 26798 21588 26850
rect 21532 26796 21588 26798
rect 21868 26124 21924 26180
rect 22428 26962 22484 26964
rect 22428 26910 22430 26962
rect 22430 26910 22482 26962
rect 22482 26910 22484 26962
rect 22428 26908 22484 26910
rect 22988 26348 23044 26404
rect 23548 26402 23604 26404
rect 23548 26350 23550 26402
rect 23550 26350 23602 26402
rect 23602 26350 23604 26402
rect 23548 26348 23604 26350
rect 23996 26348 24052 26404
rect 25228 26348 25284 26404
rect 22316 26178 22372 26180
rect 22316 26126 22318 26178
rect 22318 26126 22370 26178
rect 22370 26126 22372 26178
rect 22316 26124 22372 26126
rect 22428 25618 22484 25620
rect 22428 25566 22430 25618
rect 22430 25566 22482 25618
rect 22482 25566 22484 25618
rect 22428 25564 22484 25566
rect 21868 25394 21924 25396
rect 21868 25342 21870 25394
rect 21870 25342 21922 25394
rect 21922 25342 21924 25394
rect 21868 25340 21924 25342
rect 21532 25282 21588 25284
rect 21532 25230 21534 25282
rect 21534 25230 21586 25282
rect 21586 25230 21588 25282
rect 21532 25228 21588 25230
rect 21756 25282 21812 25284
rect 21756 25230 21758 25282
rect 21758 25230 21810 25282
rect 21810 25230 21812 25282
rect 21756 25228 21812 25230
rect 22316 25282 22372 25284
rect 22316 25230 22318 25282
rect 22318 25230 22370 25282
rect 22370 25230 22372 25282
rect 22316 25228 22372 25230
rect 24108 24834 24164 24836
rect 24108 24782 24110 24834
rect 24110 24782 24162 24834
rect 24162 24782 24164 24834
rect 24108 24780 24164 24782
rect 21644 23378 21700 23380
rect 21644 23326 21646 23378
rect 21646 23326 21698 23378
rect 21698 23326 21700 23378
rect 21644 23324 21700 23326
rect 20412 22988 20468 23044
rect 19852 22092 19908 22148
rect 19180 21868 19236 21924
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 19852 20860 19908 20916
rect 19068 20018 19124 20020
rect 19068 19966 19070 20018
rect 19070 19966 19122 20018
rect 19122 19966 19124 20018
rect 19068 19964 19124 19966
rect 19292 18956 19348 19012
rect 19628 20748 19684 20804
rect 19516 20018 19572 20020
rect 19516 19966 19518 20018
rect 19518 19966 19570 20018
rect 19570 19966 19572 20018
rect 19516 19964 19572 19966
rect 19404 18396 19460 18452
rect 20300 20748 20356 20804
rect 20412 20636 20468 20692
rect 20524 22092 20580 22148
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 20188 19964 20244 20020
rect 19852 19346 19908 19348
rect 19852 19294 19854 19346
rect 19854 19294 19906 19346
rect 19906 19294 19908 19346
rect 19852 19292 19908 19294
rect 20188 19292 20244 19348
rect 20076 19068 20132 19124
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 19516 17612 19572 17668
rect 19852 17724 19908 17780
rect 20748 21756 20804 21812
rect 21196 23100 21252 23156
rect 22316 23324 22372 23380
rect 21420 22540 21476 22596
rect 21756 23154 21812 23156
rect 21756 23102 21758 23154
rect 21758 23102 21810 23154
rect 21810 23102 21812 23154
rect 21756 23100 21812 23102
rect 21308 21756 21364 21812
rect 21196 19458 21252 19460
rect 21196 19406 21198 19458
rect 21198 19406 21250 19458
rect 21250 19406 21252 19458
rect 21196 19404 21252 19406
rect 21308 19292 21364 19348
rect 20524 18732 20580 18788
rect 20412 17836 20468 17892
rect 20300 17612 20356 17668
rect 18956 15148 19012 15204
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 15484 14924 15540 14980
rect 19516 17442 19572 17444
rect 19516 17390 19518 17442
rect 19518 17390 19570 17442
rect 19570 17390 19572 17442
rect 19516 17388 19572 17390
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 20300 16658 20356 16660
rect 20300 16606 20302 16658
rect 20302 16606 20354 16658
rect 20354 16606 20356 16658
rect 20300 16604 20356 16606
rect 20524 17724 20580 17780
rect 20524 16940 20580 16996
rect 19852 16044 19908 16100
rect 20300 16044 20356 16100
rect 20076 15874 20132 15876
rect 20076 15822 20078 15874
rect 20078 15822 20130 15874
rect 20130 15822 20132 15874
rect 20076 15820 20132 15822
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 19068 14812 19124 14868
rect 19516 15314 19572 15316
rect 19516 15262 19518 15314
rect 19518 15262 19570 15314
rect 19570 15262 19572 15314
rect 19516 15260 19572 15262
rect 19852 15202 19908 15204
rect 19852 15150 19854 15202
rect 19854 15150 19906 15202
rect 19906 15150 19908 15202
rect 19852 15148 19908 15150
rect 20188 15036 20244 15092
rect 15596 14252 15652 14308
rect 18060 14306 18116 14308
rect 18060 14254 18062 14306
rect 18062 14254 18114 14306
rect 18114 14254 18116 14306
rect 18060 14252 18116 14254
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 18620 13468 18676 13524
rect 19292 14418 19348 14420
rect 19292 14366 19294 14418
rect 19294 14366 19346 14418
rect 19346 14366 19348 14418
rect 19292 14364 19348 14366
rect 19292 13858 19348 13860
rect 19292 13806 19294 13858
rect 19294 13806 19346 13858
rect 19346 13806 19348 13858
rect 19292 13804 19348 13806
rect 20300 14530 20356 14532
rect 20300 14478 20302 14530
rect 20302 14478 20354 14530
rect 20354 14478 20356 14530
rect 20300 14476 20356 14478
rect 21756 22204 21812 22260
rect 21532 20636 21588 20692
rect 22092 22092 22148 22148
rect 23996 23772 24052 23828
rect 22540 22988 22596 23044
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 25676 24780 25732 24836
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 40012 24220 40068 24276
rect 37660 24108 37716 24164
rect 25676 24050 25732 24052
rect 25676 23998 25678 24050
rect 25678 23998 25730 24050
rect 25730 23998 25732 24050
rect 25676 23996 25732 23998
rect 25228 23436 25284 23492
rect 26124 23436 26180 23492
rect 26236 23212 26292 23268
rect 25116 22988 25172 23044
rect 26012 23042 26068 23044
rect 26012 22990 26014 23042
rect 26014 22990 26066 23042
rect 26066 22990 26068 23042
rect 26012 22988 26068 22990
rect 22540 22092 22596 22148
rect 22204 20748 22260 20804
rect 21532 19122 21588 19124
rect 21532 19070 21534 19122
rect 21534 19070 21586 19122
rect 21586 19070 21588 19122
rect 21532 19068 21588 19070
rect 21644 20076 21700 20132
rect 21308 17948 21364 18004
rect 21756 18732 21812 18788
rect 21868 19964 21924 20020
rect 21868 17890 21924 17892
rect 21868 17838 21870 17890
rect 21870 17838 21922 17890
rect 21922 17838 21924 17890
rect 21868 17836 21924 17838
rect 22764 19292 22820 19348
rect 23100 22146 23156 22148
rect 23100 22094 23102 22146
rect 23102 22094 23154 22146
rect 23154 22094 23156 22146
rect 23100 22092 23156 22094
rect 22988 21810 23044 21812
rect 22988 21758 22990 21810
rect 22990 21758 23042 21810
rect 23042 21758 23044 21810
rect 22988 21756 23044 21758
rect 23212 21756 23268 21812
rect 23660 22146 23716 22148
rect 23660 22094 23662 22146
rect 23662 22094 23714 22146
rect 23714 22094 23716 22146
rect 23660 22092 23716 22094
rect 23324 21980 23380 22036
rect 23100 21698 23156 21700
rect 23100 21646 23102 21698
rect 23102 21646 23154 21698
rect 23154 21646 23156 21698
rect 23100 21644 23156 21646
rect 22876 18956 22932 19012
rect 22988 20972 23044 21028
rect 22428 17724 22484 17780
rect 21532 17666 21588 17668
rect 21532 17614 21534 17666
rect 21534 17614 21586 17666
rect 21586 17614 21588 17666
rect 21532 17612 21588 17614
rect 21532 17164 21588 17220
rect 21644 17106 21700 17108
rect 21644 17054 21646 17106
rect 21646 17054 21698 17106
rect 21698 17054 21700 17106
rect 21644 17052 21700 17054
rect 21868 16828 21924 16884
rect 21644 16658 21700 16660
rect 21644 16606 21646 16658
rect 21646 16606 21698 16658
rect 21698 16606 21700 16658
rect 21644 16604 21700 16606
rect 23100 20748 23156 20804
rect 24780 22370 24836 22372
rect 24780 22318 24782 22370
rect 24782 22318 24834 22370
rect 24834 22318 24836 22370
rect 24780 22316 24836 22318
rect 24108 22204 24164 22260
rect 23884 22146 23940 22148
rect 23884 22094 23886 22146
rect 23886 22094 23938 22146
rect 23938 22094 23940 22146
rect 23884 22092 23940 22094
rect 26124 22370 26180 22372
rect 26124 22318 26126 22370
rect 26126 22318 26178 22370
rect 26178 22318 26180 22370
rect 26124 22316 26180 22318
rect 25004 22204 25060 22260
rect 24220 21756 24276 21812
rect 26012 21644 26068 21700
rect 28140 23212 28196 23268
rect 27132 22988 27188 23044
rect 40012 23548 40068 23604
rect 37660 23436 37716 23492
rect 27356 22370 27412 22372
rect 27356 22318 27358 22370
rect 27358 22318 27410 22370
rect 27410 22318 27412 22370
rect 27356 22316 27412 22318
rect 27020 21980 27076 22036
rect 26348 21868 26404 21924
rect 23772 20076 23828 20132
rect 23548 19292 23604 19348
rect 27020 21698 27076 21700
rect 27020 21646 27022 21698
rect 27022 21646 27074 21698
rect 27074 21646 27076 21698
rect 27020 21644 27076 21646
rect 25676 20130 25732 20132
rect 25676 20078 25678 20130
rect 25678 20078 25730 20130
rect 25730 20078 25732 20130
rect 25676 20076 25732 20078
rect 26684 20076 26740 20132
rect 24668 19852 24724 19908
rect 23436 19010 23492 19012
rect 23436 18958 23438 19010
rect 23438 18958 23490 19010
rect 23490 18958 23492 19010
rect 23436 18956 23492 18958
rect 23884 18844 23940 18900
rect 24556 19068 24612 19124
rect 22652 18396 22708 18452
rect 22876 17052 22932 17108
rect 22092 16604 22148 16660
rect 23548 17500 23604 17556
rect 24108 18396 24164 18452
rect 25340 19906 25396 19908
rect 25340 19854 25342 19906
rect 25342 19854 25394 19906
rect 25394 19854 25396 19906
rect 25340 19852 25396 19854
rect 24556 18284 24612 18340
rect 24108 17612 24164 17668
rect 24444 17778 24500 17780
rect 24444 17726 24446 17778
rect 24446 17726 24498 17778
rect 24498 17726 24500 17778
rect 24444 17724 24500 17726
rect 23436 17442 23492 17444
rect 23436 17390 23438 17442
rect 23438 17390 23490 17442
rect 23490 17390 23492 17442
rect 23436 17388 23492 17390
rect 24108 16994 24164 16996
rect 24108 16942 24110 16994
rect 24110 16942 24162 16994
rect 24162 16942 24164 16994
rect 24108 16940 24164 16942
rect 23324 16828 23380 16884
rect 22988 15820 23044 15876
rect 22988 15538 23044 15540
rect 22988 15486 22990 15538
rect 22990 15486 23042 15538
rect 23042 15486 23044 15538
rect 22988 15484 23044 15486
rect 22652 15260 22708 15316
rect 22540 15148 22596 15204
rect 21196 14476 21252 14532
rect 21644 14364 21700 14420
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 20524 13804 20580 13860
rect 24332 17554 24388 17556
rect 24332 17502 24334 17554
rect 24334 17502 24386 17554
rect 24386 17502 24388 17554
rect 24332 17500 24388 17502
rect 24556 16940 24612 16996
rect 24332 16882 24388 16884
rect 24332 16830 24334 16882
rect 24334 16830 24386 16882
rect 24386 16830 24388 16882
rect 24332 16828 24388 16830
rect 25228 18450 25284 18452
rect 25228 18398 25230 18450
rect 25230 18398 25282 18450
rect 25282 18398 25284 18450
rect 25228 18396 25284 18398
rect 23884 15202 23940 15204
rect 23884 15150 23886 15202
rect 23886 15150 23938 15202
rect 23938 15150 23940 15202
rect 23884 15148 23940 15150
rect 25116 16828 25172 16884
rect 25228 17836 25284 17892
rect 25228 17276 25284 17332
rect 25116 15874 25172 15876
rect 25116 15822 25118 15874
rect 25118 15822 25170 15874
rect 25170 15822 25172 15874
rect 25116 15820 25172 15822
rect 25900 19180 25956 19236
rect 26796 19068 26852 19124
rect 25788 18396 25844 18452
rect 25564 18284 25620 18340
rect 25564 17724 25620 17780
rect 26572 18450 26628 18452
rect 26572 18398 26574 18450
rect 26574 18398 26626 18450
rect 26626 18398 26628 18450
rect 26572 18396 26628 18398
rect 27692 22092 27748 22148
rect 27804 22204 27860 22260
rect 27244 19404 27300 19460
rect 27132 19180 27188 19236
rect 27692 19068 27748 19124
rect 26908 18956 26964 19012
rect 26012 17948 26068 18004
rect 26012 17724 26068 17780
rect 25676 17500 25732 17556
rect 25788 17612 25844 17668
rect 25900 17388 25956 17444
rect 26124 17052 26180 17108
rect 26348 17666 26404 17668
rect 26348 17614 26350 17666
rect 26350 17614 26402 17666
rect 26402 17614 26404 17666
rect 26348 17612 26404 17614
rect 26236 17164 26292 17220
rect 37660 23154 37716 23156
rect 37660 23102 37662 23154
rect 37662 23102 37714 23154
rect 37714 23102 37716 23154
rect 37660 23100 37716 23102
rect 29260 23042 29316 23044
rect 29260 22990 29262 23042
rect 29262 22990 29314 23042
rect 29314 22990 29316 23042
rect 29260 22988 29316 22990
rect 31388 23042 31444 23044
rect 31388 22990 31390 23042
rect 31390 22990 31442 23042
rect 31442 22990 31444 23042
rect 31388 22988 31444 22990
rect 28588 22482 28644 22484
rect 28588 22430 28590 22482
rect 28590 22430 28642 22482
rect 28642 22430 28644 22482
rect 28588 22428 28644 22430
rect 40012 22930 40068 22932
rect 40012 22878 40014 22930
rect 40014 22878 40066 22930
rect 40066 22878 40068 22930
rect 40012 22876 40068 22878
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 31388 22428 31444 22484
rect 28476 22146 28532 22148
rect 28476 22094 28478 22146
rect 28478 22094 28530 22146
rect 28530 22094 28532 22146
rect 28476 22092 28532 22094
rect 28140 21868 28196 21924
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 29708 19906 29764 19908
rect 29708 19854 29710 19906
rect 29710 19854 29762 19906
rect 29762 19854 29764 19906
rect 29708 19852 29764 19854
rect 29148 19458 29204 19460
rect 29148 19406 29150 19458
rect 29150 19406 29202 19458
rect 29202 19406 29204 19458
rect 29148 19404 29204 19406
rect 27244 18450 27300 18452
rect 27244 18398 27246 18450
rect 27246 18398 27298 18450
rect 27298 18398 27300 18450
rect 27244 18396 27300 18398
rect 29148 18396 29204 18452
rect 27020 17052 27076 17108
rect 29260 17554 29316 17556
rect 29260 17502 29262 17554
rect 29262 17502 29314 17554
rect 29314 17502 29316 17554
rect 29260 17500 29316 17502
rect 29708 17500 29764 17556
rect 28588 16940 28644 16996
rect 26908 16882 26964 16884
rect 26908 16830 26910 16882
rect 26910 16830 26962 16882
rect 26962 16830 26964 16882
rect 26908 16828 26964 16830
rect 25452 15484 25508 15540
rect 21868 13746 21924 13748
rect 21868 13694 21870 13746
rect 21870 13694 21922 13746
rect 21922 13694 21924 13746
rect 21868 13692 21924 13694
rect 21084 13468 21140 13524
rect 19516 13020 19572 13076
rect 20748 13074 20804 13076
rect 20748 13022 20750 13074
rect 20750 13022 20802 13074
rect 20802 13022 20804 13074
rect 20748 13020 20804 13022
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 20860 4060 20916 4116
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 16156 3276 16212 3332
rect 16940 3330 16996 3332
rect 16940 3278 16942 3330
rect 16942 3278 16994 3330
rect 16994 3278 16996 3330
rect 16940 3276 16996 3278
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 23436 13692 23492 13748
rect 25340 13746 25396 13748
rect 25340 13694 25342 13746
rect 25342 13694 25394 13746
rect 25394 13694 25396 13746
rect 25340 13692 25396 13694
rect 25788 13692 25844 13748
rect 26348 15820 26404 15876
rect 22988 13580 23044 13636
rect 24668 13634 24724 13636
rect 24668 13582 24670 13634
rect 24670 13582 24722 13634
rect 24722 13582 24724 13634
rect 24668 13580 24724 13582
rect 21644 13468 21700 13524
rect 29260 16828 29316 16884
rect 39900 20860 39956 20916
rect 40012 20188 40068 20244
rect 37884 20076 37940 20132
rect 37660 19852 37716 19908
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 40012 18226 40068 18228
rect 40012 18174 40014 18226
rect 40014 18174 40066 18226
rect 40066 18174 40068 18226
rect 40012 18172 40068 18174
rect 37660 17500 37716 17556
rect 30156 16882 30212 16884
rect 30156 16830 30158 16882
rect 30158 16830 30210 16882
rect 30210 16830 30212 16882
rect 30156 16828 30212 16830
rect 37660 16882 37716 16884
rect 37660 16830 37662 16882
rect 37662 16830 37714 16882
rect 37714 16830 37716 16882
rect 37660 16828 37716 16830
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 40012 16156 40068 16212
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 26796 13692 26852 13748
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 22092 4114 22148 4116
rect 22092 4062 22094 4114
rect 22094 4062 22146 4114
rect 22146 4062 22148 4114
rect 22092 4060 22148 4062
rect 21532 3612 21588 3668
rect 22428 3666 22484 3668
rect 22428 3614 22430 3666
rect 22430 3614 22482 3666
rect 22482 3614 22484 3666
rect 22428 3612 22484 3614
rect 24220 3612 24276 3668
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 25564 3666 25620 3668
rect 25564 3614 25566 3666
rect 25566 3614 25618 3666
rect 25618 3614 25620 3666
rect 25564 3612 25620 3614
rect 25564 3388 25620 3444
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 26796 3388 26852 3444
<< metal3 >>
rect 19506 38556 19516 38612
rect 19572 38556 20748 38612
rect 20804 38556 20814 38612
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 22866 38220 22876 38276
rect 22932 38220 25564 38276
rect 25620 38220 25630 38276
rect 26226 37884 26236 37940
rect 26292 37884 27468 37940
rect 27524 37884 27534 37940
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 17490 36652 17500 36708
rect 17556 36652 18732 36708
rect 18788 36652 18798 36708
rect 23538 36652 23548 36708
rect 23604 36652 24780 36708
rect 24836 36652 24846 36708
rect 0 36372 800 36400
rect 0 36316 1708 36372
rect 1764 36316 1774 36372
rect 0 36288 800 36316
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 16818 28812 16828 28868
rect 16884 28812 17724 28868
rect 17780 28812 17790 28868
rect 19506 28476 19516 28532
rect 19572 28476 20300 28532
rect 20356 28476 20366 28532
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 22530 27804 22540 27860
rect 22596 27804 23772 27860
rect 23828 27804 24444 27860
rect 24500 27804 24510 27860
rect 15026 27692 15036 27748
rect 15092 27692 15596 27748
rect 15652 27692 16492 27748
rect 16548 27692 16558 27748
rect 18162 27692 18172 27748
rect 18228 27692 19516 27748
rect 19572 27692 19582 27748
rect 0 27636 800 27664
rect 0 27580 4172 27636
rect 4228 27580 4238 27636
rect 0 27552 800 27580
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 1922 27132 1932 27188
rect 1988 27132 1998 27188
rect 8372 27132 12124 27188
rect 12180 27132 14476 27188
rect 14532 27132 14542 27188
rect 0 26964 800 26992
rect 1932 26964 1988 27132
rect 8372 27076 8428 27132
rect 4274 27020 4284 27076
rect 4340 27020 8428 27076
rect 14130 27020 14140 27076
rect 14196 27020 21420 27076
rect 21476 27020 21486 27076
rect 0 26908 1988 26964
rect 21746 26908 21756 26964
rect 21812 26908 22428 26964
rect 22484 26908 22494 26964
rect 0 26880 800 26908
rect 20738 26796 20748 26852
rect 20804 26796 21532 26852
rect 21588 26796 21598 26852
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 20962 26348 20972 26404
rect 21028 26348 22988 26404
rect 23044 26348 23548 26404
rect 23604 26348 23996 26404
rect 24052 26348 25228 26404
rect 25284 26348 25294 26404
rect 14690 26124 14700 26180
rect 14756 26124 15708 26180
rect 15764 26124 15774 26180
rect 16482 26124 16492 26180
rect 16548 26124 17500 26180
rect 17556 26124 19516 26180
rect 19572 26124 20524 26180
rect 20580 26124 20590 26180
rect 21858 26124 21868 26180
rect 21924 26124 22316 26180
rect 22372 26124 22382 26180
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 20178 25564 20188 25620
rect 20244 25564 22428 25620
rect 22484 25564 22494 25620
rect 4274 25452 4284 25508
rect 4340 25452 10556 25508
rect 10612 25452 13580 25508
rect 13636 25452 13646 25508
rect 15810 25452 15820 25508
rect 15876 25452 16940 25508
rect 16996 25452 17006 25508
rect 13682 25340 13692 25396
rect 13748 25340 14588 25396
rect 14644 25340 16156 25396
rect 16212 25340 16828 25396
rect 16884 25340 16894 25396
rect 18610 25340 18620 25396
rect 18676 25340 21868 25396
rect 21924 25340 21934 25396
rect 16482 25228 16492 25284
rect 16548 25228 17836 25284
rect 17892 25228 18284 25284
rect 18340 25228 18350 25284
rect 20178 25228 20188 25284
rect 20244 25228 21532 25284
rect 21588 25228 21598 25284
rect 21746 25228 21756 25284
rect 21812 25228 22316 25284
rect 22372 25228 22382 25284
rect 17042 25116 17052 25172
rect 17108 25116 17612 25172
rect 17668 25116 17678 25172
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 0 24948 800 24976
rect 0 24892 1932 24948
rect 1988 24892 1998 24948
rect 13458 24892 13468 24948
rect 13524 24892 13916 24948
rect 13972 24892 13982 24948
rect 0 24864 800 24892
rect 18274 24780 18284 24836
rect 18340 24780 19964 24836
rect 20020 24780 20030 24836
rect 24098 24780 24108 24836
rect 24164 24780 25676 24836
rect 25732 24780 25742 24836
rect 4274 24668 4284 24724
rect 4340 24668 9996 24724
rect 10052 24668 10062 24724
rect 1922 24444 1932 24500
rect 1988 24444 1998 24500
rect 0 24276 800 24304
rect 1932 24276 1988 24444
rect 12786 24332 12796 24388
rect 12852 24332 13636 24388
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 13580 24276 13636 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 41200 24276 42000 24304
rect 0 24220 1988 24276
rect 13570 24220 13580 24276
rect 13636 24220 13646 24276
rect 40002 24220 40012 24276
rect 40068 24220 42000 24276
rect 0 24192 800 24220
rect 41200 24192 42000 24220
rect 31892 24108 37660 24164
rect 37716 24108 37726 24164
rect 31892 24052 31948 24108
rect 9986 23996 9996 24052
rect 10052 23996 13692 24052
rect 13748 23996 13758 24052
rect 25666 23996 25676 24052
rect 25732 23996 31948 24052
rect 4274 23884 4284 23940
rect 4340 23884 13916 23940
rect 13972 23884 13982 23940
rect 17154 23884 17164 23940
rect 17220 23884 18508 23940
rect 18564 23884 19852 23940
rect 19908 23884 19918 23940
rect 17714 23772 17724 23828
rect 17780 23772 18172 23828
rect 18228 23772 19964 23828
rect 20020 23772 23996 23828
rect 24052 23772 24062 23828
rect 20402 23660 20412 23716
rect 20468 23660 21308 23716
rect 21364 23660 21374 23716
rect 0 23604 800 23632
rect 41200 23604 42000 23632
rect 0 23548 1932 23604
rect 1988 23548 1998 23604
rect 17490 23548 17500 23604
rect 17556 23548 18396 23604
rect 18452 23548 19628 23604
rect 19684 23548 19694 23604
rect 40002 23548 40012 23604
rect 40068 23548 42000 23604
rect 0 23520 800 23548
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 41200 23520 42000 23548
rect 25218 23436 25228 23492
rect 25284 23436 26124 23492
rect 26180 23436 26190 23492
rect 31892 23436 37660 23492
rect 37716 23436 37726 23492
rect 15922 23324 15932 23380
rect 15988 23324 17724 23380
rect 17780 23324 17790 23380
rect 21634 23324 21644 23380
rect 21700 23324 22316 23380
rect 22372 23324 22382 23380
rect 31892 23268 31948 23436
rect 13906 23212 13916 23268
rect 13972 23212 17388 23268
rect 17444 23212 17454 23268
rect 19394 23212 19404 23268
rect 19460 23212 19470 23268
rect 26226 23212 26236 23268
rect 26292 23212 28140 23268
rect 28196 23212 31948 23268
rect 19404 23156 19460 23212
rect 15362 23100 15372 23156
rect 15428 23100 20188 23156
rect 20244 23100 20254 23156
rect 20514 23100 20524 23156
rect 20580 23100 21196 23156
rect 21252 23100 21756 23156
rect 21812 23100 21822 23156
rect 31892 23100 37660 23156
rect 37716 23100 37726 23156
rect 31892 23044 31948 23100
rect 13234 22988 13244 23044
rect 13300 22988 15260 23044
rect 15316 22988 16828 23044
rect 16884 22988 16894 23044
rect 18050 22988 18060 23044
rect 18116 22988 20412 23044
rect 20468 22988 22540 23044
rect 22596 22988 22606 23044
rect 25106 22988 25116 23044
rect 25172 22988 26012 23044
rect 26068 22988 26078 23044
rect 27122 22988 27132 23044
rect 27188 22988 29260 23044
rect 29316 22988 29326 23044
rect 31378 22988 31388 23044
rect 31444 22988 31948 23044
rect 41200 22932 42000 22960
rect 14018 22876 14028 22932
rect 14084 22876 17836 22932
rect 17892 22876 18956 22932
rect 19012 22876 19022 22932
rect 40002 22876 40012 22932
rect 40068 22876 42000 22932
rect 41200 22848 42000 22876
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 12786 22540 12796 22596
rect 12852 22540 21420 22596
rect 21476 22540 21486 22596
rect 28578 22428 28588 22484
rect 28644 22428 31388 22484
rect 31444 22428 31454 22484
rect 24770 22316 24780 22372
rect 24836 22316 26124 22372
rect 26180 22316 26190 22372
rect 27346 22316 27356 22372
rect 27412 22316 27422 22372
rect 27356 22260 27412 22316
rect 17266 22204 17276 22260
rect 17332 22204 18396 22260
rect 18452 22204 18462 22260
rect 21746 22204 21756 22260
rect 21812 22204 24108 22260
rect 24164 22204 25004 22260
rect 25060 22204 25070 22260
rect 27356 22204 27804 22260
rect 27860 22204 27870 22260
rect 27356 22148 27412 22204
rect 16370 22092 16380 22148
rect 16436 22092 19852 22148
rect 19908 22092 20524 22148
rect 20580 22092 22092 22148
rect 22148 22092 22158 22148
rect 22530 22092 22540 22148
rect 22596 22092 23100 22148
rect 23156 22092 23660 22148
rect 23716 22092 23726 22148
rect 23874 22092 23884 22148
rect 23940 22092 27412 22148
rect 27682 22092 27692 22148
rect 27748 22092 28476 22148
rect 28532 22092 28542 22148
rect 23314 21980 23324 22036
rect 23380 21980 27020 22036
rect 27076 21980 27086 22036
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 18386 21868 18396 21924
rect 18452 21868 19180 21924
rect 19236 21868 19246 21924
rect 26338 21868 26348 21924
rect 26404 21868 28140 21924
rect 28196 21868 28206 21924
rect 20738 21756 20748 21812
rect 20804 21756 21308 21812
rect 21364 21756 22988 21812
rect 23044 21756 23054 21812
rect 23202 21756 23212 21812
rect 23268 21756 24220 21812
rect 24276 21756 24286 21812
rect 17042 21644 17052 21700
rect 17108 21644 17724 21700
rect 17780 21644 17790 21700
rect 23090 21644 23100 21700
rect 23156 21644 26012 21700
rect 26068 21644 27020 21700
rect 27076 21644 27086 21700
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 16594 20972 16604 21028
rect 16660 20972 17164 21028
rect 17220 20972 22988 21028
rect 23044 20972 23054 21028
rect 41200 20916 42000 20944
rect 17602 20860 17612 20916
rect 17668 20860 18060 20916
rect 18116 20860 19852 20916
rect 19908 20860 19918 20916
rect 39890 20860 39900 20916
rect 39956 20860 42000 20916
rect 41200 20832 42000 20860
rect 14802 20748 14812 20804
rect 14868 20748 16380 20804
rect 16436 20748 16446 20804
rect 17836 20748 18508 20804
rect 18564 20748 19628 20804
rect 19684 20748 20300 20804
rect 20356 20748 20366 20804
rect 22194 20748 22204 20804
rect 22260 20748 23100 20804
rect 23156 20748 23166 20804
rect 17836 20692 17892 20748
rect 17826 20636 17836 20692
rect 17892 20636 17902 20692
rect 18834 20636 18844 20692
rect 18900 20636 20412 20692
rect 20468 20636 21532 20692
rect 21588 20636 21598 20692
rect 11666 20524 11676 20580
rect 11732 20524 15372 20580
rect 15428 20524 15438 20580
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 41200 20244 42000 20272
rect 40002 20188 40012 20244
rect 40068 20188 42000 20244
rect 41200 20160 42000 20188
rect 10098 20076 10108 20132
rect 10164 20076 11004 20132
rect 11060 20076 14252 20132
rect 14308 20076 15260 20132
rect 15316 20076 15326 20132
rect 21634 20076 21644 20132
rect 21700 20076 23772 20132
rect 23828 20076 23838 20132
rect 25666 20076 25676 20132
rect 25732 20076 26684 20132
rect 26740 20076 37884 20132
rect 37940 20076 37950 20132
rect 4162 19964 4172 20020
rect 4228 19964 19068 20020
rect 19124 19964 19516 20020
rect 19572 19964 19582 20020
rect 20178 19964 20188 20020
rect 20244 19964 21868 20020
rect 21924 19964 21934 20020
rect 13794 19852 13804 19908
rect 13860 19852 14812 19908
rect 14868 19852 14878 19908
rect 18498 19852 18508 19908
rect 18564 19852 18844 19908
rect 18900 19852 18910 19908
rect 24658 19852 24668 19908
rect 24724 19852 25340 19908
rect 25396 19852 25406 19908
rect 29698 19852 29708 19908
rect 29764 19852 37660 19908
rect 37716 19852 37726 19908
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 17378 19404 17388 19460
rect 17444 19404 21196 19460
rect 21252 19404 21262 19460
rect 27234 19404 27244 19460
rect 27300 19404 29148 19460
rect 29204 19404 29214 19460
rect 12898 19292 12908 19348
rect 12964 19292 14364 19348
rect 14420 19292 14430 19348
rect 19842 19292 19852 19348
rect 19908 19292 20188 19348
rect 20244 19292 21308 19348
rect 21364 19292 21374 19348
rect 22754 19292 22764 19348
rect 22820 19292 23548 19348
rect 23604 19292 23614 19348
rect 14802 19180 14812 19236
rect 14868 19180 15484 19236
rect 15540 19180 15550 19236
rect 17042 19180 17052 19236
rect 17108 19180 18284 19236
rect 18340 19180 24836 19236
rect 25890 19180 25900 19236
rect 25956 19180 27132 19236
rect 27188 19180 27198 19236
rect 24780 19124 24836 19180
rect 10770 19068 10780 19124
rect 10836 19068 13468 19124
rect 13524 19068 17948 19124
rect 18004 19068 20076 19124
rect 20132 19068 20142 19124
rect 21522 19068 21532 19124
rect 21588 19068 24556 19124
rect 24612 19068 24622 19124
rect 24780 19068 26796 19124
rect 26852 19068 27692 19124
rect 27748 19068 27758 19124
rect 16034 18956 16044 19012
rect 16100 18956 16940 19012
rect 16996 18956 19292 19012
rect 19348 18956 20580 19012
rect 22866 18956 22876 19012
rect 22932 18956 23436 19012
rect 23492 18956 23502 19012
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 20524 18788 20580 18956
rect 26852 18900 26908 19012
rect 26964 18956 26974 19012
rect 23874 18844 23884 18900
rect 23940 18844 26908 18900
rect 20514 18732 20524 18788
rect 20580 18732 21756 18788
rect 21812 18732 21822 18788
rect 15026 18620 15036 18676
rect 15092 18620 16268 18676
rect 16324 18620 16716 18676
rect 16772 18620 16782 18676
rect 18498 18396 18508 18452
rect 18564 18396 19404 18452
rect 19460 18396 22652 18452
rect 22708 18396 22718 18452
rect 24098 18396 24108 18452
rect 24164 18396 25228 18452
rect 25284 18396 25294 18452
rect 25778 18396 25788 18452
rect 25844 18396 26572 18452
rect 26628 18396 26638 18452
rect 27234 18396 27244 18452
rect 27300 18396 29148 18452
rect 29204 18396 29214 18452
rect 24546 18284 24556 18340
rect 24612 18284 25564 18340
rect 25620 18284 25630 18340
rect 41200 18228 42000 18256
rect 16258 18172 16268 18228
rect 16324 18172 17052 18228
rect 17108 18172 17118 18228
rect 40002 18172 40012 18228
rect 40068 18172 42000 18228
rect 41200 18144 42000 18172
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 14802 17948 14812 18004
rect 14868 17948 21308 18004
rect 21364 17948 21374 18004
rect 26002 17948 26012 18004
rect 26068 17948 26078 18004
rect 26012 17892 26068 17948
rect 20402 17836 20412 17892
rect 20468 17836 21868 17892
rect 21924 17836 21934 17892
rect 25218 17836 25228 17892
rect 25284 17836 26068 17892
rect 26012 17780 26068 17836
rect 18498 17724 18508 17780
rect 18564 17724 19852 17780
rect 19908 17724 20524 17780
rect 20580 17724 22428 17780
rect 22484 17724 22494 17780
rect 24434 17724 24444 17780
rect 24500 17724 25564 17780
rect 25620 17724 25630 17780
rect 26002 17724 26012 17780
rect 26068 17724 26078 17780
rect 17602 17612 17612 17668
rect 17668 17612 18844 17668
rect 18900 17612 18910 17668
rect 19506 17612 19516 17668
rect 19572 17612 20300 17668
rect 20356 17612 21532 17668
rect 21588 17612 24108 17668
rect 24164 17612 24174 17668
rect 25778 17612 25788 17668
rect 25844 17612 26348 17668
rect 26404 17612 26414 17668
rect 14914 17500 14924 17556
rect 14980 17500 16716 17556
rect 16772 17500 16782 17556
rect 23538 17500 23548 17556
rect 23604 17500 24332 17556
rect 24388 17500 25676 17556
rect 25732 17500 25742 17556
rect 29250 17500 29260 17556
rect 29316 17500 29708 17556
rect 29764 17500 37660 17556
rect 37716 17500 37726 17556
rect 16930 17388 16940 17444
rect 16996 17388 19516 17444
rect 19572 17388 23268 17444
rect 23426 17388 23436 17444
rect 23492 17388 25900 17444
rect 25956 17388 26908 17444
rect 23212 17332 23268 17388
rect 23212 17276 25228 17332
rect 25284 17276 25294 17332
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 21420 17164 21532 17220
rect 21588 17164 26236 17220
rect 26292 17164 26302 17220
rect 21420 17108 21476 17164
rect 26852 17108 26908 17388
rect 16482 17052 16492 17108
rect 16548 17052 17388 17108
rect 17444 17052 21476 17108
rect 21634 17052 21644 17108
rect 21700 17052 22876 17108
rect 22932 17052 22942 17108
rect 26114 17052 26124 17108
rect 26180 17052 26190 17108
rect 26852 17052 27020 17108
rect 27076 17052 27086 17108
rect 26124 16996 26180 17052
rect 13682 16940 13692 16996
rect 13748 16940 14588 16996
rect 14644 16940 14654 16996
rect 18722 16940 18732 16996
rect 18788 16940 20524 16996
rect 20580 16940 23604 16996
rect 24098 16940 24108 16996
rect 24164 16940 24556 16996
rect 24612 16940 24622 16996
rect 26124 16940 28588 16996
rect 28644 16940 31948 16996
rect 23548 16884 23604 16940
rect 31892 16884 31948 16940
rect 4274 16828 4284 16884
rect 4340 16828 12236 16884
rect 12292 16828 12302 16884
rect 12898 16828 12908 16884
rect 12964 16828 14252 16884
rect 14308 16828 16156 16884
rect 16212 16828 16222 16884
rect 16370 16828 16380 16884
rect 16436 16828 18284 16884
rect 18340 16828 18350 16884
rect 21858 16828 21868 16884
rect 21924 16828 23324 16884
rect 23380 16828 23390 16884
rect 23548 16828 24332 16884
rect 24388 16828 25116 16884
rect 25172 16828 25182 16884
rect 26898 16828 26908 16884
rect 26964 16828 29260 16884
rect 29316 16828 30156 16884
rect 30212 16828 30222 16884
rect 31892 16828 37660 16884
rect 37716 16828 37726 16884
rect 15698 16716 15708 16772
rect 15764 16716 17724 16772
rect 17780 16716 18172 16772
rect 18228 16716 18238 16772
rect 16258 16604 16268 16660
rect 16324 16604 20300 16660
rect 20356 16604 21644 16660
rect 21700 16604 22092 16660
rect 22148 16604 22158 16660
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 0 16212 800 16240
rect 41200 16212 42000 16240
rect 0 16156 1932 16212
rect 1988 16156 1998 16212
rect 40002 16156 40012 16212
rect 40068 16156 42000 16212
rect 0 16128 800 16156
rect 41200 16128 42000 16156
rect 12226 16044 12236 16100
rect 12292 16044 15820 16100
rect 15876 16044 15886 16100
rect 19842 16044 19852 16100
rect 19908 16044 20300 16100
rect 20356 16044 20366 16100
rect 14466 15932 14476 15988
rect 14532 15932 16604 15988
rect 16660 15932 16670 15988
rect 16818 15820 16828 15876
rect 16884 15820 17724 15876
rect 17780 15820 20076 15876
rect 20132 15820 22988 15876
rect 23044 15820 23054 15876
rect 25106 15820 25116 15876
rect 25172 15820 26348 15876
rect 26404 15820 26414 15876
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 17266 15596 17276 15652
rect 17332 15596 17342 15652
rect 17276 15540 17332 15596
rect 17276 15484 17500 15540
rect 17556 15484 17566 15540
rect 22978 15484 22988 15540
rect 23044 15484 25452 15540
rect 25508 15484 25518 15540
rect 14242 15372 14252 15428
rect 14308 15372 17556 15428
rect 17500 15204 17556 15372
rect 18162 15260 18172 15316
rect 18228 15260 19516 15316
rect 19572 15260 22652 15316
rect 22708 15260 22718 15316
rect 15484 15148 17276 15204
rect 17332 15148 17342 15204
rect 17500 15148 18956 15204
rect 19012 15148 19852 15204
rect 19908 15148 19918 15204
rect 15484 14980 15540 15148
rect 20132 15036 20188 15260
rect 22530 15148 22540 15204
rect 22596 15148 23884 15204
rect 23940 15148 23950 15204
rect 20244 15036 20254 15092
rect 15474 14924 15484 14980
rect 15540 14924 15550 14980
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 19058 14812 19068 14868
rect 19124 14812 19134 14868
rect 19068 14420 19124 14812
rect 20290 14476 20300 14532
rect 20356 14476 21196 14532
rect 21252 14476 21262 14532
rect 19068 14364 19292 14420
rect 19348 14364 21644 14420
rect 21700 14364 21710 14420
rect 15586 14252 15596 14308
rect 15652 14252 18060 14308
rect 18116 14252 18126 14308
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 19282 13804 19292 13860
rect 19348 13804 20524 13860
rect 20580 13804 20590 13860
rect 21858 13692 21868 13748
rect 21924 13692 23436 13748
rect 23492 13692 25340 13748
rect 25396 13692 25788 13748
rect 25844 13692 26796 13748
rect 26852 13692 26862 13748
rect 22978 13580 22988 13636
rect 23044 13580 24668 13636
rect 24724 13580 24734 13636
rect 18610 13468 18620 13524
rect 18676 13468 21084 13524
rect 21140 13468 21644 13524
rect 21700 13468 21710 13524
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 19506 13020 19516 13076
rect 19572 13020 20748 13076
rect 20804 13020 20814 13076
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 20850 4060 20860 4116
rect 20916 4060 22092 4116
rect 22148 4060 22158 4116
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 21522 3612 21532 3668
rect 21588 3612 22428 3668
rect 22484 3612 22494 3668
rect 24210 3612 24220 3668
rect 24276 3612 25564 3668
rect 25620 3612 25630 3668
rect 25554 3388 25564 3444
rect 25620 3388 26796 3444
rect 26852 3388 26862 3444
rect 16146 3276 16156 3332
rect 16212 3276 16940 3332
rect 16996 3276 17006 3332
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
<< via3 >>
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
<< metal4 >>
rect 4448 38444 4768 38476
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 37660 20128 38476
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19808 34524 20128 36036
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 19808 23548 20128 25060
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 19808 21980 20128 23492
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 38444 35488 38476
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _106_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 15344 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _107_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21840 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _108_
timestamp 1698175906
transform 1 0 14112 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _109_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21952 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _110_
timestamp 1698175906
transform 1 0 22960 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _111_
timestamp 1698175906
transform -1 0 18032 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _112_
timestamp 1698175906
transform 1 0 17808 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _113_
timestamp 1698175906
transform 1 0 18032 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _114_
timestamp 1698175906
transform -1 0 20720 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _115_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 20944 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _116_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 22512 0 1 21952
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _117_
timestamp 1698175906
transform 1 0 17248 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _118_
timestamp 1698175906
transform 1 0 17360 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _119_
timestamp 1698175906
transform 1 0 19712 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _120_
timestamp 1698175906
transform 1 0 16128 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _121_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 16352 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _122_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18256 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _123_
timestamp 1698175906
transform 1 0 25088 0 -1 20384
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _124_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21168 0 1 20384
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _125_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 20720 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _126_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 24752 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _127_
timestamp 1698175906
transform -1 0 20048 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _128_
timestamp 1698175906
transform -1 0 25424 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _129_
timestamp 1698175906
transform 1 0 21168 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _130_
timestamp 1698175906
transform -1 0 24864 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _131_
timestamp 1698175906
transform 1 0 14560 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _132_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 15680 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _133_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 15344 0 -1 20384
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _134_
timestamp 1698175906
transform -1 0 14000 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _135_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18704 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _136_
timestamp 1698175906
transform -1 0 16576 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _137_
timestamp 1698175906
transform -1 0 17248 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _138_
timestamp 1698175906
transform -1 0 15120 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _139_
timestamp 1698175906
transform 1 0 19600 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _140_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 22960 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _141_
timestamp 1698175906
transform -1 0 23184 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _142_
timestamp 1698175906
transform 1 0 17920 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _143_
timestamp 1698175906
transform -1 0 17808 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _144_
timestamp 1698175906
transform -1 0 18256 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _145_
timestamp 1698175906
transform 1 0 18144 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _146_
timestamp 1698175906
transform -1 0 19152 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _147_
timestamp 1698175906
transform -1 0 18368 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _148_
timestamp 1698175906
transform 1 0 17808 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _149_
timestamp 1698175906
transform -1 0 19712 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _150_
timestamp 1698175906
transform 1 0 18816 0 -1 23520
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _151_
timestamp 1698175906
transform 1 0 19264 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _152_
timestamp 1698175906
transform -1 0 20048 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _153_
timestamp 1698175906
transform 1 0 22736 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _154_
timestamp 1698175906
transform 1 0 19040 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _155_
timestamp 1698175906
transform -1 0 24752 0 1 17248
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _156_
timestamp 1698175906
transform 1 0 18704 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _157_
timestamp 1698175906
transform -1 0 24192 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _158_
timestamp 1698175906
transform -1 0 16688 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _159_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 17696 0 1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _160_
timestamp 1698175906
transform -1 0 16016 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _161_
timestamp 1698175906
transform -1 0 14784 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _162_
timestamp 1698175906
transform -1 0 14448 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _163_
timestamp 1698175906
transform 1 0 16576 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _164_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 18144 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _165_
timestamp 1698175906
transform 1 0 22400 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _166_
timestamp 1698175906
transform 1 0 22960 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _167_
timestamp 1698175906
transform -1 0 29456 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _168_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 26208 0 -1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _169_
timestamp 1698175906
transform 1 0 25872 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _170_
timestamp 1698175906
transform 1 0 25424 0 -1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _171_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17472 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _172_
timestamp 1698175906
transform -1 0 19488 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _173_
timestamp 1698175906
transform -1 0 16688 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _174_
timestamp 1698175906
transform 1 0 21392 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _175_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 15680 0 1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _176_
timestamp 1698175906
transform -1 0 14672 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _177_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 22848 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _178_
timestamp 1698175906
transform 1 0 25872 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _179_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21168 0 1 17248
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _180_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 24416 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _181_
timestamp 1698175906
transform -1 0 29456 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _182_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 26208 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _183_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 23744 0 -1 18816
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _184_
timestamp 1698175906
transform 1 0 26880 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _185_
timestamp 1698175906
transform -1 0 20608 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _186_
timestamp 1698175906
transform 1 0 19152 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _187_
timestamp 1698175906
transform -1 0 20384 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _188_
timestamp 1698175906
transform -1 0 20272 0 -1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _189_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19712 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _190_
timestamp 1698175906
transform -1 0 21840 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _191_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19824 0 1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _192_
timestamp 1698175906
transform -1 0 28784 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _193_
timestamp 1698175906
transform -1 0 27888 0 1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _194_
timestamp 1698175906
transform -1 0 13888 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _195_
timestamp 1698175906
transform -1 0 21952 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _196_
timestamp 1698175906
transform -1 0 12992 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _197_
timestamp 1698175906
transform -1 0 22736 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _198_
timestamp 1698175906
transform 1 0 17696 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _199_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18368 0 1 23520
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _200_
timestamp 1698175906
transform 1 0 21168 0 1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _201_
timestamp 1698175906
transform 1 0 13328 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _202_
timestamp 1698175906
transform -1 0 12992 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _203_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17248 0 -1 23520
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _204_
timestamp 1698175906
transform 1 0 15792 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _205_
timestamp 1698175906
transform 1 0 23296 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _206_
timestamp 1698175906
transform 1 0 23856 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _207_
timestamp 1698175906
transform 1 0 23408 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _208_
timestamp 1698175906
transform -1 0 22624 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _209_
timestamp 1698175906
transform 1 0 19712 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _210_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 20720 0 -1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _211_
timestamp 1698175906
transform 1 0 21168 0 1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _212_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 23632 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _213_
timestamp 1698175906
transform 1 0 23296 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _214_
timestamp 1698175906
transform 1 0 10752 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _215_
timestamp 1698175906
transform 1 0 9856 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _216_
timestamp 1698175906
transform 1 0 12656 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _217_
timestamp 1698175906
transform 1 0 14560 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _218_
timestamp 1698175906
transform 1 0 16240 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _219_
timestamp 1698175906
transform 1 0 17248 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _220_
timestamp 1698175906
transform 1 0 21616 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _221_
timestamp 1698175906
transform 1 0 13776 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _222_
timestamp 1698175906
transform -1 0 15232 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _223_
timestamp 1698175906
transform 1 0 26656 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _224_
timestamp 1698175906
transform 1 0 25536 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _225_
timestamp 1698175906
transform -1 0 15344 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _226_
timestamp 1698175906
transform 1 0 25088 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _227_
timestamp 1698175906
transform 1 0 26656 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _228_
timestamp 1698175906
transform 1 0 17696 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _229_
timestamp 1698175906
transform 1 0 18368 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _230_
timestamp 1698175906
transform 1 0 28336 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _231_
timestamp 1698175906
transform -1 0 13664 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _232_
timestamp 1698175906
transform 1 0 20720 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _233_
timestamp 1698175906
transform -1 0 13104 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _234_
timestamp 1698175906
transform -1 0 17024 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _235_
timestamp 1698175906
transform 1 0 22624 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _236_
timestamp 1698175906
transform -1 0 23296 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _241_
timestamp 1698175906
transform -1 0 24640 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__212__CLK dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 27104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__213__CLK
timestamp 1698175906
transform 1 0 26768 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__214__CLK
timestamp 1698175906
transform 1 0 14224 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__215__CLK
timestamp 1698175906
transform 1 0 13104 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__216__CLK
timestamp 1698175906
transform 1 0 16128 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__217__CLK
timestamp 1698175906
transform 1 0 18032 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__218__CLK
timestamp 1698175906
transform 1 0 19488 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__219__CLK
timestamp 1698175906
transform 1 0 20496 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__220__CLK
timestamp 1698175906
transform 1 0 25312 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__221__CLK
timestamp 1698175906
transform 1 0 17472 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__222__CLK
timestamp 1698175906
transform -1 0 15680 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__223__CLK
timestamp 1698175906
transform 1 0 30128 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__224__CLK
timestamp 1698175906
transform 1 0 29232 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__225__CLK
timestamp 1698175906
transform 1 0 15568 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__226__CLK
timestamp 1698175906
transform 1 0 28336 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__227__CLK
timestamp 1698175906
transform 1 0 30128 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__228__CLK
timestamp 1698175906
transform -1 0 21168 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__229__CLK
timestamp 1698175906
transform 1 0 21616 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__230__CLK
timestamp 1698175906
transform 1 0 28112 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__231__CLK
timestamp 1698175906
transform 1 0 13888 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__232__CLK
timestamp 1698175906
transform 1 0 23968 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__233__CLK
timestamp 1698175906
transform 1 0 13216 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__234__CLK
timestamp 1698175906
transform 1 0 17024 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__235__CLK
timestamp 1698175906
transform 1 0 26096 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__236__CLK
timestamp 1698175906
transform 1 0 23520 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1698175906
transform 1 0 19040 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19264 0 -1 20384
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1698175906
transform -1 0 22848 0 -1 21952
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1698175906
transform 1 0 23072 0 1 20384
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1568 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698175906
transform 1 0 5376 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698175906
transform 1 0 9184 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698175906
transform 1 0 12992 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_142 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17248 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_158 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19040 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_166 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19936 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_172
timestamp 1698175906
transform 1 0 20608 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_176 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21056 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_232
timestamp 1698175906
transform 1 0 27328 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_236
timestamp 1698175906
transform 1 0 27776 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_240
timestamp 1698175906
transform 1 0 28224 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_274
timestamp 1698175906
transform 1 0 32032 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_308
timestamp 1698175906
transform 1 0 35840 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_342
timestamp 1698175906
transform 1 0 39648 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_346
timestamp 1698175906
transform 1 0 40096 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_348 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 40320 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1568 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698175906
transform 1 0 8736 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698175906
transform 1 0 9408 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698175906
transform 1 0 16576 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_142
timestamp 1698175906
transform 1 0 17248 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_174
timestamp 1698175906
transform 1 0 20832 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_201
timestamp 1698175906
transform 1 0 23856 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_209
timestamp 1698175906
transform 1 0 24752 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_212
timestamp 1698175906
transform 1 0 25088 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_216
timestamp 1698175906
transform 1 0 25536 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_243
timestamp 1698175906
transform 1 0 28560 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_275
timestamp 1698175906
transform 1 0 32144 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_279
timestamp 1698175906
transform 1 0 32592 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_282
timestamp 1698175906
transform 1 0 32928 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_346
timestamp 1698175906
transform 1 0 40096 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_348
timestamp 1698175906
transform 1 0 40320 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698175906
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698175906
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698175906
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698175906
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_107
timestamp 1698175906
transform 1 0 13328 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_171
timestamp 1698175906
transform 1 0 20496 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_177
timestamp 1698175906
transform 1 0 21168 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_241
timestamp 1698175906
transform 1 0 28336 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698175906
transform 1 0 29008 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698175906
transform 1 0 36176 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_317
timestamp 1698175906
transform 1 0 36848 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698175906
transform 1 0 1568 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698175906
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698175906
transform 1 0 9408 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698175906
transform 1 0 16576 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_142
timestamp 1698175906
transform 1 0 17248 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_206
timestamp 1698175906
transform 1 0 24416 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_212
timestamp 1698175906
transform 1 0 25088 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_276
timestamp 1698175906
transform 1 0 32256 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_282
timestamp 1698175906
transform 1 0 32928 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_346
timestamp 1698175906
transform 1 0 40096 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_348
timestamp 1698175906
transform 1 0 40320 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698175906
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698175906
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698175906
transform 1 0 5488 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698175906
transform 1 0 12656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_107
timestamp 1698175906
transform 1 0 13328 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698175906
transform 1 0 20496 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_177
timestamp 1698175906
transform 1 0 21168 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_241
timestamp 1698175906
transform 1 0 28336 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698175906
transform 1 0 29008 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698175906
transform 1 0 36176 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_317
timestamp 1698175906
transform 1 0 36848 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698175906
transform 1 0 1568 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698175906
transform 1 0 8736 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698175906
transform 1 0 9408 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698175906
transform 1 0 16576 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_142
timestamp 1698175906
transform 1 0 17248 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_206
timestamp 1698175906
transform 1 0 24416 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_212
timestamp 1698175906
transform 1 0 25088 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698175906
transform 1 0 32256 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_282
timestamp 1698175906
transform 1 0 32928 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_346
timestamp 1698175906
transform 1 0 40096 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_348
timestamp 1698175906
transform 1 0 40320 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698175906
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698175906
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698175906
transform 1 0 5488 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698175906
transform 1 0 12656 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_107
timestamp 1698175906
transform 1 0 13328 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_171
timestamp 1698175906
transform 1 0 20496 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_177
timestamp 1698175906
transform 1 0 21168 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_241
timestamp 1698175906
transform 1 0 28336 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_247
timestamp 1698175906
transform 1 0 29008 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_311
timestamp 1698175906
transform 1 0 36176 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_317
timestamp 1698175906
transform 1 0 36848 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698175906
transform 1 0 1568 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698175906
transform 1 0 8736 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_72
timestamp 1698175906
transform 1 0 9408 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698175906
transform 1 0 16576 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_142
timestamp 1698175906
transform 1 0 17248 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_206
timestamp 1698175906
transform 1 0 24416 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_212
timestamp 1698175906
transform 1 0 25088 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_276
timestamp 1698175906
transform 1 0 32256 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_282
timestamp 1698175906
transform 1 0 32928 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_346
timestamp 1698175906
transform 1 0 40096 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_348
timestamp 1698175906
transform 1 0 40320 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698175906
transform 1 0 1568 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698175906
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_37
timestamp 1698175906
transform 1 0 5488 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_101
timestamp 1698175906
transform 1 0 12656 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_107
timestamp 1698175906
transform 1 0 13328 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_171
timestamp 1698175906
transform 1 0 20496 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_177
timestamp 1698175906
transform 1 0 21168 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_241
timestamp 1698175906
transform 1 0 28336 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_247
timestamp 1698175906
transform 1 0 29008 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_311
timestamp 1698175906
transform 1 0 36176 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_317
timestamp 1698175906
transform 1 0 36848 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698175906
transform 1 0 1568 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698175906
transform 1 0 8736 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_72
timestamp 1698175906
transform 1 0 9408 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_136
timestamp 1698175906
transform 1 0 16576 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_142
timestamp 1698175906
transform 1 0 17248 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_206
timestamp 1698175906
transform 1 0 24416 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_212
timestamp 1698175906
transform 1 0 25088 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_276
timestamp 1698175906
transform 1 0 32256 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_282
timestamp 1698175906
transform 1 0 32928 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_346
timestamp 1698175906
transform 1 0 40096 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_348
timestamp 1698175906
transform 1 0 40320 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698175906
transform 1 0 1568 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698175906
transform 1 0 5152 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_37
timestamp 1698175906
transform 1 0 5488 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698175906
transform 1 0 12656 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_107
timestamp 1698175906
transform 1 0 13328 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_171
timestamp 1698175906
transform 1 0 20496 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_177
timestamp 1698175906
transform 1 0 21168 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_241
timestamp 1698175906
transform 1 0 28336 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_247
timestamp 1698175906
transform 1 0 29008 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_311
timestamp 1698175906
transform 1 0 36176 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_317
timestamp 1698175906
transform 1 0 36848 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2
timestamp 1698175906
transform 1 0 1568 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698175906
transform 1 0 8736 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_72
timestamp 1698175906
transform 1 0 9408 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698175906
transform 1 0 16576 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_11_142
timestamp 1698175906
transform 1 0 17248 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_174
timestamp 1698175906
transform 1 0 20832 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_11_177
timestamp 1698175906
transform 1 0 21168 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_209
timestamp 1698175906
transform 1 0 24752 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_212
timestamp 1698175906
transform 1 0 25088 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_276
timestamp 1698175906
transform 1 0 32256 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_282
timestamp 1698175906
transform 1 0 32928 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_346
timestamp 1698175906
transform 1 0 40096 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_348
timestamp 1698175906
transform 1 0 40320 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698175906
transform 1 0 1568 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698175906
transform 1 0 5152 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_37
timestamp 1698175906
transform 1 0 5488 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698175906
transform 1 0 12656 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_107
timestamp 1698175906
transform 1 0 13328 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_139
timestamp 1698175906
transform 1 0 16912 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_143
timestamp 1698175906
transform 1 0 17360 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_145
timestamp 1698175906
transform 1 0 17584 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_177
timestamp 1698175906
transform 1 0 21168 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_183
timestamp 1698175906
transform 1 0 21840 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_215
timestamp 1698175906
transform 1 0 25424 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_231
timestamp 1698175906
transform 1 0 27216 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_239
timestamp 1698175906
transform 1 0 28112 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_243
timestamp 1698175906
transform 1 0 28560 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_247
timestamp 1698175906
transform 1 0 29008 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_311
timestamp 1698175906
transform 1 0 36176 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_317
timestamp 1698175906
transform 1 0 36848 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_2
timestamp 1698175906
transform 1 0 1568 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_66
timestamp 1698175906
transform 1 0 8736 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_72
timestamp 1698175906
transform 1 0 9408 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_136
timestamp 1698175906
transform 1 0 16576 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_142
timestamp 1698175906
transform 1 0 17248 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_150
timestamp 1698175906
transform 1 0 18144 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_212
timestamp 1698175906
transform 1 0 25088 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_216
timestamp 1698175906
transform 1 0 25536 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_282
timestamp 1698175906
transform 1 0 32928 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_346
timestamp 1698175906
transform 1 0 40096 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_348
timestamp 1698175906
transform 1 0 40320 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698175906
transform 1 0 1568 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698175906
transform 1 0 5152 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_37
timestamp 1698175906
transform 1 0 5488 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_101
timestamp 1698175906
transform 1 0 12656 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_107
timestamp 1698175906
transform 1 0 13328 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_115
timestamp 1698175906
transform 1 0 14224 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_117
timestamp 1698175906
transform 1 0 14448 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_147
timestamp 1698175906
transform 1 0 17808 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_151
timestamp 1698175906
transform 1 0 18256 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_183
timestamp 1698175906
transform 1 0 21840 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_225
timestamp 1698175906
transform 1 0 26544 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_229
timestamp 1698175906
transform 1 0 26992 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_247
timestamp 1698175906
transform 1 0 29008 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_311
timestamp 1698175906
transform 1 0 36176 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_317
timestamp 1698175906
transform 1 0 36848 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_2
timestamp 1698175906
transform 1 0 1568 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_66
timestamp 1698175906
transform 1 0 8736 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_72
timestamp 1698175906
transform 1 0 9408 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_88
timestamp 1698175906
transform 1 0 11200 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_125
timestamp 1698175906
transform 1 0 15344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_129
timestamp 1698175906
transform 1 0 15792 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_137
timestamp 1698175906
transform 1 0 16688 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_139
timestamp 1698175906
transform 1 0 16912 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_147
timestamp 1698175906
transform 1 0 17808 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_155
timestamp 1698175906
transform 1 0 18704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_169
timestamp 1698175906
transform 1 0 20272 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_185
timestamp 1698175906
transform 1 0 22064 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_195
timestamp 1698175906
transform 1 0 23184 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_204
timestamp 1698175906
transform 1 0 24192 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_208
timestamp 1698175906
transform 1 0 24640 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_212
timestamp 1698175906
transform 1 0 25088 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_276
timestamp 1698175906
transform 1 0 32256 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_282
timestamp 1698175906
transform 1 0 32928 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_346
timestamp 1698175906
transform 1 0 40096 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_348
timestamp 1698175906
transform 1 0 40320 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_2
timestamp 1698175906
transform 1 0 1568 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698175906
transform 1 0 5152 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_37
timestamp 1698175906
transform 1 0 5488 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_101
timestamp 1698175906
transform 1 0 12656 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_107
timestamp 1698175906
transform 1 0 13328 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_111
timestamp 1698175906
transform 1 0 13776 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_119
timestamp 1698175906
transform 1 0 14672 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_127
timestamp 1698175906
transform 1 0 15568 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_140
timestamp 1698175906
transform 1 0 17024 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_153
timestamp 1698175906
transform 1 0 18480 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_161
timestamp 1698175906
transform 1 0 19376 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_170
timestamp 1698175906
transform 1 0 20384 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_174
timestamp 1698175906
transform 1 0 20832 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_177
timestamp 1698175906
transform 1 0 21168 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_209
timestamp 1698175906
transform 1 0 24752 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_215
timestamp 1698175906
transform 1 0 25424 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_247
timestamp 1698175906
transform 1 0 29008 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_251
timestamp 1698175906
transform 1 0 29456 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_317
timestamp 1698175906
transform 1 0 36848 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_28
timestamp 1698175906
transform 1 0 4480 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_60
timestamp 1698175906
transform 1 0 8064 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_68
timestamp 1698175906
transform 1 0 8960 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_72
timestamp 1698175906
transform 1 0 9408 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_88
timestamp 1698175906
transform 1 0 11200 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_96
timestamp 1698175906
transform 1 0 12096 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_100
timestamp 1698175906
transform 1 0 12544 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_130
timestamp 1698175906
transform 1 0 15904 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_134
timestamp 1698175906
transform 1 0 16352 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_138
timestamp 1698175906
transform 1 0 16800 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_150
timestamp 1698175906
transform 1 0 18144 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_158
timestamp 1698175906
transform 1 0 19040 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_162
timestamp 1698175906
transform 1 0 19488 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_172
timestamp 1698175906
transform 1 0 20608 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_176
timestamp 1698175906
transform 1 0 21056 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_178
timestamp 1698175906
transform 1 0 21280 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_184
timestamp 1698175906
transform 1 0 21952 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_200
timestamp 1698175906
transform 1 0 23744 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_212
timestamp 1698175906
transform 1 0 25088 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_214
timestamp 1698175906
transform 1 0 25312 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_224
timestamp 1698175906
transform 1 0 26432 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_255
timestamp 1698175906
transform 1 0 29904 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_259
timestamp 1698175906
transform 1 0 30352 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_275
timestamp 1698175906
transform 1 0 32144 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_279
timestamp 1698175906
transform 1 0 32592 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_282
timestamp 1698175906
transform 1 0 32928 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_314
timestamp 1698175906
transform 1 0 36512 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_322
timestamp 1698175906
transform 1 0 37408 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_2
timestamp 1698175906
transform 1 0 1568 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698175906
transform 1 0 5152 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_37
timestamp 1698175906
transform 1 0 5488 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_101
timestamp 1698175906
transform 1 0 12656 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_107
timestamp 1698175906
transform 1 0 13328 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_115
timestamp 1698175906
transform 1 0 14224 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_117
timestamp 1698175906
transform 1 0 14448 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_123
timestamp 1698175906
transform 1 0 15120 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_142
timestamp 1698175906
transform 1 0 17248 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_146
timestamp 1698175906
transform 1 0 17696 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_148
timestamp 1698175906
transform 1 0 17920 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_173
timestamp 1698175906
transform 1 0 20720 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_199
timestamp 1698175906
transform 1 0 23632 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_201
timestamp 1698175906
transform 1 0 23856 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_209
timestamp 1698175906
transform 1 0 24752 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_217
timestamp 1698175906
transform 1 0 25648 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_224
timestamp 1698175906
transform 1 0 26432 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_240
timestamp 1698175906
transform 1 0 28224 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_244
timestamp 1698175906
transform 1 0 28672 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_251
timestamp 1698175906
transform 1 0 29456 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_317
timestamp 1698175906
transform 1 0 36848 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_2
timestamp 1698175906
transform 1 0 1568 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_66
timestamp 1698175906
transform 1 0 8736 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_72
timestamp 1698175906
transform 1 0 9408 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_104
timestamp 1698175906
transform 1 0 12992 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_107
timestamp 1698175906
transform 1 0 13328 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_123
timestamp 1698175906
transform 1 0 15120 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_136
timestamp 1698175906
transform 1 0 16576 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_142
timestamp 1698175906
transform 1 0 17248 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_200
timestamp 1698175906
transform 1 0 23744 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_208
timestamp 1698175906
transform 1 0 24640 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_234
timestamp 1698175906
transform 1 0 27552 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_266
timestamp 1698175906
transform 1 0 31136 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_274
timestamp 1698175906
transform 1 0 32032 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_278
timestamp 1698175906
transform 1 0 32480 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_282
timestamp 1698175906
transform 1 0 32928 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_314
timestamp 1698175906
transform 1 0 36512 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_322
timestamp 1698175906
transform 1 0 37408 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_2
timestamp 1698175906
transform 1 0 1568 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698175906
transform 1 0 5152 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_37
timestamp 1698175906
transform 1 0 5488 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_69
timestamp 1698175906
transform 1 0 9072 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_73
timestamp 1698175906
transform 1 0 9520 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_75
timestamp 1698175906
transform 1 0 9744 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_113
timestamp 1698175906
transform 1 0 14000 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_117
timestamp 1698175906
transform 1 0 14448 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_124
timestamp 1698175906
transform 1 0 15232 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_133
timestamp 1698175906
transform 1 0 16240 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_135
timestamp 1698175906
transform 1 0 16464 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_142
timestamp 1698175906
transform 1 0 17248 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_144
timestamp 1698175906
transform 1 0 17472 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_149
timestamp 1698175906
transform 1 0 18032 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_157
timestamp 1698175906
transform 1 0 18928 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_172
timestamp 1698175906
transform 1 0 20608 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_174
timestamp 1698175906
transform 1 0 20832 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_228
timestamp 1698175906
transform 1 0 26880 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_232
timestamp 1698175906
transform 1 0 27328 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_240
timestamp 1698175906
transform 1 0 28224 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_244
timestamp 1698175906
transform 1 0 28672 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_251
timestamp 1698175906
transform 1 0 29456 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_317
timestamp 1698175906
transform 1 0 36848 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_2
timestamp 1698175906
transform 1 0 1568 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_66
timestamp 1698175906
transform 1 0 8736 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_72
timestamp 1698175906
transform 1 0 9408 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_80
timestamp 1698175906
transform 1 0 10304 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_125
timestamp 1698175906
transform 1 0 15344 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_129
timestamp 1698175906
transform 1 0 15792 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_131
timestamp 1698175906
transform 1 0 16016 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_142
timestamp 1698175906
transform 1 0 17248 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_146
timestamp 1698175906
transform 1 0 17696 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_155
timestamp 1698175906
transform 1 0 18704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_157
timestamp 1698175906
transform 1 0 18928 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_219
timestamp 1698175906
transform 1 0 25872 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_223
timestamp 1698175906
transform 1 0 26320 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_225
timestamp 1698175906
transform 1 0 26544 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_255
timestamp 1698175906
transform 1 0 29904 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_259
timestamp 1698175906
transform 1 0 30352 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_275
timestamp 1698175906
transform 1 0 32144 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_279
timestamp 1698175906
transform 1 0 32592 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_282
timestamp 1698175906
transform 1 0 32928 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_346
timestamp 1698175906
transform 1 0 40096 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_348
timestamp 1698175906
transform 1 0 40320 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_2
timestamp 1698175906
transform 1 0 1568 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698175906
transform 1 0 5152 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_37
timestamp 1698175906
transform 1 0 5488 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_101
timestamp 1698175906
transform 1 0 12656 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_107
timestamp 1698175906
transform 1 0 13328 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_111
timestamp 1698175906
transform 1 0 13776 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_113
timestamp 1698175906
transform 1 0 14000 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_122
timestamp 1698175906
transform 1 0 15008 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_128
timestamp 1698175906
transform 1 0 15680 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_132
timestamp 1698175906
transform 1 0 16128 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_172
timestamp 1698175906
transform 1 0 20608 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_174
timestamp 1698175906
transform 1 0 20832 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_191
timestamp 1698175906
transform 1 0 22736 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_193
timestamp 1698175906
transform 1 0 22960 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_244
timestamp 1698175906
transform 1 0 28672 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_247
timestamp 1698175906
transform 1 0 29008 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_311
timestamp 1698175906
transform 1 0 36176 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_317
timestamp 1698175906
transform 1 0 36848 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_321
timestamp 1698175906
transform 1 0 37296 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_2
timestamp 1698175906
transform 1 0 1568 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_66
timestamp 1698175906
transform 1 0 8736 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_72
timestamp 1698175906
transform 1 0 9408 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_136
timestamp 1698175906
transform 1 0 16576 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_200
timestamp 1698175906
transform 1 0 23744 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_209
timestamp 1698175906
transform 1 0 24752 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_212
timestamp 1698175906
transform 1 0 25088 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_238
timestamp 1698175906
transform 1 0 28000 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_270
timestamp 1698175906
transform 1 0 31584 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_278
timestamp 1698175906
transform 1 0 32480 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_282
timestamp 1698175906
transform 1 0 32928 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_314
timestamp 1698175906
transform 1 0 36512 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_322
timestamp 1698175906
transform 1 0 37408 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_2
timestamp 1698175906
transform 1 0 1568 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698175906
transform 1 0 5152 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_37
timestamp 1698175906
transform 1 0 5488 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_101
timestamp 1698175906
transform 1 0 12656 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_107
timestamp 1698175906
transform 1 0 13328 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_123
timestamp 1698175906
transform 1 0 15120 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_127
timestamp 1698175906
transform 1 0 15568 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_133
timestamp 1698175906
transform 1 0 16240 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_137
timestamp 1698175906
transform 1 0 16688 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_139
timestamp 1698175906
transform 1 0 16912 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_142
timestamp 1698175906
transform 1 0 17248 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_144
timestamp 1698175906
transform 1 0 17472 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_162
timestamp 1698175906
transform 1 0 19488 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_204
timestamp 1698175906
transform 1 0 24192 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_214
timestamp 1698175906
transform 1 0 25312 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_218
timestamp 1698175906
transform 1 0 25760 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_225
timestamp 1698175906
transform 1 0 26544 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_237
timestamp 1698175906
transform 1 0 27888 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_247
timestamp 1698175906
transform 1 0 29008 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_311
timestamp 1698175906
transform 1 0 36176 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_317
timestamp 1698175906
transform 1 0 36848 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_2
timestamp 1698175906
transform 1 0 1568 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_66
timestamp 1698175906
transform 1 0 8736 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_72
timestamp 1698175906
transform 1 0 9408 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_88
timestamp 1698175906
transform 1 0 11200 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_96
timestamp 1698175906
transform 1 0 12096 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_98
timestamp 1698175906
transform 1 0 12320 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_104
timestamp 1698175906
transform 1 0 12992 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_108
timestamp 1698175906
transform 1 0 13440 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_110
timestamp 1698175906
transform 1 0 13664 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_153
timestamp 1698175906
transform 1 0 18480 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_155
timestamp 1698175906
transform 1 0 18704 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_188
timestamp 1698175906
transform 1 0 22400 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_196
timestamp 1698175906
transform 1 0 23296 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_205
timestamp 1698175906
transform 1 0 24304 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_209
timestamp 1698175906
transform 1 0 24752 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_270
timestamp 1698175906
transform 1 0 31584 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_278
timestamp 1698175906
transform 1 0 32480 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_282
timestamp 1698175906
transform 1 0 32928 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_314
timestamp 1698175906
transform 1 0 36512 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_322
timestamp 1698175906
transform 1 0 37408 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_28
timestamp 1698175906
transform 1 0 4480 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_32
timestamp 1698175906
transform 1 0 4928 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698175906
transform 1 0 5152 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_37
timestamp 1698175906
transform 1 0 5488 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_69
timestamp 1698175906
transform 1 0 9072 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_73
timestamp 1698175906
transform 1 0 9520 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_75
timestamp 1698175906
transform 1 0 9744 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_115
timestamp 1698175906
transform 1 0 14224 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_131
timestamp 1698175906
transform 1 0 16016 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_139
timestamp 1698175906
transform 1 0 16912 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_143
timestamp 1698175906
transform 1 0 17360 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_145
timestamp 1698175906
transform 1 0 17584 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_177
timestamp 1698175906
transform 1 0 21168 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_185
timestamp 1698175906
transform 1 0 22064 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_189
timestamp 1698175906
transform 1 0 22512 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_219
timestamp 1698175906
transform 1 0 25872 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_223
timestamp 1698175906
transform 1 0 26320 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_239
timestamp 1698175906
transform 1 0 28112 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_243
timestamp 1698175906
transform 1 0 28560 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_247
timestamp 1698175906
transform 1 0 29008 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_311
timestamp 1698175906
transform 1 0 36176 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_317
timestamp 1698175906
transform 1 0 36848 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_321
timestamp 1698175906
transform 1 0 37296 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_28
timestamp 1698175906
transform 1 0 4480 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_60
timestamp 1698175906
transform 1 0 8064 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_68
timestamp 1698175906
transform 1 0 8960 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_72
timestamp 1698175906
transform 1 0 9408 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_80
timestamp 1698175906
transform 1 0 10304 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_110
timestamp 1698175906
transform 1 0 13664 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_114
timestamp 1698175906
transform 1 0 14112 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_130
timestamp 1698175906
transform 1 0 15904 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_138
timestamp 1698175906
transform 1 0 16800 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_142
timestamp 1698175906
transform 1 0 17248 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_158
timestamp 1698175906
transform 1 0 19040 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_162
timestamp 1698175906
transform 1 0 19488 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_169
timestamp 1698175906
transform 1 0 20272 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_206
timestamp 1698175906
transform 1 0 24416 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_212
timestamp 1698175906
transform 1 0 25088 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_276
timestamp 1698175906
transform 1 0 32256 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_282
timestamp 1698175906
transform 1 0 32928 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_314
timestamp 1698175906
transform 1 0 36512 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_322
timestamp 1698175906
transform 1 0 37408 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_28
timestamp 1698175906
transform 1 0 4480 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_32
timestamp 1698175906
transform 1 0 4928 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698175906
transform 1 0 5152 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_37
timestamp 1698175906
transform 1 0 5488 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_69
timestamp 1698175906
transform 1 0 9072 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_85
timestamp 1698175906
transform 1 0 10864 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_93
timestamp 1698175906
transform 1 0 11760 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_97
timestamp 1698175906
transform 1 0 12208 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_104
timestamp 1698175906
transform 1 0 12992 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_112
timestamp 1698175906
transform 1 0 13888 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_114
timestamp 1698175906
transform 1 0 14112 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_120
timestamp 1698175906
transform 1 0 14784 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_124
timestamp 1698175906
transform 1 0 15232 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_126
timestamp 1698175906
transform 1 0 15456 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_146
timestamp 1698175906
transform 1 0 17696 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_156
timestamp 1698175906
transform 1 0 18816 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_172
timestamp 1698175906
transform 1 0 20608 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_174
timestamp 1698175906
transform 1 0 20832 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_190
timestamp 1698175906
transform 1 0 22624 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_222
timestamp 1698175906
transform 1 0 26208 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_238
timestamp 1698175906
transform 1 0 28000 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_242
timestamp 1698175906
transform 1 0 28448 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_244
timestamp 1698175906
transform 1 0 28672 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_247
timestamp 1698175906
transform 1 0 29008 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_311
timestamp 1698175906
transform 1 0 36176 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_317
timestamp 1698175906
transform 1 0 36848 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_2
timestamp 1698175906
transform 1 0 1568 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_66
timestamp 1698175906
transform 1 0 8736 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_72
timestamp 1698175906
transform 1 0 9408 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_104
timestamp 1698175906
transform 1 0 12992 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_108
timestamp 1698175906
transform 1 0 13440 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_110
timestamp 1698175906
transform 1 0 13664 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_142
timestamp 1698175906
transform 1 0 17248 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_146
timestamp 1698175906
transform 1 0 17696 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_164
timestamp 1698175906
transform 1 0 19712 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_166
timestamp 1698175906
transform 1 0 19936 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_196
timestamp 1698175906
transform 1 0 23296 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_200
timestamp 1698175906
transform 1 0 23744 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_208
timestamp 1698175906
transform 1 0 24640 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_212
timestamp 1698175906
transform 1 0 25088 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_276
timestamp 1698175906
transform 1 0 32256 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_282
timestamp 1698175906
transform 1 0 32928 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_346
timestamp 1698175906
transform 1 0 40096 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_348
timestamp 1698175906
transform 1 0 40320 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_28
timestamp 1698175906
transform 1 0 4480 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_32
timestamp 1698175906
transform 1 0 4928 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698175906
transform 1 0 5152 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_37
timestamp 1698175906
transform 1 0 5488 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_101
timestamp 1698175906
transform 1 0 12656 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_107
timestamp 1698175906
transform 1 0 13328 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_111
timestamp 1698175906
transform 1 0 13776 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_117
timestamp 1698175906
transform 1 0 14448 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_167
timestamp 1698175906
transform 1 0 20048 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_173
timestamp 1698175906
transform 1 0 20720 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_186
timestamp 1698175906
transform 1 0 22176 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_191
timestamp 1698175906
transform 1 0 22736 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_199
timestamp 1698175906
transform 1 0 23632 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_201
timestamp 1698175906
transform 1 0 23856 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_204
timestamp 1698175906
transform 1 0 24192 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_236
timestamp 1698175906
transform 1 0 27776 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_244
timestamp 1698175906
transform 1 0 28672 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_247
timestamp 1698175906
transform 1 0 29008 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_311
timestamp 1698175906
transform 1 0 36176 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_317
timestamp 1698175906
transform 1 0 36848 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_2
timestamp 1698175906
transform 1 0 1568 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_66
timestamp 1698175906
transform 1 0 8736 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_72
timestamp 1698175906
transform 1 0 9408 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_88
timestamp 1698175906
transform 1 0 11200 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_92
timestamp 1698175906
transform 1 0 11648 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_94
timestamp 1698175906
transform 1 0 11872 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_124
timestamp 1698175906
transform 1 0 15232 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_128
timestamp 1698175906
transform 1 0 15680 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_136
timestamp 1698175906
transform 1 0 16576 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_171
timestamp 1698175906
transform 1 0 20496 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_208
timestamp 1698175906
transform 1 0 24640 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_212
timestamp 1698175906
transform 1 0 25088 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_276
timestamp 1698175906
transform 1 0 32256 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_282
timestamp 1698175906
transform 1 0 32928 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_346
timestamp 1698175906
transform 1 0 40096 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_348
timestamp 1698175906
transform 1 0 40320 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_2
timestamp 1698175906
transform 1 0 1568 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698175906
transform 1 0 5152 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_37
timestamp 1698175906
transform 1 0 5488 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_101
timestamp 1698175906
transform 1 0 12656 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_107
timestamp 1698175906
transform 1 0 13328 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_139
timestamp 1698175906
transform 1 0 16912 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_152
timestamp 1698175906
transform 1 0 18368 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_159
timestamp 1698175906
transform 1 0 19152 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_165
timestamp 1698175906
transform 1 0 19824 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_173
timestamp 1698175906
transform 1 0 20720 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_177
timestamp 1698175906
transform 1 0 21168 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_241
timestamp 1698175906
transform 1 0 28336 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_247
timestamp 1698175906
transform 1 0 29008 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_311
timestamp 1698175906
transform 1 0 36176 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_317
timestamp 1698175906
transform 1 0 36848 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_2
timestamp 1698175906
transform 1 0 1568 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_66
timestamp 1698175906
transform 1 0 8736 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_72
timestamp 1698175906
transform 1 0 9408 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_136
timestamp 1698175906
transform 1 0 16576 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_142
timestamp 1698175906
transform 1 0 17248 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_206
timestamp 1698175906
transform 1 0 24416 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_212
timestamp 1698175906
transform 1 0 25088 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_276
timestamp 1698175906
transform 1 0 32256 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_282
timestamp 1698175906
transform 1 0 32928 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_346
timestamp 1698175906
transform 1 0 40096 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_348
timestamp 1698175906
transform 1 0 40320 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698175906
transform 1 0 1568 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698175906
transform 1 0 5152 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_37
timestamp 1698175906
transform 1 0 5488 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_101
timestamp 1698175906
transform 1 0 12656 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_107
timestamp 1698175906
transform 1 0 13328 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_171
timestamp 1698175906
transform 1 0 20496 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_177
timestamp 1698175906
transform 1 0 21168 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_241
timestamp 1698175906
transform 1 0 28336 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_247
timestamp 1698175906
transform 1 0 29008 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_311
timestamp 1698175906
transform 1 0 36176 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_317
timestamp 1698175906
transform 1 0 36848 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2
timestamp 1698175906
transform 1 0 1568 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_66
timestamp 1698175906
transform 1 0 8736 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_72
timestamp 1698175906
transform 1 0 9408 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_136
timestamp 1698175906
transform 1 0 16576 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_142
timestamp 1698175906
transform 1 0 17248 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_206
timestamp 1698175906
transform 1 0 24416 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_212
timestamp 1698175906
transform 1 0 25088 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_276
timestamp 1698175906
transform 1 0 32256 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_282
timestamp 1698175906
transform 1 0 32928 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_346
timestamp 1698175906
transform 1 0 40096 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_348
timestamp 1698175906
transform 1 0 40320 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_2
timestamp 1698175906
transform 1 0 1568 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698175906
transform 1 0 5152 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_37
timestamp 1698175906
transform 1 0 5488 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_101
timestamp 1698175906
transform 1 0 12656 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_107
timestamp 1698175906
transform 1 0 13328 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_171
timestamp 1698175906
transform 1 0 20496 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_177
timestamp 1698175906
transform 1 0 21168 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_241
timestamp 1698175906
transform 1 0 28336 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_247
timestamp 1698175906
transform 1 0 29008 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_311
timestamp 1698175906
transform 1 0 36176 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_317
timestamp 1698175906
transform 1 0 36848 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2
timestamp 1698175906
transform 1 0 1568 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_66
timestamp 1698175906
transform 1 0 8736 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_72
timestamp 1698175906
transform 1 0 9408 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_136
timestamp 1698175906
transform 1 0 16576 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_142
timestamp 1698175906
transform 1 0 17248 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_206
timestamp 1698175906
transform 1 0 24416 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_212
timestamp 1698175906
transform 1 0 25088 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_276
timestamp 1698175906
transform 1 0 32256 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_282
timestamp 1698175906
transform 1 0 32928 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_346
timestamp 1698175906
transform 1 0 40096 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_348
timestamp 1698175906
transform 1 0 40320 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698175906
transform 1 0 1568 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698175906
transform 1 0 5152 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_37
timestamp 1698175906
transform 1 0 5488 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_101
timestamp 1698175906
transform 1 0 12656 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_107
timestamp 1698175906
transform 1 0 13328 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_171
timestamp 1698175906
transform 1 0 20496 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_177
timestamp 1698175906
transform 1 0 21168 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_241
timestamp 1698175906
transform 1 0 28336 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_247
timestamp 1698175906
transform 1 0 29008 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_311
timestamp 1698175906
transform 1 0 36176 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_317
timestamp 1698175906
transform 1 0 36848 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_2
timestamp 1698175906
transform 1 0 1568 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_66
timestamp 1698175906
transform 1 0 8736 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_72
timestamp 1698175906
transform 1 0 9408 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_136
timestamp 1698175906
transform 1 0 16576 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_142
timestamp 1698175906
transform 1 0 17248 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_206
timestamp 1698175906
transform 1 0 24416 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_212
timestamp 1698175906
transform 1 0 25088 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_276
timestamp 1698175906
transform 1 0 32256 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_282
timestamp 1698175906
transform 1 0 32928 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_346
timestamp 1698175906
transform 1 0 40096 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_348
timestamp 1698175906
transform 1 0 40320 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698175906
transform 1 0 1568 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698175906
transform 1 0 5152 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_37
timestamp 1698175906
transform 1 0 5488 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_101
timestamp 1698175906
transform 1 0 12656 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_107
timestamp 1698175906
transform 1 0 13328 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_171
timestamp 1698175906
transform 1 0 20496 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_177
timestamp 1698175906
transform 1 0 21168 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_241
timestamp 1698175906
transform 1 0 28336 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_247
timestamp 1698175906
transform 1 0 29008 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_311
timestamp 1698175906
transform 1 0 36176 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_317
timestamp 1698175906
transform 1 0 36848 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2
timestamp 1698175906
transform 1 0 1568 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1698175906
transform 1 0 8736 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_72
timestamp 1698175906
transform 1 0 9408 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_136
timestamp 1698175906
transform 1 0 16576 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_142
timestamp 1698175906
transform 1 0 17248 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_206
timestamp 1698175906
transform 1 0 24416 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_212
timestamp 1698175906
transform 1 0 25088 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_276
timestamp 1698175906
transform 1 0 32256 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_282
timestamp 1698175906
transform 1 0 32928 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_346
timestamp 1698175906
transform 1 0 40096 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_348
timestamp 1698175906
transform 1 0 40320 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_6
timestamp 1698175906
transform 1 0 2016 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_22
timestamp 1698175906
transform 1 0 3808 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_30
timestamp 1698175906
transform 1 0 4704 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698175906
transform 1 0 5152 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_37
timestamp 1698175906
transform 1 0 5488 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_101
timestamp 1698175906
transform 1 0 12656 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_107
timestamp 1698175906
transform 1 0 13328 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_139
timestamp 1698175906
transform 1 0 16912 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_143
timestamp 1698175906
transform 1 0 17360 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_171
timestamp 1698175906
transform 1 0 20496 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_177
timestamp 1698175906
transform 1 0 21168 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_193
timestamp 1698175906
transform 1 0 22960 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_197
timestamp 1698175906
transform 1 0 23408 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_225
timestamp 1698175906
transform 1 0 26544 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_241
timestamp 1698175906
transform 1 0 28336 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_247
timestamp 1698175906
transform 1 0 29008 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_311
timestamp 1698175906
transform 1 0 36176 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_317
timestamp 1698175906
transform 1 0 36848 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_2
timestamp 1698175906
transform 1 0 1568 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_66
timestamp 1698175906
transform 1 0 8736 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_72
timestamp 1698175906
transform 1 0 9408 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_136
timestamp 1698175906
transform 1 0 16576 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_142
timestamp 1698175906
transform 1 0 17248 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_150
timestamp 1698175906
transform 1 0 18144 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_155
timestamp 1698175906
transform 1 0 18704 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_189
timestamp 1698175906
transform 1 0 22512 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_205
timestamp 1698175906
transform 1 0 24304 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_209
timestamp 1698175906
transform 1 0 24752 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_212
timestamp 1698175906
transform 1 0 25088 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_276
timestamp 1698175906
transform 1 0 32256 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_282
timestamp 1698175906
transform 1 0 32928 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_346
timestamp 1698175906
transform 1 0 40096 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_348
timestamp 1698175906
transform 1 0 40320 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_2
timestamp 1698175906
transform 1 0 1568 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_36
timestamp 1698175906
transform 1 0 5376 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_70
timestamp 1698175906
transform 1 0 9184 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_104
timestamp 1698175906
transform 1 0 12992 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_138
timestamp 1698175906
transform 1 0 16800 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_142
timestamp 1698175906
transform 1 0 17248 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_172
timestamp 1698175906
transform 1 0 20608 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_176
timestamp 1698175906
transform 1 0 21056 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_236
timestamp 1698175906
transform 1 0 27776 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_240
timestamp 1698175906
transform 1 0 28224 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_274
timestamp 1698175906
transform 1 0 32032 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_308
timestamp 1698175906
transform 1 0 35840 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_342
timestamp 1698175906
transform 1 0 39648 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_346
timestamp 1698175906
transform 1 0 40096 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_348
timestamp 1698175906
transform 1 0 40320 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita4_23 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 17248 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita4_24
timestamp 1698175906
transform -1 0 27776 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita4_25
timestamp 1698175906
transform -1 0 2016 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita4_26
timestamp 1698175906
transform -1 0 18704 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 20944 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output2
timestamp 1698175906
transform 1 0 37520 0 1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output3
timestamp 1698175906
transform 1 0 21280 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output4
timestamp 1698175906
transform 1 0 21280 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output5
timestamp 1698175906
transform 1 0 23632 0 1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output6
timestamp 1698175906
transform 1 0 24416 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output7
timestamp 1698175906
transform -1 0 4480 0 -1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output8
timestamp 1698175906
transform -1 0 4480 0 1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output9
timestamp 1698175906
transform 1 0 37520 0 -1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output10
timestamp 1698175906
transform 1 0 37520 0 1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output11
timestamp 1698175906
transform -1 0 4480 0 -1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output12
timestamp 1698175906
transform 1 0 37520 0 -1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output13
timestamp 1698175906
transform -1 0 4480 0 1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output14
timestamp 1698175906
transform 1 0 37520 0 -1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output15
timestamp 1698175906
transform 1 0 37520 0 -1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output16
timestamp 1698175906
transform -1 0 4480 0 1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output17
timestamp 1698175906
transform 1 0 17584 0 1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output18
timestamp 1698175906
transform 1 0 24416 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output19
timestamp 1698175906
transform 1 0 19600 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output20
timestamp 1698175906
transform -1 0 20384 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output21
timestamp 1698175906
transform 1 0 25648 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output22
timestamp 1698175906
transform 1 0 37520 0 -1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_45 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698175906
transform -1 0 40656 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_46
timestamp 1698175906
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698175906
transform -1 0 40656 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_47
timestamp 1698175906
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698175906
transform -1 0 40656 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_48
timestamp 1698175906
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698175906
transform -1 0 40656 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_49
timestamp 1698175906
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698175906
transform -1 0 40656 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_50
timestamp 1698175906
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698175906
transform -1 0 40656 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_51
timestamp 1698175906
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698175906
transform -1 0 40656 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_52
timestamp 1698175906
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698175906
transform -1 0 40656 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_53
timestamp 1698175906
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698175906
transform -1 0 40656 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_54
timestamp 1698175906
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698175906
transform -1 0 40656 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_55
timestamp 1698175906
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698175906
transform -1 0 40656 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_56
timestamp 1698175906
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698175906
transform -1 0 40656 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_57
timestamp 1698175906
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698175906
transform -1 0 40656 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_58
timestamp 1698175906
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698175906
transform -1 0 40656 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_59
timestamp 1698175906
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698175906
transform -1 0 40656 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_60
timestamp 1698175906
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698175906
transform -1 0 40656 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_61
timestamp 1698175906
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698175906
transform -1 0 40656 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_62
timestamp 1698175906
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698175906
transform -1 0 40656 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_63
timestamp 1698175906
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698175906
transform -1 0 40656 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_64
timestamp 1698175906
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698175906
transform -1 0 40656 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_65
timestamp 1698175906
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698175906
transform -1 0 40656 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_66
timestamp 1698175906
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698175906
transform -1 0 40656 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_67
timestamp 1698175906
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698175906
transform -1 0 40656 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_68
timestamp 1698175906
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698175906
transform -1 0 40656 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_69
timestamp 1698175906
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698175906
transform -1 0 40656 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_70
timestamp 1698175906
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698175906
transform -1 0 40656 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_71
timestamp 1698175906
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698175906
transform -1 0 40656 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_72
timestamp 1698175906
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698175906
transform -1 0 40656 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_73
timestamp 1698175906
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698175906
transform -1 0 40656 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_74
timestamp 1698175906
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698175906
transform -1 0 40656 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_75
timestamp 1698175906
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698175906
transform -1 0 40656 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_76
timestamp 1698175906
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698175906
transform -1 0 40656 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_77
timestamp 1698175906
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698175906
transform -1 0 40656 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_78
timestamp 1698175906
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698175906
transform -1 0 40656 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_79
timestamp 1698175906
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698175906
transform -1 0 40656 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_80
timestamp 1698175906
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698175906
transform -1 0 40656 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_81
timestamp 1698175906
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698175906
transform -1 0 40656 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_82
timestamp 1698175906
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698175906
transform -1 0 40656 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_83
timestamp 1698175906
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698175906
transform -1 0 40656 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_84
timestamp 1698175906
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698175906
transform -1 0 40656 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_85
timestamp 1698175906
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698175906
transform -1 0 40656 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_86
timestamp 1698175906
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698175906
transform -1 0 40656 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_87
timestamp 1698175906
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698175906
transform -1 0 40656 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_88
timestamp 1698175906
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698175906
transform -1 0 40656 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_89
timestamp 1698175906
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698175906
transform -1 0 40656 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_90 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_91
timestamp 1698175906
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_92
timestamp 1698175906
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_93
timestamp 1698175906
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_94
timestamp 1698175906
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_95
timestamp 1698175906
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_96
timestamp 1698175906
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_97
timestamp 1698175906
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_98
timestamp 1698175906
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_99
timestamp 1698175906
transform 1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_100
timestamp 1698175906
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_101
timestamp 1698175906
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_102
timestamp 1698175906
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_103
timestamp 1698175906
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_104
timestamp 1698175906
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_105
timestamp 1698175906
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_106
timestamp 1698175906
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_107
timestamp 1698175906
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_108
timestamp 1698175906
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_109
timestamp 1698175906
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_110
timestamp 1698175906
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_111
timestamp 1698175906
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_112
timestamp 1698175906
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_113
timestamp 1698175906
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_114
timestamp 1698175906
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_115
timestamp 1698175906
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_116
timestamp 1698175906
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_117
timestamp 1698175906
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_118
timestamp 1698175906
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_119
timestamp 1698175906
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_120
timestamp 1698175906
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_121
timestamp 1698175906
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_122
timestamp 1698175906
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_123
timestamp 1698175906
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_124
timestamp 1698175906
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_125
timestamp 1698175906
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_126
timestamp 1698175906
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_127
timestamp 1698175906
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_128
timestamp 1698175906
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_129
timestamp 1698175906
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_130
timestamp 1698175906
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_131
timestamp 1698175906
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_132
timestamp 1698175906
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_133
timestamp 1698175906
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_134
timestamp 1698175906
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_135
timestamp 1698175906
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_136
timestamp 1698175906
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_137
timestamp 1698175906
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_138
timestamp 1698175906
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_139
timestamp 1698175906
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_140
timestamp 1698175906
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_141
timestamp 1698175906
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_142
timestamp 1698175906
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_143
timestamp 1698175906
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_144
timestamp 1698175906
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_145
timestamp 1698175906
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_146
timestamp 1698175906
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_147
timestamp 1698175906
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_148
timestamp 1698175906
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_149
timestamp 1698175906
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_150
timestamp 1698175906
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_151
timestamp 1698175906
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_152
timestamp 1698175906
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_153
timestamp 1698175906
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_154
timestamp 1698175906
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_155
timestamp 1698175906
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_156
timestamp 1698175906
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_157
timestamp 1698175906
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_158
timestamp 1698175906
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_159
timestamp 1698175906
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_160
timestamp 1698175906
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_161
timestamp 1698175906
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_162
timestamp 1698175906
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_163
timestamp 1698175906
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_164
timestamp 1698175906
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_165
timestamp 1698175906
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_166
timestamp 1698175906
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_167
timestamp 1698175906
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_168
timestamp 1698175906
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_169
timestamp 1698175906
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_170
timestamp 1698175906
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_171
timestamp 1698175906
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_172
timestamp 1698175906
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_173
timestamp 1698175906
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_174
timestamp 1698175906
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_175
timestamp 1698175906
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_176
timestamp 1698175906
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_177
timestamp 1698175906
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_178
timestamp 1698175906
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_179
timestamp 1698175906
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_180
timestamp 1698175906
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_181
timestamp 1698175906
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_182
timestamp 1698175906
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_183
timestamp 1698175906
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_184
timestamp 1698175906
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_185
timestamp 1698175906
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_186
timestamp 1698175906
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_187
timestamp 1698175906
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_188
timestamp 1698175906
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_189
timestamp 1698175906
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_190
timestamp 1698175906
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_191
timestamp 1698175906
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_192
timestamp 1698175906
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_193
timestamp 1698175906
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_194
timestamp 1698175906
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_195
timestamp 1698175906
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_196
timestamp 1698175906
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_197
timestamp 1698175906
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_198
timestamp 1698175906
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_199
timestamp 1698175906
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_200
timestamp 1698175906
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_201
timestamp 1698175906
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_202
timestamp 1698175906
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_203
timestamp 1698175906
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_204
timestamp 1698175906
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_205
timestamp 1698175906
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_206
timestamp 1698175906
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_207
timestamp 1698175906
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_208
timestamp 1698175906
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_209
timestamp 1698175906
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_210
timestamp 1698175906
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_211
timestamp 1698175906
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_212
timestamp 1698175906
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_213
timestamp 1698175906
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_214
timestamp 1698175906
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_215
timestamp 1698175906
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_216
timestamp 1698175906
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_217
timestamp 1698175906
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_218
timestamp 1698175906
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_219
timestamp 1698175906
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_220
timestamp 1698175906
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_221
timestamp 1698175906
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_222
timestamp 1698175906
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_223
timestamp 1698175906
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_224
timestamp 1698175906
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_225
timestamp 1698175906
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_226
timestamp 1698175906
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_227
timestamp 1698175906
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_228
timestamp 1698175906
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_229
timestamp 1698175906
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_230
timestamp 1698175906
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_231
timestamp 1698175906
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_232
timestamp 1698175906
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_233
timestamp 1698175906
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_234
timestamp 1698175906
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_235
timestamp 1698175906
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_236
timestamp 1698175906
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_237
timestamp 1698175906
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_238
timestamp 1698175906
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_239
timestamp 1698175906
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_240
timestamp 1698175906
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_241
timestamp 1698175906
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_242
timestamp 1698175906
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_243
timestamp 1698175906
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_244
timestamp 1698175906
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_245
timestamp 1698175906
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_246
timestamp 1698175906
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_247
timestamp 1698175906
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_248
timestamp 1698175906
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_249
timestamp 1698175906
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_250
timestamp 1698175906
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_251
timestamp 1698175906
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_252
timestamp 1698175906
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_253
timestamp 1698175906
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_254
timestamp 1698175906
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_255
timestamp 1698175906
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_256
timestamp 1698175906
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_257
timestamp 1698175906
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_258
timestamp 1698175906
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_259
timestamp 1698175906
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_260
timestamp 1698175906
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_261
timestamp 1698175906
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_262
timestamp 1698175906
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_263
timestamp 1698175906
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_264
timestamp 1698175906
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_265
timestamp 1698175906
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_266
timestamp 1698175906
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_267
timestamp 1698175906
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_268
timestamp 1698175906
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_269
timestamp 1698175906
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_270
timestamp 1698175906
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_271
timestamp 1698175906
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_272
timestamp 1698175906
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_273
timestamp 1698175906
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_274
timestamp 1698175906
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_275
timestamp 1698175906
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_276
timestamp 1698175906
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_277
timestamp 1698175906
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_278
timestamp 1698175906
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_279
timestamp 1698175906
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_280
timestamp 1698175906
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_281
timestamp 1698175906
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_282
timestamp 1698175906
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_283
timestamp 1698175906
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_284
timestamp 1698175906
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_285
timestamp 1698175906
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_286
timestamp 1698175906
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_287
timestamp 1698175906
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_288
timestamp 1698175906
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_289
timestamp 1698175906
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_290
timestamp 1698175906
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_291
timestamp 1698175906
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_292
timestamp 1698175906
transform 1 0 32704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_293
timestamp 1698175906
transform 1 0 5152 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_294
timestamp 1698175906
transform 1 0 8960 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_295
timestamp 1698175906
transform 1 0 12768 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_296
timestamp 1698175906
transform 1 0 16576 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_297
timestamp 1698175906
transform 1 0 20384 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_298
timestamp 1698175906
transform 1 0 24192 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_299
timestamp 1698175906
transform 1 0 28000 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_300
timestamp 1698175906
transform 1 0 31808 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_301
timestamp 1698175906
transform 1 0 35616 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_302
timestamp 1698175906
transform 1 0 39424 0 1 37632
box -86 -86 310 870
<< labels >>
flabel metal3 s 0 27552 800 27664 0 FreeSans 448 0 0 0 clk
port 0 nsew signal input
flabel metal2 s 16128 0 16240 800 0 FreeSans 448 90 0 0 segm[0]
port 1 nsew signal tristate
flabel metal2 s 20832 0 20944 800 0 FreeSans 448 90 0 0 segm[10]
port 2 nsew signal tristate
flabel metal3 s 41200 20160 42000 20272 0 FreeSans 448 0 0 0 segm[11]
port 3 nsew signal tristate
flabel metal2 s 22176 41200 22288 42000 0 FreeSans 448 90 0 0 segm[12]
port 4 nsew signal tristate
flabel metal2 s 21504 0 21616 800 0 FreeSans 448 90 0 0 segm[13]
port 5 nsew signal tristate
flabel metal2 s 23520 41200 23632 42000 0 FreeSans 448 90 0 0 segm[1]
port 6 nsew signal tristate
flabel metal2 s 26208 41200 26320 42000 0 FreeSans 448 90 0 0 segm[2]
port 7 nsew signal tristate
flabel metal3 s 0 36288 800 36400 0 FreeSans 448 0 0 0 segm[3]
port 8 nsew signal tristate
flabel metal2 s 22848 41200 22960 42000 0 FreeSans 448 90 0 0 segm[4]
port 9 nsew signal tristate
flabel metal2 s 18144 41200 18256 42000 0 FreeSans 448 90 0 0 segm[5]
port 10 nsew signal tristate
flabel metal3 s 0 24192 800 24304 0 FreeSans 448 0 0 0 segm[6]
port 11 nsew signal tristate
flabel metal3 s 0 23520 800 23632 0 FreeSans 448 0 0 0 segm[7]
port 12 nsew signal tristate
flabel metal3 s 41200 24192 42000 24304 0 FreeSans 448 0 0 0 segm[8]
port 13 nsew signal tristate
flabel metal3 s 41200 23520 42000 23632 0 FreeSans 448 0 0 0 segm[9]
port 14 nsew signal tristate
flabel metal3 s 0 16128 800 16240 0 FreeSans 448 0 0 0 sel[0]
port 15 nsew signal tristate
flabel metal3 s 41200 22848 42000 22960 0 FreeSans 448 0 0 0 sel[10]
port 16 nsew signal tristate
flabel metal3 s 0 24864 800 24976 0 FreeSans 448 0 0 0 sel[11]
port 17 nsew signal tristate
flabel metal3 s 41200 16128 42000 16240 0 FreeSans 448 0 0 0 sel[1]
port 18 nsew signal tristate
flabel metal3 s 41200 18144 42000 18256 0 FreeSans 448 0 0 0 sel[2]
port 19 nsew signal tristate
flabel metal3 s 0 26880 800 26992 0 FreeSans 448 0 0 0 sel[3]
port 20 nsew signal tristate
flabel metal2 s 17472 41200 17584 42000 0 FreeSans 448 90 0 0 sel[4]
port 21 nsew signal tristate
flabel metal2 s 24192 0 24304 800 0 FreeSans 448 90 0 0 sel[5]
port 22 nsew signal tristate
flabel metal2 s 19488 41200 19600 42000 0 FreeSans 448 90 0 0 sel[6]
port 23 nsew signal tristate
flabel metal2 s 18816 41200 18928 42000 0 FreeSans 448 90 0 0 sel[7]
port 24 nsew signal tristate
flabel metal2 s 25536 0 25648 800 0 FreeSans 448 90 0 0 sel[8]
port 25 nsew signal tristate
flabel metal3 s 41200 20832 42000 20944 0 FreeSans 448 0 0 0 sel[9]
port 26 nsew signal tristate
flabel metal4 s 4448 3076 4768 38476 0 FreeSans 1280 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 35168 3076 35488 38476 0 FreeSans 1280 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 19808 3076 20128 38476 0 FreeSans 1280 90 0 0 vss
port 28 nsew ground bidirectional
rlabel metal1 21000 38416 21000 38416 0 vdd
rlabel metal1 21000 37632 21000 37632 0 vss
rlabel metal2 27608 17248 27608 17248 0 _000_
rlabel metal2 26488 16296 26488 16296 0 _001_
rlabel metal2 14392 15624 14392 15624 0 _002_
rlabel metal2 25144 22792 25144 22792 0 _003_
rlabel metal2 27384 20804 27384 20804 0 _004_
rlabel metal2 18704 13048 18704 13048 0 _005_
rlabel metal2 20552 14056 20552 14056 0 _006_
rlabel metal2 27160 22736 27160 22736 0 _007_
rlabel metal2 12488 23968 12488 23968 0 _008_
rlabel metal2 21672 27440 21672 27440 0 _009_
rlabel metal2 12152 24640 12152 24640 0 _010_
rlabel metal2 16072 22792 16072 22792 0 _011_
rlabel metal2 23688 23576 23688 23576 0 _012_
rlabel metal2 21896 25872 21896 25872 0 _013_
rlabel metal2 24528 19320 24528 19320 0 _014_
rlabel metal2 24248 14868 24248 14868 0 _015_
rlabel metal3 19432 23184 19432 23184 0 _016_
rlabel metal2 18032 20664 18032 20664 0 _017_
rlabel metal2 13608 16912 13608 16912 0 _018_
rlabel metal2 15512 14784 15512 14784 0 _019_
rlabel metal2 17192 27776 17192 27776 0 _020_
rlabel metal2 19544 27384 19544 27384 0 _021_
rlabel metal3 23240 15176 23240 15176 0 _022_
rlabel metal2 15736 25928 15736 25928 0 _023_
rlabel metal2 14168 27496 14168 27496 0 _024_
rlabel metal2 25592 17360 25592 17360 0 _025_
rlabel metal2 21672 14896 21672 14896 0 _026_
rlabel metal2 16856 25424 16856 25424 0 _027_
rlabel metal2 16968 25536 16968 25536 0 _028_
rlabel metal2 14280 26208 14280 26208 0 _029_
rlabel metal2 27664 21112 27664 21112 0 _030_
rlabel metal2 26264 17528 26264 17528 0 _031_
rlabel metal2 22904 17248 22904 17248 0 _032_
rlabel metal3 27384 22232 27384 22232 0 _033_
rlabel metal2 29176 18144 29176 18144 0 _034_
rlabel metal2 25816 17360 25816 17360 0 _035_
rlabel metal2 19208 22120 19208 22120 0 _036_
rlabel metal3 17528 15288 17528 15288 0 _037_
rlabel metal2 15960 17024 15960 17024 0 _038_
rlabel metal3 18312 16632 18312 16632 0 _039_
rlabel metal3 15568 15960 15568 15960 0 _040_
rlabel metal2 26040 21952 26040 21952 0 _041_
rlabel metal3 25480 22344 25480 22344 0 _042_
rlabel metal2 23800 21616 23800 21616 0 _043_
rlabel metal3 28224 19432 28224 19432 0 _044_
rlabel metal2 27384 21784 27384 21784 0 _045_
rlabel metal2 27048 22064 27048 22064 0 _046_
rlabel metal2 20216 15288 20216 15288 0 _047_
rlabel metal2 19432 14952 19432 14952 0 _048_
rlabel metal2 19208 15680 19208 15680 0 _049_
rlabel metal2 20552 18984 20552 18984 0 _050_
rlabel metal2 21280 14616 21280 14616 0 _051_
rlabel metal3 28112 22120 28112 22120 0 _052_
rlabel metal2 12712 23744 12712 23744 0 _053_
rlabel metal2 21448 22848 21448 22848 0 _054_
rlabel metal3 22120 26936 22120 26936 0 _055_
rlabel metal3 22008 23800 22008 23800 0 _056_
rlabel metal3 21168 26824 21168 26824 0 _057_
rlabel metal2 13608 24136 13608 24136 0 _058_
rlabel metal2 15960 22904 15960 22904 0 _059_
rlabel metal2 23576 22792 23576 22792 0 _060_
rlabel metal2 24136 23800 24136 23800 0 _061_
rlabel metal3 22064 25256 22064 25256 0 _062_
rlabel metal2 20216 25088 20216 25088 0 _063_
rlabel metal2 20440 23520 20440 23520 0 _064_
rlabel metal2 20440 18648 20440 18648 0 _065_
rlabel metal2 22456 22120 22456 22120 0 _066_
rlabel metal2 19880 22232 19880 22232 0 _067_
rlabel metal2 22120 20776 22120 20776 0 _068_
rlabel metal3 23184 18984 23184 18984 0 _069_
rlabel metal2 17752 20832 17752 20832 0 _070_
rlabel metal3 18704 19880 18704 19880 0 _071_
rlabel metal2 22512 17640 22512 17640 0 _072_
rlabel metal2 20776 22008 20776 22008 0 _073_
rlabel metal2 20440 22792 20440 22792 0 _074_
rlabel metal2 24248 21728 24248 21728 0 _075_
rlabel metal3 24248 15512 24248 15512 0 _076_
rlabel metal2 19880 20832 19880 20832 0 _077_
rlabel metal2 19600 20776 19600 20776 0 _078_
rlabel metal2 23016 19824 23016 19824 0 _079_
rlabel metal3 17864 22232 17864 22232 0 _080_
rlabel metal2 20216 16184 20216 16184 0 _081_
rlabel metal2 24696 20720 24696 20720 0 _082_
rlabel metal2 21000 21952 21000 21952 0 _083_
rlabel metal2 24136 21896 24136 21896 0 _084_
rlabel metal3 18256 17416 18256 17416 0 _085_
rlabel metal2 24920 16464 24920 16464 0 _086_
rlabel metal2 21560 19712 21560 19712 0 _087_
rlabel metal2 16744 18816 16744 18816 0 _088_
rlabel metal2 13888 19208 13888 19208 0 _089_
rlabel metal2 14168 26992 14168 26992 0 _090_
rlabel metal2 17080 17920 17080 17920 0 _091_
rlabel metal3 15848 17528 15848 17528 0 _092_
rlabel metal2 20048 22232 20048 22232 0 _093_
rlabel metal2 17696 28056 17696 28056 0 _094_
rlabel metal2 20328 14280 20328 14280 0 _095_
rlabel metal2 17640 15904 17640 15904 0 _096_
rlabel metal3 17416 25256 17416 25256 0 _097_
rlabel metal2 19432 27720 19432 27720 0 _098_
rlabel metal2 18200 28560 18200 28560 0 _099_
rlabel metal2 22792 18928 22792 18928 0 _100_
rlabel metal3 17864 23912 17864 23912 0 _101_
rlabel metal2 19712 26936 19712 26936 0 _102_
rlabel metal2 19768 27048 19768 27048 0 _103_
rlabel metal2 23240 14784 23240 14784 0 _104_
rlabel metal2 24136 17976 24136 17976 0 _105_
rlabel metal3 2478 27608 2478 27608 0 clk
rlabel metal2 23240 20440 23240 20440 0 clknet_0_clk
rlabel metal2 21672 13272 21672 13272 0 clknet_1_0__leaf_clk
rlabel metal2 28168 22008 28168 22008 0 clknet_1_1__leaf_clk
rlabel metal2 14840 19600 14840 19600 0 dut4.count\[0\]
rlabel metal2 14392 19656 14392 19656 0 dut4.count\[1\]
rlabel metal3 16744 16744 16744 16744 0 dut4.count\[2\]
rlabel metal2 17584 14616 17584 14616 0 dut4.count\[3\]
rlabel metal2 21112 6356 21112 6356 0 net1
rlabel metal2 28168 23128 28168 23128 0 net10
rlabel metal2 12264 16016 12264 16016 0 net11
rlabel metal2 31416 22736 31416 22736 0 net12
rlabel metal2 10584 25032 10584 25032 0 net13
rlabel metal2 28616 16576 28616 16576 0 net14
rlabel metal2 29736 17136 29736 17136 0 net15
rlabel metal3 6356 27048 6356 27048 0 net16
rlabel metal2 16856 27496 16856 27496 0 net17
rlabel metal2 24584 5964 24584 5964 0 net18
rlabel metal2 20328 28112 20328 28112 0 net19
rlabel metal2 29288 19600 29288 19600 0 net2
rlabel metal2 19320 27720 19320 27720 0 net20
rlabel metal2 25816 6356 25816 6356 0 net21
rlabel metal2 37912 20832 37912 20832 0 net22
rlabel metal2 16184 2030 16184 2030 0 net23
rlabel metal3 26880 37912 26880 37912 0 net24
rlabel metal3 1246 36344 1246 36344 0 net25
rlabel metal2 18312 37464 18312 37464 0 net26
rlabel metal2 20832 31920 20832 31920 0 net3
rlabel metal2 21448 13944 21448 13944 0 net4
rlabel metal2 24136 32256 24136 32256 0 net5
rlabel metal3 24136 27832 24136 27832 0 net6
rlabel metal2 10024 24360 10024 24360 0 net7
rlabel metal2 13944 23464 13944 23464 0 net8
rlabel metal3 31920 24080 31920 24080 0 net9
rlabel metal2 20888 2422 20888 2422 0 segm[10]
rlabel metal2 40040 20552 40040 20552 0 segm[11]
rlabel metal2 22232 39746 22232 39746 0 segm[12]
rlabel metal2 21560 2198 21560 2198 0 segm[13]
rlabel metal2 23576 38962 23576 38962 0 segm[1]
rlabel metal2 22904 39746 22904 39746 0 segm[4]
rlabel metal3 1358 24248 1358 24248 0 segm[6]
rlabel metal3 1358 23576 1358 23576 0 segm[7]
rlabel metal2 40040 24360 40040 24360 0 segm[8]
rlabel metal2 40040 23800 40040 23800 0 segm[9]
rlabel metal3 1358 16184 1358 16184 0 sel[0]
rlabel metal3 40642 22904 40642 22904 0 sel[10]
rlabel metal3 1358 24920 1358 24920 0 sel[11]
rlabel metal2 40040 16408 40040 16408 0 sel[1]
rlabel metal3 40642 18200 40642 18200 0 sel[2]
rlabel metal3 1358 26936 1358 26936 0 sel[3]
rlabel metal2 17528 38962 17528 38962 0 sel[4]
rlabel metal2 24248 2198 24248 2198 0 sel[5]
rlabel metal2 20776 38024 20776 38024 0 sel[6]
rlabel metal2 18872 39690 18872 39690 0 sel[7]
rlabel metal2 25592 2086 25592 2086 0 sel[8]
rlabel metal2 39928 21168 39928 21168 0 sel[9]
<< properties >>
string FIXED_BBOX 0 0 42000 42000
<< end >>
