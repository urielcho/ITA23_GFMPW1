magic
tech gf180mcuD
magscale 1 5
timestamp 1699642920
<< metal1 >>
rect 672 19221 20328 19238
rect 672 19195 2239 19221
rect 2265 19195 2291 19221
rect 2317 19195 2343 19221
rect 2369 19195 17599 19221
rect 17625 19195 17651 19221
rect 17677 19195 17703 19221
rect 17729 19195 20328 19221
rect 672 19178 20328 19195
rect 11047 19137 11073 19143
rect 11047 19105 11073 19111
rect 12783 19137 12809 19143
rect 12783 19105 12809 19111
rect 9417 19055 9423 19081
rect 9449 19055 9455 19081
rect 9025 18999 9031 19025
rect 9057 18999 9063 19025
rect 10649 18999 10655 19025
rect 10681 18999 10687 19025
rect 12273 18999 12279 19025
rect 12305 18999 12311 19025
rect 672 18829 20328 18846
rect 672 18803 9919 18829
rect 9945 18803 9971 18829
rect 9997 18803 10023 18829
rect 10049 18803 20328 18829
rect 672 18786 20328 18803
rect 10711 18745 10737 18751
rect 10711 18713 10737 18719
rect 13399 18745 13425 18751
rect 13399 18713 13425 18719
rect 20119 18689 20145 18695
rect 20119 18657 20145 18663
rect 10369 18607 10375 18633
rect 10401 18607 10407 18633
rect 13001 18607 13007 18633
rect 13033 18607 13039 18633
rect 672 18437 20328 18454
rect 672 18411 2239 18437
rect 2265 18411 2291 18437
rect 2317 18411 2343 18437
rect 2369 18411 17599 18437
rect 17625 18411 17651 18437
rect 17677 18411 17703 18437
rect 17729 18411 20328 18437
rect 672 18394 20328 18411
rect 672 18045 20328 18062
rect 672 18019 9919 18045
rect 9945 18019 9971 18045
rect 9997 18019 10023 18045
rect 10049 18019 20328 18045
rect 672 18002 20328 18019
rect 672 17653 20328 17670
rect 672 17627 2239 17653
rect 2265 17627 2291 17653
rect 2317 17627 2343 17653
rect 2369 17627 17599 17653
rect 17625 17627 17651 17653
rect 17677 17627 17703 17653
rect 17729 17627 20328 17653
rect 672 17610 20328 17627
rect 20119 17345 20145 17351
rect 20119 17313 20145 17319
rect 672 17261 20328 17278
rect 672 17235 9919 17261
rect 9945 17235 9971 17261
rect 9997 17235 10023 17261
rect 10049 17235 20328 17261
rect 672 17218 20328 17235
rect 672 16869 20328 16886
rect 672 16843 2239 16869
rect 2265 16843 2291 16869
rect 2317 16843 2343 16869
rect 2369 16843 17599 16869
rect 17625 16843 17651 16869
rect 17677 16843 17703 16869
rect 17729 16843 20328 16869
rect 672 16826 20328 16843
rect 672 16477 20328 16494
rect 672 16451 9919 16477
rect 9945 16451 9971 16477
rect 9997 16451 10023 16477
rect 10049 16451 20328 16477
rect 672 16434 20328 16451
rect 672 16085 20328 16102
rect 672 16059 2239 16085
rect 2265 16059 2291 16085
rect 2317 16059 2343 16085
rect 2369 16059 17599 16085
rect 17625 16059 17651 16085
rect 17677 16059 17703 16085
rect 17729 16059 20328 16085
rect 672 16042 20328 16059
rect 672 15693 20328 15710
rect 672 15667 9919 15693
rect 9945 15667 9971 15693
rect 9997 15667 10023 15693
rect 10049 15667 20328 15693
rect 672 15650 20328 15667
rect 672 15301 20328 15318
rect 672 15275 2239 15301
rect 2265 15275 2291 15301
rect 2317 15275 2343 15301
rect 2369 15275 17599 15301
rect 17625 15275 17651 15301
rect 17677 15275 17703 15301
rect 17729 15275 20328 15301
rect 672 15258 20328 15275
rect 672 14909 20328 14926
rect 672 14883 9919 14909
rect 9945 14883 9971 14909
rect 9997 14883 10023 14909
rect 10049 14883 20328 14909
rect 672 14866 20328 14883
rect 672 14517 20328 14534
rect 672 14491 2239 14517
rect 2265 14491 2291 14517
rect 2317 14491 2343 14517
rect 2369 14491 17599 14517
rect 17625 14491 17651 14517
rect 17677 14491 17703 14517
rect 17729 14491 20328 14517
rect 672 14474 20328 14491
rect 672 14125 20328 14142
rect 672 14099 9919 14125
rect 9945 14099 9971 14125
rect 9997 14099 10023 14125
rect 10049 14099 20328 14125
rect 672 14082 20328 14099
rect 18937 13903 18943 13929
rect 18969 13903 18975 13929
rect 12951 13873 12977 13879
rect 19945 13847 19951 13873
rect 19977 13847 19983 13873
rect 12951 13841 12977 13847
rect 672 13733 20328 13750
rect 672 13707 2239 13733
rect 2265 13707 2291 13733
rect 2317 13707 2343 13733
rect 2369 13707 17599 13733
rect 17625 13707 17651 13733
rect 17677 13707 17703 13733
rect 17729 13707 20328 13733
rect 672 13690 20328 13707
rect 967 13593 993 13599
rect 20007 13593 20033 13599
rect 10369 13567 10375 13593
rect 10401 13567 10407 13593
rect 12777 13567 12783 13593
rect 12809 13567 12815 13593
rect 967 13561 993 13567
rect 20007 13561 20033 13567
rect 12895 13537 12921 13543
rect 2137 13511 2143 13537
rect 2169 13511 2175 13537
rect 8969 13511 8975 13537
rect 9001 13511 9007 13537
rect 10761 13511 10767 13537
rect 10793 13511 10799 13537
rect 11377 13511 11383 13537
rect 11409 13511 11415 13537
rect 12895 13505 12921 13511
rect 13343 13537 13369 13543
rect 18825 13511 18831 13537
rect 18857 13511 18863 13537
rect 13343 13505 13369 13511
rect 8751 13481 8777 13487
rect 11103 13481 11129 13487
rect 9305 13455 9311 13481
rect 9337 13455 9343 13481
rect 10649 13455 10655 13481
rect 10681 13455 10687 13481
rect 8751 13449 8777 13455
rect 11103 13449 11129 13455
rect 11159 13481 11185 13487
rect 13007 13481 13033 13487
rect 11713 13455 11719 13481
rect 11745 13455 11751 13481
rect 11159 13449 11185 13455
rect 13007 13449 13033 13455
rect 13063 13481 13089 13487
rect 13063 13449 13089 13455
rect 13399 13481 13425 13487
rect 13399 13449 13425 13455
rect 10991 13425 11017 13431
rect 10991 13393 11017 13399
rect 13511 13425 13537 13431
rect 13511 13393 13537 13399
rect 672 13341 20328 13358
rect 672 13315 9919 13341
rect 9945 13315 9971 13341
rect 9997 13315 10023 13341
rect 10049 13315 20328 13341
rect 672 13298 20328 13315
rect 9703 13257 9729 13263
rect 9703 13225 9729 13231
rect 9927 13257 9953 13263
rect 11831 13257 11857 13263
rect 10089 13231 10095 13257
rect 10121 13231 10127 13257
rect 9927 13225 9953 13231
rect 11831 13225 11857 13231
rect 9199 13201 9225 13207
rect 9199 13169 9225 13175
rect 11943 13201 11969 13207
rect 11943 13169 11969 13175
rect 11999 13201 12025 13207
rect 11999 13169 12025 13175
rect 12951 13201 12977 13207
rect 12951 13169 12977 13175
rect 13007 13201 13033 13207
rect 13007 13169 13033 13175
rect 14799 13201 14825 13207
rect 14961 13175 14967 13201
rect 14993 13175 14999 13201
rect 14799 13169 14825 13175
rect 9143 13145 9169 13151
rect 2137 13119 2143 13145
rect 2169 13119 2175 13145
rect 8017 13119 8023 13145
rect 8049 13119 8055 13145
rect 9143 13113 9169 13119
rect 9311 13145 9337 13151
rect 9311 13113 9337 13119
rect 9647 13145 9673 13151
rect 9647 13113 9673 13119
rect 9815 13145 9841 13151
rect 12839 13145 12865 13151
rect 10313 13119 10319 13145
rect 10345 13119 10351 13145
rect 13169 13119 13175 13145
rect 13201 13119 13207 13145
rect 18825 13119 18831 13145
rect 18857 13119 18863 13145
rect 9815 13113 9841 13119
rect 12839 13113 12865 13119
rect 8303 13089 8329 13095
rect 12223 13089 12249 13095
rect 6617 13063 6623 13089
rect 6649 13063 6655 13089
rect 7681 13063 7687 13089
rect 7713 13063 7719 13089
rect 10649 13063 10655 13089
rect 10681 13063 10687 13089
rect 11713 13063 11719 13089
rect 11745 13063 11751 13089
rect 8303 13057 8329 13063
rect 12223 13057 12249 13063
rect 12727 13089 12753 13095
rect 13561 13063 13567 13089
rect 13593 13063 13599 13089
rect 14625 13063 14631 13089
rect 14657 13063 14663 13089
rect 12727 13057 12753 13063
rect 967 13033 993 13039
rect 967 13001 993 13007
rect 20007 13033 20033 13039
rect 20007 13001 20033 13007
rect 672 12949 20328 12966
rect 672 12923 2239 12949
rect 2265 12923 2291 12949
rect 2317 12923 2343 12949
rect 2369 12923 17599 12949
rect 17625 12923 17651 12949
rect 17677 12923 17703 12949
rect 17729 12923 20328 12949
rect 672 12906 20328 12923
rect 10095 12865 10121 12871
rect 10095 12833 10121 12839
rect 7295 12809 7321 12815
rect 10375 12809 10401 12815
rect 7569 12783 7575 12809
rect 7601 12783 7607 12809
rect 9473 12783 9479 12809
rect 9505 12783 9511 12809
rect 13505 12783 13511 12809
rect 13537 12783 13543 12809
rect 7295 12777 7321 12783
rect 10375 12777 10401 12783
rect 7631 12753 7657 12759
rect 9815 12753 9841 12759
rect 8017 12727 8023 12753
rect 8049 12727 8055 12753
rect 7631 12721 7657 12727
rect 9815 12721 9841 12727
rect 10151 12753 10177 12759
rect 10151 12721 10177 12727
rect 10879 12753 10905 12759
rect 10879 12721 10905 12727
rect 11047 12753 11073 12759
rect 13623 12753 13649 12759
rect 12105 12727 12111 12753
rect 12137 12727 12143 12753
rect 11047 12721 11073 12727
rect 13623 12721 13649 12727
rect 13791 12753 13817 12759
rect 13791 12721 13817 12727
rect 6847 12697 6873 12703
rect 6847 12665 6873 12671
rect 7351 12697 7377 12703
rect 7351 12665 7377 12671
rect 7855 12697 7881 12703
rect 8409 12671 8415 12697
rect 8441 12671 8447 12697
rect 12441 12671 12447 12697
rect 12473 12671 12479 12697
rect 7855 12665 7881 12671
rect 6903 12641 6929 12647
rect 6903 12609 6929 12615
rect 7575 12641 7601 12647
rect 7575 12609 7601 12615
rect 7743 12641 7769 12647
rect 7743 12609 7769 12615
rect 9927 12641 9953 12647
rect 9927 12609 9953 12615
rect 10039 12641 10065 12647
rect 10039 12609 10065 12615
rect 10991 12641 11017 12647
rect 10991 12609 11017 12615
rect 13735 12641 13761 12647
rect 13735 12609 13761 12615
rect 14015 12641 14041 12647
rect 14015 12609 14041 12615
rect 672 12557 20328 12574
rect 672 12531 9919 12557
rect 9945 12531 9971 12557
rect 9997 12531 10023 12557
rect 10049 12531 20328 12557
rect 672 12514 20328 12531
rect 7631 12473 7657 12479
rect 7631 12441 7657 12447
rect 7743 12473 7769 12479
rect 7743 12441 7769 12447
rect 9031 12473 9057 12479
rect 12559 12473 12585 12479
rect 9417 12447 9423 12473
rect 9449 12447 9455 12473
rect 9031 12441 9057 12447
rect 12559 12441 12585 12447
rect 12671 12417 12697 12423
rect 7009 12391 7015 12417
rect 7041 12391 7047 12417
rect 12671 12385 12697 12391
rect 12727 12417 12753 12423
rect 12727 12385 12753 12391
rect 7687 12361 7713 12367
rect 7401 12335 7407 12361
rect 7433 12335 7439 12361
rect 7687 12329 7713 12335
rect 7799 12361 7825 12367
rect 8975 12361 9001 12367
rect 7905 12335 7911 12361
rect 7937 12335 7943 12361
rect 7799 12329 7825 12335
rect 8975 12329 9001 12335
rect 9087 12361 9113 12367
rect 9087 12329 9113 12335
rect 9311 12361 9337 12367
rect 9815 12361 9841 12367
rect 9529 12335 9535 12361
rect 9561 12335 9567 12361
rect 9311 12329 9337 12335
rect 9815 12329 9841 12335
rect 5945 12279 5951 12305
rect 5977 12279 5983 12305
rect 672 12165 20328 12182
rect 672 12139 2239 12165
rect 2265 12139 2291 12165
rect 2317 12139 2343 12165
rect 2369 12139 17599 12165
rect 17625 12139 17651 12165
rect 17677 12139 17703 12165
rect 17729 12139 20328 12165
rect 672 12122 20328 12139
rect 967 12025 993 12031
rect 967 11993 993 11999
rect 7687 12025 7713 12031
rect 7687 11993 7713 11999
rect 12391 12025 12417 12031
rect 12391 11993 12417 11999
rect 7463 11969 7489 11975
rect 2137 11943 2143 11969
rect 2169 11943 2175 11969
rect 7463 11937 7489 11943
rect 9759 11969 9785 11975
rect 9759 11937 9785 11943
rect 7407 11913 7433 11919
rect 7407 11881 7433 11887
rect 9591 11913 9617 11919
rect 9591 11881 9617 11887
rect 7295 11857 7321 11863
rect 7295 11825 7321 11831
rect 9647 11857 9673 11863
rect 9647 11825 9673 11831
rect 672 11773 20328 11790
rect 672 11747 9919 11773
rect 9945 11747 9971 11773
rect 9997 11747 10023 11773
rect 10049 11747 20328 11773
rect 672 11730 20328 11747
rect 7351 11689 7377 11695
rect 7351 11657 7377 11663
rect 8919 11689 8945 11695
rect 8919 11657 8945 11663
rect 10207 11689 10233 11695
rect 10207 11657 10233 11663
rect 10319 11689 10345 11695
rect 10319 11657 10345 11663
rect 14631 11689 14657 11695
rect 14631 11657 14657 11663
rect 8863 11633 8889 11639
rect 8863 11601 8889 11607
rect 12727 11633 12753 11639
rect 12727 11601 12753 11607
rect 7519 11577 7545 11583
rect 7121 11551 7127 11577
rect 7153 11551 7159 11577
rect 7519 11545 7545 11551
rect 7631 11577 7657 11583
rect 7631 11545 7657 11551
rect 7743 11577 7769 11583
rect 10151 11577 10177 11583
rect 9025 11551 9031 11577
rect 9057 11551 9063 11577
rect 7743 11545 7769 11551
rect 10151 11545 10177 11551
rect 11999 11577 12025 11583
rect 11999 11545 12025 11551
rect 12111 11577 12137 11583
rect 12783 11577 12809 11583
rect 12273 11551 12279 11577
rect 12305 11551 12311 11577
rect 13001 11551 13007 11577
rect 13033 11551 13039 11577
rect 18825 11551 18831 11577
rect 18857 11551 18863 11577
rect 12111 11545 12137 11551
rect 12783 11545 12809 11551
rect 7575 11521 7601 11527
rect 5665 11495 5671 11521
rect 5697 11495 5703 11521
rect 6729 11495 6735 11521
rect 6761 11495 6767 11521
rect 7575 11489 7601 11495
rect 9871 11521 9897 11527
rect 9871 11489 9897 11495
rect 12055 11521 12081 11527
rect 13337 11495 13343 11521
rect 13369 11495 13375 11521
rect 14401 11495 14407 11521
rect 14433 11495 14439 11521
rect 12055 11489 12081 11495
rect 9927 11465 9953 11471
rect 9927 11433 9953 11439
rect 12727 11465 12753 11471
rect 12727 11433 12753 11439
rect 20007 11465 20033 11471
rect 20007 11433 20033 11439
rect 672 11381 20328 11398
rect 672 11355 2239 11381
rect 2265 11355 2291 11381
rect 2317 11355 2343 11381
rect 2369 11355 17599 11381
rect 17625 11355 17651 11381
rect 17677 11355 17703 11381
rect 17729 11355 20328 11381
rect 672 11338 20328 11355
rect 10151 11297 10177 11303
rect 10151 11265 10177 11271
rect 967 11241 993 11247
rect 13343 11241 13369 11247
rect 9025 11215 9031 11241
rect 9057 11215 9063 11241
rect 12217 11215 12223 11241
rect 12249 11215 12255 11241
rect 967 11209 993 11215
rect 13343 11209 13369 11215
rect 20007 11241 20033 11247
rect 20007 11209 20033 11215
rect 7071 11185 7097 11191
rect 2137 11159 2143 11185
rect 2169 11159 2175 11185
rect 7071 11153 7097 11159
rect 7295 11185 7321 11191
rect 7295 11153 7321 11159
rect 7631 11185 7657 11191
rect 12671 11185 12697 11191
rect 13231 11185 13257 11191
rect 7961 11159 7967 11185
rect 7993 11159 7999 11185
rect 8633 11159 8639 11185
rect 8665 11159 8671 11185
rect 8857 11159 8863 11185
rect 8889 11159 8895 11185
rect 9921 11159 9927 11185
rect 9953 11159 9959 11185
rect 10817 11159 10823 11185
rect 10849 11159 10855 11185
rect 12553 11159 12559 11185
rect 12585 11159 12591 11185
rect 12889 11159 12895 11185
rect 12921 11159 12927 11185
rect 7631 11153 7657 11159
rect 12671 11153 12697 11159
rect 13231 11153 13257 11159
rect 13791 11185 13817 11191
rect 18825 11159 18831 11185
rect 18857 11159 18863 11185
rect 13791 11153 13817 11159
rect 7799 11129 7825 11135
rect 13511 11129 13537 11135
rect 8689 11103 8695 11129
rect 8721 11103 8727 11129
rect 8969 11103 8975 11129
rect 9001 11103 9007 11129
rect 9249 11103 9255 11129
rect 9281 11103 9287 11129
rect 9809 11103 9815 11129
rect 9841 11103 9847 11129
rect 11153 11103 11159 11129
rect 11185 11103 11191 11129
rect 7799 11097 7825 11103
rect 13511 11097 13537 11103
rect 13623 11129 13649 11135
rect 13623 11097 13649 11103
rect 7351 11073 7377 11079
rect 7351 11041 7377 11047
rect 7407 11073 7433 11079
rect 7407 11041 7433 11047
rect 7743 11073 7769 11079
rect 7743 11041 7769 11047
rect 9423 11073 9449 11079
rect 9423 11041 9449 11047
rect 10319 11073 10345 11079
rect 10319 11041 10345 11047
rect 12727 11073 12753 11079
rect 12727 11041 12753 11047
rect 12783 11073 12809 11079
rect 13679 11073 13705 11079
rect 13057 11047 13063 11073
rect 13089 11047 13095 11073
rect 12783 11041 12809 11047
rect 13679 11041 13705 11047
rect 672 10989 20328 11006
rect 672 10963 9919 10989
rect 9945 10963 9971 10989
rect 9997 10963 10023 10989
rect 10049 10963 20328 10989
rect 672 10946 20328 10963
rect 8751 10905 8777 10911
rect 11159 10905 11185 10911
rect 8241 10879 8247 10905
rect 8273 10879 8279 10905
rect 10033 10879 10039 10905
rect 10065 10879 10071 10905
rect 8751 10873 8777 10879
rect 11159 10873 11185 10879
rect 11495 10905 11521 10911
rect 11495 10873 11521 10879
rect 11887 10905 11913 10911
rect 11887 10873 11913 10879
rect 11999 10905 12025 10911
rect 11999 10873 12025 10879
rect 12167 10905 12193 10911
rect 12167 10873 12193 10879
rect 12671 10905 12697 10911
rect 12671 10873 12697 10879
rect 7463 10849 7489 10855
rect 6785 10823 6791 10849
rect 6817 10823 6823 10849
rect 7463 10817 7489 10823
rect 7967 10849 7993 10855
rect 7967 10817 7993 10823
rect 8023 10849 8049 10855
rect 10319 10849 10345 10855
rect 9697 10823 9703 10849
rect 9729 10823 9735 10849
rect 9921 10823 9927 10849
rect 9953 10823 9959 10849
rect 8023 10817 8049 10823
rect 10319 10817 10345 10823
rect 10599 10849 10625 10855
rect 10599 10817 10625 10823
rect 11047 10849 11073 10855
rect 11047 10817 11073 10823
rect 11775 10849 11801 10855
rect 11775 10817 11801 10823
rect 12727 10849 12753 10855
rect 12727 10817 12753 10823
rect 12783 10849 12809 10855
rect 12889 10823 12895 10849
rect 12921 10823 12927 10849
rect 13673 10823 13679 10849
rect 13705 10823 13711 10849
rect 12783 10817 12809 10823
rect 7743 10793 7769 10799
rect 10263 10793 10289 10799
rect 7121 10767 7127 10793
rect 7153 10767 7159 10793
rect 7569 10767 7575 10793
rect 7601 10767 7607 10793
rect 8353 10767 8359 10793
rect 8385 10767 8391 10793
rect 8801 10767 8807 10793
rect 8833 10767 8839 10793
rect 9529 10767 9535 10793
rect 9561 10767 9567 10793
rect 7743 10761 7769 10767
rect 10263 10761 10289 10767
rect 10543 10793 10569 10799
rect 10543 10761 10569 10767
rect 10711 10793 10737 10799
rect 10711 10761 10737 10767
rect 10991 10793 11017 10799
rect 10991 10761 11017 10767
rect 11271 10793 11297 10799
rect 11271 10761 11297 10767
rect 11383 10793 11409 10799
rect 11383 10761 11409 10767
rect 12111 10793 12137 10799
rect 12111 10761 12137 10767
rect 12335 10793 12361 10799
rect 12335 10761 12361 10767
rect 12615 10793 12641 10799
rect 13337 10767 13343 10793
rect 13369 10767 13375 10793
rect 12615 10761 12641 10767
rect 9311 10737 9337 10743
rect 5721 10711 5727 10737
rect 5753 10711 5759 10737
rect 7513 10711 7519 10737
rect 7545 10711 7551 10737
rect 8857 10711 8863 10737
rect 8889 10711 8895 10737
rect 9311 10705 9337 10711
rect 11327 10737 11353 10743
rect 14737 10711 14743 10737
rect 14769 10711 14775 10737
rect 11327 10705 11353 10711
rect 8023 10681 8049 10687
rect 8023 10649 8049 10655
rect 10319 10681 10345 10687
rect 10319 10649 10345 10655
rect 672 10597 20328 10614
rect 672 10571 2239 10597
rect 2265 10571 2291 10597
rect 2317 10571 2343 10597
rect 2369 10571 17599 10597
rect 17625 10571 17651 10597
rect 17677 10571 17703 10597
rect 17729 10571 20328 10597
rect 672 10554 20328 10571
rect 7295 10457 7321 10463
rect 7625 10431 7631 10457
rect 7657 10431 7663 10457
rect 7295 10425 7321 10431
rect 10375 10401 10401 10407
rect 10033 10375 10039 10401
rect 10065 10375 10071 10401
rect 10375 10369 10401 10375
rect 10655 10401 10681 10407
rect 10873 10375 10879 10401
rect 10905 10375 10911 10401
rect 11153 10375 11159 10401
rect 11185 10375 11191 10401
rect 10655 10369 10681 10375
rect 13393 10319 13399 10345
rect 13425 10319 13431 10345
rect 10319 10289 10345 10295
rect 10319 10257 10345 10263
rect 672 10205 20328 10222
rect 672 10179 9919 10205
rect 9945 10179 9971 10205
rect 9997 10179 10023 10205
rect 10049 10179 20328 10205
rect 672 10162 20328 10179
rect 8303 10121 8329 10127
rect 13001 10095 13007 10121
rect 13033 10095 13039 10121
rect 8303 10089 8329 10095
rect 7071 10065 7097 10071
rect 7071 10033 7097 10039
rect 7407 10065 7433 10071
rect 7407 10033 7433 10039
rect 7743 10065 7769 10071
rect 7743 10033 7769 10039
rect 8023 10065 8049 10071
rect 12279 10065 12305 10071
rect 11153 10039 11159 10065
rect 11185 10039 11191 10065
rect 8023 10033 8049 10039
rect 12279 10033 12305 10039
rect 12727 10065 12753 10071
rect 12727 10033 12753 10039
rect 12839 10065 12865 10071
rect 12839 10033 12865 10039
rect 6903 10009 6929 10015
rect 7687 10009 7713 10015
rect 7233 9983 7239 10009
rect 7265 9983 7271 10009
rect 6903 9977 6929 9983
rect 7687 9977 7713 9983
rect 7967 10009 7993 10015
rect 12223 10009 12249 10015
rect 8409 9983 8415 10009
rect 8441 9983 8447 10009
rect 9025 9983 9031 10009
rect 9057 9983 9063 10009
rect 9193 9983 9199 10009
rect 9225 9983 9231 10009
rect 9417 9983 9423 10009
rect 9449 9983 9455 10009
rect 12609 9983 12615 10009
rect 12641 9983 12647 10009
rect 13113 9983 13119 10009
rect 13145 9983 13151 10009
rect 13561 9983 13567 10009
rect 13593 9983 13599 10009
rect 7967 9977 7993 9983
rect 12223 9977 12249 9983
rect 6567 9953 6593 9959
rect 6567 9921 6593 9927
rect 13399 9953 13425 9959
rect 13953 9927 13959 9953
rect 13985 9927 13991 9953
rect 15017 9927 15023 9953
rect 15049 9927 15055 9953
rect 13399 9921 13425 9927
rect 7239 9897 7265 9903
rect 7239 9865 7265 9871
rect 7743 9897 7769 9903
rect 7743 9865 7769 9871
rect 8023 9897 8049 9903
rect 8023 9865 8049 9871
rect 8247 9897 8273 9903
rect 12279 9897 12305 9903
rect 9193 9871 9199 9897
rect 9225 9871 9231 9897
rect 8247 9865 8273 9871
rect 12279 9865 12305 9871
rect 12895 9897 12921 9903
rect 12895 9865 12921 9871
rect 672 9813 20328 9830
rect 672 9787 2239 9813
rect 2265 9787 2291 9813
rect 2317 9787 2343 9813
rect 2369 9787 17599 9813
rect 17625 9787 17651 9813
rect 17677 9787 17703 9813
rect 17729 9787 20328 9813
rect 672 9770 20328 9787
rect 7071 9729 7097 9735
rect 7071 9697 7097 9703
rect 11439 9729 11465 9735
rect 11439 9697 11465 9703
rect 12111 9729 12137 9735
rect 12111 9697 12137 9703
rect 967 9673 993 9679
rect 13343 9673 13369 9679
rect 4993 9647 4999 9673
rect 5025 9647 5031 9673
rect 7905 9647 7911 9673
rect 7937 9647 7943 9673
rect 967 9641 993 9647
rect 13343 9641 13369 9647
rect 13399 9673 13425 9679
rect 13735 9673 13761 9679
rect 13561 9647 13567 9673
rect 13593 9647 13599 9673
rect 13399 9641 13425 9647
rect 13735 9641 13761 9647
rect 13959 9673 13985 9679
rect 13959 9641 13985 9647
rect 14687 9673 14713 9679
rect 14687 9641 14713 9647
rect 20007 9673 20033 9679
rect 20007 9641 20033 9647
rect 7127 9617 7153 9623
rect 2137 9591 2143 9617
rect 2169 9591 2175 9617
rect 6393 9591 6399 9617
rect 6425 9591 6431 9617
rect 6953 9591 6959 9617
rect 6985 9591 6991 9617
rect 7127 9585 7153 9591
rect 7295 9617 7321 9623
rect 8639 9617 8665 9623
rect 9871 9617 9897 9623
rect 8017 9591 8023 9617
rect 8049 9591 8055 9617
rect 8745 9591 8751 9617
rect 8777 9591 8783 9617
rect 9249 9591 9255 9617
rect 9281 9591 9287 9617
rect 9417 9591 9423 9617
rect 9449 9591 9455 9617
rect 7295 9585 7321 9591
rect 8639 9585 8665 9591
rect 9871 9585 9897 9591
rect 10207 9617 10233 9623
rect 10207 9585 10233 9591
rect 10823 9617 10849 9623
rect 10823 9585 10849 9591
rect 11047 9617 11073 9623
rect 11047 9585 11073 9591
rect 11607 9617 11633 9623
rect 14631 9617 14657 9623
rect 11825 9591 11831 9617
rect 11857 9591 11863 9617
rect 12385 9591 12391 9617
rect 12417 9591 12423 9617
rect 12497 9591 12503 9617
rect 12529 9591 12535 9617
rect 14065 9591 14071 9617
rect 14097 9591 14103 9617
rect 18825 9591 18831 9617
rect 18857 9591 18863 9617
rect 11607 9585 11633 9591
rect 14631 9585 14657 9591
rect 8807 9561 8833 9567
rect 10655 9561 10681 9567
rect 6057 9535 6063 9561
rect 6089 9535 6095 9561
rect 7625 9535 7631 9561
rect 7657 9535 7663 9561
rect 9025 9535 9031 9561
rect 9057 9535 9063 9561
rect 9697 9535 9703 9561
rect 9729 9535 9735 9561
rect 8807 9529 8833 9535
rect 10655 9529 10681 9535
rect 11719 9561 11745 9567
rect 11719 9529 11745 9535
rect 13287 9561 13313 9567
rect 13287 9529 13313 9535
rect 13903 9561 13929 9567
rect 13903 9529 13929 9535
rect 6903 9505 6929 9511
rect 6903 9473 6929 9479
rect 7463 9505 7489 9511
rect 7463 9473 7489 9479
rect 7911 9505 7937 9511
rect 13063 9505 13089 9511
rect 9473 9479 9479 9505
rect 9505 9479 9511 9505
rect 10369 9479 10375 9505
rect 10401 9479 10407 9505
rect 7911 9473 7937 9479
rect 13063 9473 13089 9479
rect 13623 9505 13649 9511
rect 13623 9473 13649 9479
rect 672 9421 20328 9438
rect 672 9395 9919 9421
rect 9945 9395 9971 9421
rect 9997 9395 10023 9421
rect 10049 9395 20328 9421
rect 672 9378 20328 9395
rect 6791 9337 6817 9343
rect 6791 9305 6817 9311
rect 7519 9337 7545 9343
rect 8919 9337 8945 9343
rect 7905 9311 7911 9337
rect 7937 9311 7943 9337
rect 7519 9305 7545 9311
rect 8919 9305 8945 9311
rect 11103 9337 11129 9343
rect 11103 9305 11129 9311
rect 11327 9337 11353 9343
rect 11327 9305 11353 9311
rect 11439 9337 11465 9343
rect 11439 9305 11465 9311
rect 11551 9337 11577 9343
rect 12111 9337 12137 9343
rect 11769 9311 11775 9337
rect 11801 9311 11807 9337
rect 11551 9305 11577 9311
rect 12111 9305 12137 9311
rect 8695 9281 8721 9287
rect 7121 9255 7127 9281
rect 7153 9255 7159 9281
rect 8017 9255 8023 9281
rect 8049 9255 8055 9281
rect 9977 9255 9983 9281
rect 10009 9255 10015 9281
rect 10481 9255 10487 9281
rect 10513 9255 10519 9281
rect 12273 9255 12279 9281
rect 12305 9255 12311 9281
rect 8695 9249 8721 9255
rect 6735 9225 6761 9231
rect 5049 9199 5055 9225
rect 5081 9199 5087 9225
rect 6735 9193 6761 9199
rect 6959 9225 6985 9231
rect 6959 9193 6985 9199
rect 7407 9225 7433 9231
rect 8975 9225 9001 9231
rect 9591 9225 9617 9231
rect 7681 9199 7687 9225
rect 7713 9199 7719 9225
rect 8185 9199 8191 9225
rect 8217 9199 8223 9225
rect 8801 9199 8807 9225
rect 8833 9199 8839 9225
rect 9417 9199 9423 9225
rect 9449 9199 9455 9225
rect 9753 9199 9759 9225
rect 9785 9199 9791 9225
rect 10145 9199 10151 9225
rect 10177 9199 10183 9225
rect 10369 9199 10375 9225
rect 10401 9199 10407 9225
rect 10929 9199 10935 9225
rect 10961 9199 10967 9225
rect 11881 9199 11887 9225
rect 11913 9199 11919 9225
rect 13113 9199 13119 9225
rect 13145 9199 13151 9225
rect 18825 9199 18831 9225
rect 18857 9199 18863 9225
rect 7407 9193 7433 9199
rect 8975 9193 9001 9199
rect 9591 9193 9617 9199
rect 7463 9169 7489 9175
rect 5385 9143 5391 9169
rect 5417 9143 5423 9169
rect 6449 9143 6455 9169
rect 6481 9143 6487 9169
rect 7463 9137 7489 9143
rect 9311 9169 9337 9175
rect 11383 9169 11409 9175
rect 9697 9143 9703 9169
rect 9729 9143 9735 9169
rect 9311 9137 9337 9143
rect 11383 9137 11409 9143
rect 12951 9169 12977 9175
rect 13505 9143 13511 9169
rect 13537 9143 13543 9169
rect 14569 9143 14575 9169
rect 14601 9143 14607 9169
rect 12951 9137 12977 9143
rect 9255 9113 9281 9119
rect 9255 9081 9281 9087
rect 20007 9113 20033 9119
rect 20007 9081 20033 9087
rect 672 9029 20328 9046
rect 672 9003 2239 9029
rect 2265 9003 2291 9029
rect 2317 9003 2343 9029
rect 2369 9003 17599 9029
rect 17625 9003 17651 9029
rect 17677 9003 17703 9029
rect 17729 9003 20328 9029
rect 672 8986 20328 9003
rect 7127 8945 7153 8951
rect 8695 8945 8721 8951
rect 8017 8919 8023 8945
rect 8049 8919 8055 8945
rect 7127 8913 7153 8919
rect 8695 8913 8721 8919
rect 13791 8945 13817 8951
rect 13791 8913 13817 8919
rect 7631 8889 7657 8895
rect 8185 8863 8191 8889
rect 8217 8863 8223 8889
rect 7631 8857 7657 8863
rect 6791 8833 6817 8839
rect 6791 8801 6817 8807
rect 8135 8833 8161 8839
rect 9087 8833 9113 8839
rect 8521 8807 8527 8833
rect 8553 8807 8559 8833
rect 8135 8801 8161 8807
rect 9087 8801 9113 8807
rect 9255 8833 9281 8839
rect 9255 8801 9281 8807
rect 9871 8833 9897 8839
rect 9871 8801 9897 8807
rect 9983 8833 10009 8839
rect 9983 8801 10009 8807
rect 10207 8833 10233 8839
rect 10207 8801 10233 8807
rect 10655 8833 10681 8839
rect 10655 8801 10681 8807
rect 13063 8833 13089 8839
rect 13287 8833 13313 8839
rect 13847 8833 13873 8839
rect 13169 8807 13175 8833
rect 13201 8807 13207 8833
rect 13337 8807 13343 8833
rect 13369 8807 13375 8833
rect 13953 8807 13959 8833
rect 13985 8807 13991 8833
rect 13063 8801 13089 8807
rect 13287 8801 13313 8807
rect 13847 8801 13873 8807
rect 6847 8777 6873 8783
rect 6847 8745 6873 8751
rect 7127 8777 7153 8783
rect 7127 8745 7153 8751
rect 7183 8777 7209 8783
rect 7183 8745 7209 8751
rect 9143 8777 9169 8783
rect 9143 8745 9169 8751
rect 10711 8777 10737 8783
rect 10711 8745 10737 8751
rect 6455 8721 6481 8727
rect 6455 8689 6481 8695
rect 6959 8721 6985 8727
rect 6959 8689 6985 8695
rect 7351 8721 7377 8727
rect 7351 8689 7377 8695
rect 8639 8721 8665 8727
rect 8639 8689 8665 8695
rect 9927 8721 9953 8727
rect 9927 8689 9953 8695
rect 10823 8721 10849 8727
rect 10823 8689 10849 8695
rect 13455 8721 13481 8727
rect 13455 8689 13481 8695
rect 672 8637 20328 8654
rect 672 8611 9919 8637
rect 9945 8611 9971 8637
rect 9997 8611 10023 8637
rect 10049 8611 20328 8637
rect 672 8594 20328 8611
rect 7239 8553 7265 8559
rect 8247 8553 8273 8559
rect 7737 8527 7743 8553
rect 7769 8527 7775 8553
rect 10593 8527 10599 8553
rect 10625 8527 10631 8553
rect 7239 8521 7265 8527
rect 8247 8521 8273 8527
rect 7351 8497 7377 8503
rect 7905 8471 7911 8497
rect 7937 8471 7943 8497
rect 8409 8471 8415 8497
rect 8441 8471 8447 8497
rect 10705 8471 10711 8497
rect 10737 8471 10743 8497
rect 7351 8465 7377 8471
rect 7407 8441 7433 8447
rect 8079 8441 8105 8447
rect 7625 8415 7631 8441
rect 7657 8415 7663 8441
rect 7407 8409 7433 8415
rect 8079 8409 8105 8415
rect 8863 8441 8889 8447
rect 8863 8409 8889 8415
rect 9143 8441 9169 8447
rect 10033 8415 10039 8441
rect 10065 8415 10071 8441
rect 10201 8415 10207 8441
rect 10233 8415 10239 8441
rect 10649 8415 10655 8441
rect 10681 8415 10687 8441
rect 9143 8409 9169 8415
rect 13007 8385 13033 8391
rect 13007 8353 13033 8359
rect 672 8245 20328 8262
rect 672 8219 2239 8245
rect 2265 8219 2291 8245
rect 2317 8219 2343 8245
rect 2369 8219 17599 8245
rect 17625 8219 17651 8245
rect 17677 8219 17703 8245
rect 17729 8219 20328 8245
rect 672 8202 20328 8219
rect 7687 8161 7713 8167
rect 7687 8129 7713 8135
rect 7855 8161 7881 8167
rect 7855 8129 7881 8135
rect 7631 8105 7657 8111
rect 7631 8073 7657 8079
rect 7911 8105 7937 8111
rect 7911 8073 7937 8079
rect 20007 8105 20033 8111
rect 20007 8073 20033 8079
rect 7295 8049 7321 8055
rect 12727 8049 12753 8055
rect 9529 8023 9535 8049
rect 9561 8023 9567 8049
rect 7295 8017 7321 8023
rect 12727 8017 12753 8023
rect 12895 8049 12921 8055
rect 12895 8017 12921 8023
rect 13287 8049 13313 8055
rect 18937 8023 18943 8049
rect 18969 8023 18975 8049
rect 13287 8017 13313 8023
rect 13007 7993 13033 7999
rect 7457 7967 7463 7993
rect 7489 7967 7495 7993
rect 13007 7961 13033 7967
rect 13119 7993 13145 7999
rect 13119 7961 13145 7967
rect 13567 7993 13593 7999
rect 13567 7961 13593 7967
rect 13791 7993 13817 7999
rect 13791 7961 13817 7967
rect 11271 7937 11297 7943
rect 12783 7937 12809 7943
rect 9417 7911 9423 7937
rect 9449 7911 9455 7937
rect 11433 7911 11439 7937
rect 11465 7911 11471 7937
rect 11271 7905 11297 7911
rect 12783 7905 12809 7911
rect 12839 7937 12865 7943
rect 12839 7905 12865 7911
rect 13231 7937 13257 7943
rect 13231 7905 13257 7911
rect 13399 7937 13425 7943
rect 13399 7905 13425 7911
rect 13511 7937 13537 7943
rect 13511 7905 13537 7911
rect 672 7853 20328 7870
rect 672 7827 9919 7853
rect 9945 7827 9971 7853
rect 9997 7827 10023 7853
rect 10049 7827 20328 7853
rect 672 7810 20328 7827
rect 9647 7769 9673 7775
rect 11271 7769 11297 7775
rect 9473 7743 9479 7769
rect 9505 7743 9511 7769
rect 10481 7743 10487 7769
rect 10513 7743 10519 7769
rect 9647 7737 9673 7743
rect 11271 7737 11297 7743
rect 12111 7769 12137 7775
rect 12111 7737 12137 7743
rect 12223 7769 12249 7775
rect 12223 7737 12249 7743
rect 10767 7713 10793 7719
rect 5945 7687 5951 7713
rect 5977 7687 5983 7713
rect 10767 7681 10793 7687
rect 10879 7713 10905 7719
rect 10879 7681 10905 7687
rect 11383 7713 11409 7719
rect 11383 7681 11409 7687
rect 11999 7713 12025 7719
rect 13169 7687 13175 7713
rect 13201 7687 13207 7713
rect 11999 7681 12025 7687
rect 11103 7657 11129 7663
rect 5609 7631 5615 7657
rect 5641 7631 5647 7657
rect 10369 7631 10375 7657
rect 10401 7631 10407 7657
rect 11103 7625 11129 7631
rect 11327 7657 11353 7663
rect 11327 7625 11353 7631
rect 11495 7657 11521 7663
rect 11495 7625 11521 7631
rect 11607 7657 11633 7663
rect 12329 7631 12335 7657
rect 12361 7631 12367 7657
rect 12777 7631 12783 7657
rect 12809 7631 12815 7657
rect 18825 7631 18831 7657
rect 18857 7631 18863 7657
rect 11607 7625 11633 7631
rect 7239 7601 7265 7607
rect 7009 7575 7015 7601
rect 7041 7575 7047 7601
rect 7239 7569 7265 7575
rect 10991 7601 11017 7607
rect 10991 7569 11017 7575
rect 12167 7601 12193 7607
rect 14463 7601 14489 7607
rect 14233 7575 14239 7601
rect 14265 7575 14271 7601
rect 12167 7569 12193 7575
rect 14463 7569 14489 7575
rect 20007 7601 20033 7607
rect 20007 7569 20033 7575
rect 672 7461 20328 7478
rect 672 7435 2239 7461
rect 2265 7435 2291 7461
rect 2317 7435 2343 7461
rect 2369 7435 17599 7461
rect 17625 7435 17651 7461
rect 17677 7435 17703 7461
rect 17729 7435 20328 7461
rect 672 7418 20328 7435
rect 14295 7321 14321 7327
rect 8185 7295 8191 7321
rect 8217 7295 8223 7321
rect 11041 7295 11047 7321
rect 11073 7295 11079 7321
rect 12105 7295 12111 7321
rect 12137 7295 12143 7321
rect 13001 7295 13007 7321
rect 13033 7295 13039 7321
rect 14065 7295 14071 7321
rect 14097 7295 14103 7321
rect 14295 7289 14321 7295
rect 9199 7265 9225 7271
rect 6785 7239 6791 7265
rect 6817 7239 6823 7265
rect 9199 7233 9225 7239
rect 9255 7265 9281 7271
rect 9255 7233 9281 7239
rect 9367 7265 9393 7271
rect 9367 7233 9393 7239
rect 9423 7265 9449 7271
rect 9423 7233 9449 7239
rect 9647 7265 9673 7271
rect 9647 7233 9673 7239
rect 9759 7265 9785 7271
rect 9759 7233 9785 7239
rect 10039 7265 10065 7271
rect 10039 7233 10065 7239
rect 10375 7265 10401 7271
rect 12335 7265 12361 7271
rect 10705 7239 10711 7265
rect 10737 7239 10743 7265
rect 12609 7239 12615 7265
rect 12641 7239 12647 7265
rect 10375 7233 10401 7239
rect 12335 7233 12361 7239
rect 9927 7209 9953 7215
rect 7121 7183 7127 7209
rect 7153 7183 7159 7209
rect 9927 7177 9953 7183
rect 10263 7209 10289 7215
rect 10263 7177 10289 7183
rect 8415 7153 8441 7159
rect 8415 7121 8441 7127
rect 8975 7153 9001 7159
rect 8975 7121 9001 7127
rect 9311 7153 9337 7159
rect 9311 7121 9337 7127
rect 9703 7153 9729 7159
rect 9703 7121 9729 7127
rect 10151 7153 10177 7159
rect 10151 7121 10177 7127
rect 672 7069 20328 7086
rect 672 7043 9919 7069
rect 9945 7043 9971 7069
rect 9997 7043 10023 7069
rect 10049 7043 20328 7069
rect 672 7026 20328 7043
rect 11601 6959 11607 6985
rect 11633 6959 11639 6985
rect 8247 6929 8273 6935
rect 11439 6929 11465 6935
rect 9585 6903 9591 6929
rect 9617 6903 9623 6929
rect 8247 6897 8273 6903
rect 11439 6897 11465 6903
rect 8415 6873 8441 6879
rect 8919 6873 8945 6879
rect 8745 6847 8751 6873
rect 8777 6847 8783 6873
rect 8415 6841 8441 6847
rect 8919 6841 8945 6847
rect 9031 6873 9057 6879
rect 12167 6873 12193 6879
rect 9249 6847 9255 6873
rect 9281 6847 9287 6873
rect 11545 6847 11551 6873
rect 11577 6847 11583 6873
rect 11825 6847 11831 6873
rect 11857 6847 11863 6873
rect 9031 6841 9057 6847
rect 12167 6841 12193 6847
rect 12223 6817 12249 6823
rect 10649 6791 10655 6817
rect 10681 6791 10687 6817
rect 12223 6785 12249 6791
rect 11713 6735 11719 6761
rect 11745 6735 11751 6761
rect 672 6677 20328 6694
rect 672 6651 2239 6677
rect 2265 6651 2291 6677
rect 2317 6651 2343 6677
rect 2369 6651 17599 6677
rect 17625 6651 17651 6677
rect 17677 6651 17703 6677
rect 17729 6651 20328 6677
rect 672 6634 20328 6651
rect 9311 6593 9337 6599
rect 9311 6561 9337 6567
rect 9367 6537 9393 6543
rect 8073 6511 8079 6537
rect 8105 6511 8111 6537
rect 9137 6511 9143 6537
rect 9169 6511 9175 6537
rect 9367 6505 9393 6511
rect 9647 6537 9673 6543
rect 12951 6537 12977 6543
rect 11601 6511 11607 6537
rect 11633 6511 11639 6537
rect 12665 6511 12671 6537
rect 12697 6511 12703 6537
rect 9647 6505 9673 6511
rect 12951 6505 12977 6511
rect 7737 6455 7743 6481
rect 7769 6455 7775 6481
rect 11209 6455 11215 6481
rect 11241 6455 11247 6481
rect 672 6285 20328 6302
rect 672 6259 9919 6285
rect 9945 6259 9971 6285
rect 9997 6259 10023 6285
rect 10049 6259 20328 6285
rect 672 6242 20328 6259
rect 672 5893 20328 5910
rect 672 5867 2239 5893
rect 2265 5867 2291 5893
rect 2317 5867 2343 5893
rect 2369 5867 17599 5893
rect 17625 5867 17651 5893
rect 17677 5867 17703 5893
rect 17729 5867 20328 5893
rect 672 5850 20328 5867
rect 672 5501 20328 5518
rect 672 5475 9919 5501
rect 9945 5475 9971 5501
rect 9997 5475 10023 5501
rect 10049 5475 20328 5501
rect 672 5458 20328 5475
rect 672 5109 20328 5126
rect 672 5083 2239 5109
rect 2265 5083 2291 5109
rect 2317 5083 2343 5109
rect 2369 5083 17599 5109
rect 17625 5083 17651 5109
rect 17677 5083 17703 5109
rect 17729 5083 20328 5109
rect 672 5066 20328 5083
rect 672 4717 20328 4734
rect 672 4691 9919 4717
rect 9945 4691 9971 4717
rect 9997 4691 10023 4717
rect 10049 4691 20328 4717
rect 672 4674 20328 4691
rect 672 4325 20328 4342
rect 672 4299 2239 4325
rect 2265 4299 2291 4325
rect 2317 4299 2343 4325
rect 2369 4299 17599 4325
rect 17625 4299 17651 4325
rect 17677 4299 17703 4325
rect 17729 4299 20328 4325
rect 672 4282 20328 4299
rect 672 3933 20328 3950
rect 672 3907 9919 3933
rect 9945 3907 9971 3933
rect 9997 3907 10023 3933
rect 10049 3907 20328 3933
rect 672 3890 20328 3907
rect 672 3541 20328 3558
rect 672 3515 2239 3541
rect 2265 3515 2291 3541
rect 2317 3515 2343 3541
rect 2369 3515 17599 3541
rect 17625 3515 17651 3541
rect 17677 3515 17703 3541
rect 17729 3515 20328 3541
rect 672 3498 20328 3515
rect 672 3149 20328 3166
rect 672 3123 9919 3149
rect 9945 3123 9971 3149
rect 9997 3123 10023 3149
rect 10049 3123 20328 3149
rect 672 3106 20328 3123
rect 672 2757 20328 2774
rect 672 2731 2239 2757
rect 2265 2731 2291 2757
rect 2317 2731 2343 2757
rect 2369 2731 17599 2757
rect 17625 2731 17651 2757
rect 17677 2731 17703 2757
rect 17729 2731 20328 2757
rect 672 2714 20328 2731
rect 672 2365 20328 2382
rect 672 2339 9919 2365
rect 9945 2339 9971 2365
rect 9997 2339 10023 2365
rect 10049 2339 20328 2365
rect 672 2322 20328 2339
rect 12609 2143 12615 2169
rect 12641 2143 12647 2169
rect 13119 2057 13145 2063
rect 13119 2025 13145 2031
rect 672 1973 20328 1990
rect 672 1947 2239 1973
rect 2265 1947 2291 1973
rect 2317 1947 2343 1973
rect 2369 1947 17599 1973
rect 17625 1947 17651 1973
rect 17677 1947 17703 1973
rect 17729 1947 20328 1973
rect 672 1930 20328 1947
rect 9311 1833 9337 1839
rect 9311 1801 9337 1807
rect 11047 1833 11073 1839
rect 11047 1801 11073 1807
rect 12783 1833 12809 1839
rect 12783 1801 12809 1807
rect 8801 1751 8807 1777
rect 8833 1751 8839 1777
rect 10537 1751 10543 1777
rect 10569 1751 10575 1777
rect 12273 1751 12279 1777
rect 12305 1751 12311 1777
rect 17599 1665 17625 1671
rect 17599 1633 17625 1639
rect 672 1581 20328 1598
rect 672 1555 9919 1581
rect 9945 1555 9971 1581
rect 9997 1555 10023 1581
rect 10049 1555 20328 1581
rect 672 1538 20328 1555
<< via1 >>
rect 2239 19195 2265 19221
rect 2291 19195 2317 19221
rect 2343 19195 2369 19221
rect 17599 19195 17625 19221
rect 17651 19195 17677 19221
rect 17703 19195 17729 19221
rect 11047 19111 11073 19137
rect 12783 19111 12809 19137
rect 9423 19055 9449 19081
rect 9031 18999 9057 19025
rect 10655 18999 10681 19025
rect 12279 18999 12305 19025
rect 9919 18803 9945 18829
rect 9971 18803 9997 18829
rect 10023 18803 10049 18829
rect 10711 18719 10737 18745
rect 13399 18719 13425 18745
rect 20119 18663 20145 18689
rect 10375 18607 10401 18633
rect 13007 18607 13033 18633
rect 2239 18411 2265 18437
rect 2291 18411 2317 18437
rect 2343 18411 2369 18437
rect 17599 18411 17625 18437
rect 17651 18411 17677 18437
rect 17703 18411 17729 18437
rect 9919 18019 9945 18045
rect 9971 18019 9997 18045
rect 10023 18019 10049 18045
rect 2239 17627 2265 17653
rect 2291 17627 2317 17653
rect 2343 17627 2369 17653
rect 17599 17627 17625 17653
rect 17651 17627 17677 17653
rect 17703 17627 17729 17653
rect 20119 17319 20145 17345
rect 9919 17235 9945 17261
rect 9971 17235 9997 17261
rect 10023 17235 10049 17261
rect 2239 16843 2265 16869
rect 2291 16843 2317 16869
rect 2343 16843 2369 16869
rect 17599 16843 17625 16869
rect 17651 16843 17677 16869
rect 17703 16843 17729 16869
rect 9919 16451 9945 16477
rect 9971 16451 9997 16477
rect 10023 16451 10049 16477
rect 2239 16059 2265 16085
rect 2291 16059 2317 16085
rect 2343 16059 2369 16085
rect 17599 16059 17625 16085
rect 17651 16059 17677 16085
rect 17703 16059 17729 16085
rect 9919 15667 9945 15693
rect 9971 15667 9997 15693
rect 10023 15667 10049 15693
rect 2239 15275 2265 15301
rect 2291 15275 2317 15301
rect 2343 15275 2369 15301
rect 17599 15275 17625 15301
rect 17651 15275 17677 15301
rect 17703 15275 17729 15301
rect 9919 14883 9945 14909
rect 9971 14883 9997 14909
rect 10023 14883 10049 14909
rect 2239 14491 2265 14517
rect 2291 14491 2317 14517
rect 2343 14491 2369 14517
rect 17599 14491 17625 14517
rect 17651 14491 17677 14517
rect 17703 14491 17729 14517
rect 9919 14099 9945 14125
rect 9971 14099 9997 14125
rect 10023 14099 10049 14125
rect 18943 13903 18969 13929
rect 12951 13847 12977 13873
rect 19951 13847 19977 13873
rect 2239 13707 2265 13733
rect 2291 13707 2317 13733
rect 2343 13707 2369 13733
rect 17599 13707 17625 13733
rect 17651 13707 17677 13733
rect 17703 13707 17729 13733
rect 967 13567 993 13593
rect 10375 13567 10401 13593
rect 12783 13567 12809 13593
rect 20007 13567 20033 13593
rect 2143 13511 2169 13537
rect 8975 13511 9001 13537
rect 10767 13511 10793 13537
rect 11383 13511 11409 13537
rect 12895 13511 12921 13537
rect 13343 13511 13369 13537
rect 18831 13511 18857 13537
rect 8751 13455 8777 13481
rect 9311 13455 9337 13481
rect 10655 13455 10681 13481
rect 11103 13455 11129 13481
rect 11159 13455 11185 13481
rect 11719 13455 11745 13481
rect 13007 13455 13033 13481
rect 13063 13455 13089 13481
rect 13399 13455 13425 13481
rect 10991 13399 11017 13425
rect 13511 13399 13537 13425
rect 9919 13315 9945 13341
rect 9971 13315 9997 13341
rect 10023 13315 10049 13341
rect 9703 13231 9729 13257
rect 9927 13231 9953 13257
rect 10095 13231 10121 13257
rect 11831 13231 11857 13257
rect 9199 13175 9225 13201
rect 11943 13175 11969 13201
rect 11999 13175 12025 13201
rect 12951 13175 12977 13201
rect 13007 13175 13033 13201
rect 14799 13175 14825 13201
rect 14967 13175 14993 13201
rect 2143 13119 2169 13145
rect 8023 13119 8049 13145
rect 9143 13119 9169 13145
rect 9311 13119 9337 13145
rect 9647 13119 9673 13145
rect 9815 13119 9841 13145
rect 10319 13119 10345 13145
rect 12839 13119 12865 13145
rect 13175 13119 13201 13145
rect 18831 13119 18857 13145
rect 6623 13063 6649 13089
rect 7687 13063 7713 13089
rect 8303 13063 8329 13089
rect 10655 13063 10681 13089
rect 11719 13063 11745 13089
rect 12223 13063 12249 13089
rect 12727 13063 12753 13089
rect 13567 13063 13593 13089
rect 14631 13063 14657 13089
rect 967 13007 993 13033
rect 20007 13007 20033 13033
rect 2239 12923 2265 12949
rect 2291 12923 2317 12949
rect 2343 12923 2369 12949
rect 17599 12923 17625 12949
rect 17651 12923 17677 12949
rect 17703 12923 17729 12949
rect 10095 12839 10121 12865
rect 7295 12783 7321 12809
rect 7575 12783 7601 12809
rect 9479 12783 9505 12809
rect 10375 12783 10401 12809
rect 13511 12783 13537 12809
rect 7631 12727 7657 12753
rect 8023 12727 8049 12753
rect 9815 12727 9841 12753
rect 10151 12727 10177 12753
rect 10879 12727 10905 12753
rect 11047 12727 11073 12753
rect 12111 12727 12137 12753
rect 13623 12727 13649 12753
rect 13791 12727 13817 12753
rect 6847 12671 6873 12697
rect 7351 12671 7377 12697
rect 7855 12671 7881 12697
rect 8415 12671 8441 12697
rect 12447 12671 12473 12697
rect 6903 12615 6929 12641
rect 7575 12615 7601 12641
rect 7743 12615 7769 12641
rect 9927 12615 9953 12641
rect 10039 12615 10065 12641
rect 10991 12615 11017 12641
rect 13735 12615 13761 12641
rect 14015 12615 14041 12641
rect 9919 12531 9945 12557
rect 9971 12531 9997 12557
rect 10023 12531 10049 12557
rect 7631 12447 7657 12473
rect 7743 12447 7769 12473
rect 9031 12447 9057 12473
rect 9423 12447 9449 12473
rect 12559 12447 12585 12473
rect 7015 12391 7041 12417
rect 12671 12391 12697 12417
rect 12727 12391 12753 12417
rect 7407 12335 7433 12361
rect 7687 12335 7713 12361
rect 7799 12335 7825 12361
rect 7911 12335 7937 12361
rect 8975 12335 9001 12361
rect 9087 12335 9113 12361
rect 9311 12335 9337 12361
rect 9535 12335 9561 12361
rect 9815 12335 9841 12361
rect 5951 12279 5977 12305
rect 2239 12139 2265 12165
rect 2291 12139 2317 12165
rect 2343 12139 2369 12165
rect 17599 12139 17625 12165
rect 17651 12139 17677 12165
rect 17703 12139 17729 12165
rect 967 11999 993 12025
rect 7687 11999 7713 12025
rect 12391 11999 12417 12025
rect 2143 11943 2169 11969
rect 7463 11943 7489 11969
rect 9759 11943 9785 11969
rect 7407 11887 7433 11913
rect 9591 11887 9617 11913
rect 7295 11831 7321 11857
rect 9647 11831 9673 11857
rect 9919 11747 9945 11773
rect 9971 11747 9997 11773
rect 10023 11747 10049 11773
rect 7351 11663 7377 11689
rect 8919 11663 8945 11689
rect 10207 11663 10233 11689
rect 10319 11663 10345 11689
rect 14631 11663 14657 11689
rect 8863 11607 8889 11633
rect 12727 11607 12753 11633
rect 7127 11551 7153 11577
rect 7519 11551 7545 11577
rect 7631 11551 7657 11577
rect 7743 11551 7769 11577
rect 9031 11551 9057 11577
rect 10151 11551 10177 11577
rect 11999 11551 12025 11577
rect 12111 11551 12137 11577
rect 12279 11551 12305 11577
rect 12783 11551 12809 11577
rect 13007 11551 13033 11577
rect 18831 11551 18857 11577
rect 5671 11495 5697 11521
rect 6735 11495 6761 11521
rect 7575 11495 7601 11521
rect 9871 11495 9897 11521
rect 12055 11495 12081 11521
rect 13343 11495 13369 11521
rect 14407 11495 14433 11521
rect 9927 11439 9953 11465
rect 12727 11439 12753 11465
rect 20007 11439 20033 11465
rect 2239 11355 2265 11381
rect 2291 11355 2317 11381
rect 2343 11355 2369 11381
rect 17599 11355 17625 11381
rect 17651 11355 17677 11381
rect 17703 11355 17729 11381
rect 10151 11271 10177 11297
rect 967 11215 993 11241
rect 9031 11215 9057 11241
rect 12223 11215 12249 11241
rect 13343 11215 13369 11241
rect 20007 11215 20033 11241
rect 2143 11159 2169 11185
rect 7071 11159 7097 11185
rect 7295 11159 7321 11185
rect 7631 11159 7657 11185
rect 7967 11159 7993 11185
rect 8639 11159 8665 11185
rect 8863 11159 8889 11185
rect 9927 11159 9953 11185
rect 10823 11159 10849 11185
rect 12559 11159 12585 11185
rect 12671 11159 12697 11185
rect 12895 11159 12921 11185
rect 13231 11159 13257 11185
rect 13791 11159 13817 11185
rect 18831 11159 18857 11185
rect 7799 11103 7825 11129
rect 8695 11103 8721 11129
rect 8975 11103 9001 11129
rect 9255 11103 9281 11129
rect 9815 11103 9841 11129
rect 11159 11103 11185 11129
rect 13511 11103 13537 11129
rect 13623 11103 13649 11129
rect 7351 11047 7377 11073
rect 7407 11047 7433 11073
rect 7743 11047 7769 11073
rect 9423 11047 9449 11073
rect 10319 11047 10345 11073
rect 12727 11047 12753 11073
rect 12783 11047 12809 11073
rect 13063 11047 13089 11073
rect 13679 11047 13705 11073
rect 9919 10963 9945 10989
rect 9971 10963 9997 10989
rect 10023 10963 10049 10989
rect 8247 10879 8273 10905
rect 8751 10879 8777 10905
rect 10039 10879 10065 10905
rect 11159 10879 11185 10905
rect 11495 10879 11521 10905
rect 11887 10879 11913 10905
rect 11999 10879 12025 10905
rect 12167 10879 12193 10905
rect 12671 10879 12697 10905
rect 6791 10823 6817 10849
rect 7463 10823 7489 10849
rect 7967 10823 7993 10849
rect 8023 10823 8049 10849
rect 9703 10823 9729 10849
rect 9927 10823 9953 10849
rect 10319 10823 10345 10849
rect 10599 10823 10625 10849
rect 11047 10823 11073 10849
rect 11775 10823 11801 10849
rect 12727 10823 12753 10849
rect 12783 10823 12809 10849
rect 12895 10823 12921 10849
rect 13679 10823 13705 10849
rect 7127 10767 7153 10793
rect 7575 10767 7601 10793
rect 7743 10767 7769 10793
rect 8359 10767 8385 10793
rect 8807 10767 8833 10793
rect 9535 10767 9561 10793
rect 10263 10767 10289 10793
rect 10543 10767 10569 10793
rect 10711 10767 10737 10793
rect 10991 10767 11017 10793
rect 11271 10767 11297 10793
rect 11383 10767 11409 10793
rect 12111 10767 12137 10793
rect 12335 10767 12361 10793
rect 12615 10767 12641 10793
rect 13343 10767 13369 10793
rect 5727 10711 5753 10737
rect 7519 10711 7545 10737
rect 8863 10711 8889 10737
rect 9311 10711 9337 10737
rect 11327 10711 11353 10737
rect 14743 10711 14769 10737
rect 8023 10655 8049 10681
rect 10319 10655 10345 10681
rect 2239 10571 2265 10597
rect 2291 10571 2317 10597
rect 2343 10571 2369 10597
rect 17599 10571 17625 10597
rect 17651 10571 17677 10597
rect 17703 10571 17729 10597
rect 7295 10431 7321 10457
rect 7631 10431 7657 10457
rect 10039 10375 10065 10401
rect 10375 10375 10401 10401
rect 10655 10375 10681 10401
rect 10879 10375 10905 10401
rect 11159 10375 11185 10401
rect 13399 10319 13425 10345
rect 10319 10263 10345 10289
rect 9919 10179 9945 10205
rect 9971 10179 9997 10205
rect 10023 10179 10049 10205
rect 8303 10095 8329 10121
rect 13007 10095 13033 10121
rect 7071 10039 7097 10065
rect 7407 10039 7433 10065
rect 7743 10039 7769 10065
rect 8023 10039 8049 10065
rect 11159 10039 11185 10065
rect 12279 10039 12305 10065
rect 12727 10039 12753 10065
rect 12839 10039 12865 10065
rect 6903 9983 6929 10009
rect 7239 9983 7265 10009
rect 7687 9983 7713 10009
rect 7967 9983 7993 10009
rect 8415 9983 8441 10009
rect 9031 9983 9057 10009
rect 9199 9983 9225 10009
rect 9423 9983 9449 10009
rect 12223 9983 12249 10009
rect 12615 9983 12641 10009
rect 13119 9983 13145 10009
rect 13567 9983 13593 10009
rect 6567 9927 6593 9953
rect 13399 9927 13425 9953
rect 13959 9927 13985 9953
rect 15023 9927 15049 9953
rect 7239 9871 7265 9897
rect 7743 9871 7769 9897
rect 8023 9871 8049 9897
rect 8247 9871 8273 9897
rect 9199 9871 9225 9897
rect 12279 9871 12305 9897
rect 12895 9871 12921 9897
rect 2239 9787 2265 9813
rect 2291 9787 2317 9813
rect 2343 9787 2369 9813
rect 17599 9787 17625 9813
rect 17651 9787 17677 9813
rect 17703 9787 17729 9813
rect 7071 9703 7097 9729
rect 11439 9703 11465 9729
rect 12111 9703 12137 9729
rect 967 9647 993 9673
rect 4999 9647 5025 9673
rect 7911 9647 7937 9673
rect 13343 9647 13369 9673
rect 13399 9647 13425 9673
rect 13567 9647 13593 9673
rect 13735 9647 13761 9673
rect 13959 9647 13985 9673
rect 14687 9647 14713 9673
rect 20007 9647 20033 9673
rect 2143 9591 2169 9617
rect 6399 9591 6425 9617
rect 6959 9591 6985 9617
rect 7127 9591 7153 9617
rect 7295 9591 7321 9617
rect 8023 9591 8049 9617
rect 8639 9591 8665 9617
rect 8751 9591 8777 9617
rect 9255 9591 9281 9617
rect 9423 9591 9449 9617
rect 9871 9591 9897 9617
rect 10207 9591 10233 9617
rect 10823 9591 10849 9617
rect 11047 9591 11073 9617
rect 11607 9591 11633 9617
rect 11831 9591 11857 9617
rect 12391 9591 12417 9617
rect 12503 9591 12529 9617
rect 14071 9591 14097 9617
rect 14631 9591 14657 9617
rect 18831 9591 18857 9617
rect 6063 9535 6089 9561
rect 7631 9535 7657 9561
rect 8807 9535 8833 9561
rect 9031 9535 9057 9561
rect 9703 9535 9729 9561
rect 10655 9535 10681 9561
rect 11719 9535 11745 9561
rect 13287 9535 13313 9561
rect 13903 9535 13929 9561
rect 6903 9479 6929 9505
rect 7463 9479 7489 9505
rect 7911 9479 7937 9505
rect 9479 9479 9505 9505
rect 10375 9479 10401 9505
rect 13063 9479 13089 9505
rect 13623 9479 13649 9505
rect 9919 9395 9945 9421
rect 9971 9395 9997 9421
rect 10023 9395 10049 9421
rect 6791 9311 6817 9337
rect 7519 9311 7545 9337
rect 7911 9311 7937 9337
rect 8919 9311 8945 9337
rect 11103 9311 11129 9337
rect 11327 9311 11353 9337
rect 11439 9311 11465 9337
rect 11551 9311 11577 9337
rect 11775 9311 11801 9337
rect 12111 9311 12137 9337
rect 7127 9255 7153 9281
rect 8023 9255 8049 9281
rect 8695 9255 8721 9281
rect 9983 9255 10009 9281
rect 10487 9255 10513 9281
rect 12279 9255 12305 9281
rect 5055 9199 5081 9225
rect 6735 9199 6761 9225
rect 6959 9199 6985 9225
rect 7407 9199 7433 9225
rect 7687 9199 7713 9225
rect 8191 9199 8217 9225
rect 8807 9199 8833 9225
rect 8975 9199 9001 9225
rect 9423 9199 9449 9225
rect 9591 9199 9617 9225
rect 9759 9199 9785 9225
rect 10151 9199 10177 9225
rect 10375 9199 10401 9225
rect 10935 9199 10961 9225
rect 11887 9199 11913 9225
rect 13119 9199 13145 9225
rect 18831 9199 18857 9225
rect 5391 9143 5417 9169
rect 6455 9143 6481 9169
rect 7463 9143 7489 9169
rect 9311 9143 9337 9169
rect 9703 9143 9729 9169
rect 11383 9143 11409 9169
rect 12951 9143 12977 9169
rect 13511 9143 13537 9169
rect 14575 9143 14601 9169
rect 9255 9087 9281 9113
rect 20007 9087 20033 9113
rect 2239 9003 2265 9029
rect 2291 9003 2317 9029
rect 2343 9003 2369 9029
rect 17599 9003 17625 9029
rect 17651 9003 17677 9029
rect 17703 9003 17729 9029
rect 7127 8919 7153 8945
rect 8023 8919 8049 8945
rect 8695 8919 8721 8945
rect 13791 8919 13817 8945
rect 7631 8863 7657 8889
rect 8191 8863 8217 8889
rect 6791 8807 6817 8833
rect 8135 8807 8161 8833
rect 8527 8807 8553 8833
rect 9087 8807 9113 8833
rect 9255 8807 9281 8833
rect 9871 8807 9897 8833
rect 9983 8807 10009 8833
rect 10207 8807 10233 8833
rect 10655 8807 10681 8833
rect 13063 8807 13089 8833
rect 13175 8807 13201 8833
rect 13287 8807 13313 8833
rect 13343 8807 13369 8833
rect 13847 8807 13873 8833
rect 13959 8807 13985 8833
rect 6847 8751 6873 8777
rect 7127 8751 7153 8777
rect 7183 8751 7209 8777
rect 9143 8751 9169 8777
rect 10711 8751 10737 8777
rect 6455 8695 6481 8721
rect 6959 8695 6985 8721
rect 7351 8695 7377 8721
rect 8639 8695 8665 8721
rect 9927 8695 9953 8721
rect 10823 8695 10849 8721
rect 13455 8695 13481 8721
rect 9919 8611 9945 8637
rect 9971 8611 9997 8637
rect 10023 8611 10049 8637
rect 7239 8527 7265 8553
rect 7743 8527 7769 8553
rect 8247 8527 8273 8553
rect 10599 8527 10625 8553
rect 7351 8471 7377 8497
rect 7911 8471 7937 8497
rect 8415 8471 8441 8497
rect 10711 8471 10737 8497
rect 7407 8415 7433 8441
rect 7631 8415 7657 8441
rect 8079 8415 8105 8441
rect 8863 8415 8889 8441
rect 9143 8415 9169 8441
rect 10039 8415 10065 8441
rect 10207 8415 10233 8441
rect 10655 8415 10681 8441
rect 13007 8359 13033 8385
rect 2239 8219 2265 8245
rect 2291 8219 2317 8245
rect 2343 8219 2369 8245
rect 17599 8219 17625 8245
rect 17651 8219 17677 8245
rect 17703 8219 17729 8245
rect 7687 8135 7713 8161
rect 7855 8135 7881 8161
rect 7631 8079 7657 8105
rect 7911 8079 7937 8105
rect 20007 8079 20033 8105
rect 7295 8023 7321 8049
rect 9535 8023 9561 8049
rect 12727 8023 12753 8049
rect 12895 8023 12921 8049
rect 13287 8023 13313 8049
rect 18943 8023 18969 8049
rect 7463 7967 7489 7993
rect 13007 7967 13033 7993
rect 13119 7967 13145 7993
rect 13567 7967 13593 7993
rect 13791 7967 13817 7993
rect 9423 7911 9449 7937
rect 11271 7911 11297 7937
rect 11439 7911 11465 7937
rect 12783 7911 12809 7937
rect 12839 7911 12865 7937
rect 13231 7911 13257 7937
rect 13399 7911 13425 7937
rect 13511 7911 13537 7937
rect 9919 7827 9945 7853
rect 9971 7827 9997 7853
rect 10023 7827 10049 7853
rect 9479 7743 9505 7769
rect 9647 7743 9673 7769
rect 10487 7743 10513 7769
rect 11271 7743 11297 7769
rect 12111 7743 12137 7769
rect 12223 7743 12249 7769
rect 5951 7687 5977 7713
rect 10767 7687 10793 7713
rect 10879 7687 10905 7713
rect 11383 7687 11409 7713
rect 11999 7687 12025 7713
rect 13175 7687 13201 7713
rect 5615 7631 5641 7657
rect 10375 7631 10401 7657
rect 11103 7631 11129 7657
rect 11327 7631 11353 7657
rect 11495 7631 11521 7657
rect 11607 7631 11633 7657
rect 12335 7631 12361 7657
rect 12783 7631 12809 7657
rect 18831 7631 18857 7657
rect 7015 7575 7041 7601
rect 7239 7575 7265 7601
rect 10991 7575 11017 7601
rect 12167 7575 12193 7601
rect 14239 7575 14265 7601
rect 14463 7575 14489 7601
rect 20007 7575 20033 7601
rect 2239 7435 2265 7461
rect 2291 7435 2317 7461
rect 2343 7435 2369 7461
rect 17599 7435 17625 7461
rect 17651 7435 17677 7461
rect 17703 7435 17729 7461
rect 8191 7295 8217 7321
rect 11047 7295 11073 7321
rect 12111 7295 12137 7321
rect 13007 7295 13033 7321
rect 14071 7295 14097 7321
rect 14295 7295 14321 7321
rect 6791 7239 6817 7265
rect 9199 7239 9225 7265
rect 9255 7239 9281 7265
rect 9367 7239 9393 7265
rect 9423 7239 9449 7265
rect 9647 7239 9673 7265
rect 9759 7239 9785 7265
rect 10039 7239 10065 7265
rect 10375 7239 10401 7265
rect 10711 7239 10737 7265
rect 12335 7239 12361 7265
rect 12615 7239 12641 7265
rect 7127 7183 7153 7209
rect 9927 7183 9953 7209
rect 10263 7183 10289 7209
rect 8415 7127 8441 7153
rect 8975 7127 9001 7153
rect 9311 7127 9337 7153
rect 9703 7127 9729 7153
rect 10151 7127 10177 7153
rect 9919 7043 9945 7069
rect 9971 7043 9997 7069
rect 10023 7043 10049 7069
rect 11607 6959 11633 6985
rect 8247 6903 8273 6929
rect 9591 6903 9617 6929
rect 11439 6903 11465 6929
rect 8415 6847 8441 6873
rect 8751 6847 8777 6873
rect 8919 6847 8945 6873
rect 9031 6847 9057 6873
rect 9255 6847 9281 6873
rect 11551 6847 11577 6873
rect 11831 6847 11857 6873
rect 12167 6847 12193 6873
rect 10655 6791 10681 6817
rect 12223 6791 12249 6817
rect 11719 6735 11745 6761
rect 2239 6651 2265 6677
rect 2291 6651 2317 6677
rect 2343 6651 2369 6677
rect 17599 6651 17625 6677
rect 17651 6651 17677 6677
rect 17703 6651 17729 6677
rect 9311 6567 9337 6593
rect 8079 6511 8105 6537
rect 9143 6511 9169 6537
rect 9367 6511 9393 6537
rect 9647 6511 9673 6537
rect 11607 6511 11633 6537
rect 12671 6511 12697 6537
rect 12951 6511 12977 6537
rect 7743 6455 7769 6481
rect 11215 6455 11241 6481
rect 9919 6259 9945 6285
rect 9971 6259 9997 6285
rect 10023 6259 10049 6285
rect 2239 5867 2265 5893
rect 2291 5867 2317 5893
rect 2343 5867 2369 5893
rect 17599 5867 17625 5893
rect 17651 5867 17677 5893
rect 17703 5867 17729 5893
rect 9919 5475 9945 5501
rect 9971 5475 9997 5501
rect 10023 5475 10049 5501
rect 2239 5083 2265 5109
rect 2291 5083 2317 5109
rect 2343 5083 2369 5109
rect 17599 5083 17625 5109
rect 17651 5083 17677 5109
rect 17703 5083 17729 5109
rect 9919 4691 9945 4717
rect 9971 4691 9997 4717
rect 10023 4691 10049 4717
rect 2239 4299 2265 4325
rect 2291 4299 2317 4325
rect 2343 4299 2369 4325
rect 17599 4299 17625 4325
rect 17651 4299 17677 4325
rect 17703 4299 17729 4325
rect 9919 3907 9945 3933
rect 9971 3907 9997 3933
rect 10023 3907 10049 3933
rect 2239 3515 2265 3541
rect 2291 3515 2317 3541
rect 2343 3515 2369 3541
rect 17599 3515 17625 3541
rect 17651 3515 17677 3541
rect 17703 3515 17729 3541
rect 9919 3123 9945 3149
rect 9971 3123 9997 3149
rect 10023 3123 10049 3149
rect 2239 2731 2265 2757
rect 2291 2731 2317 2757
rect 2343 2731 2369 2757
rect 17599 2731 17625 2757
rect 17651 2731 17677 2757
rect 17703 2731 17729 2757
rect 9919 2339 9945 2365
rect 9971 2339 9997 2365
rect 10023 2339 10049 2365
rect 12615 2143 12641 2169
rect 13119 2031 13145 2057
rect 2239 1947 2265 1973
rect 2291 1947 2317 1973
rect 2343 1947 2369 1973
rect 17599 1947 17625 1973
rect 17651 1947 17677 1973
rect 17703 1947 17729 1973
rect 9311 1807 9337 1833
rect 11047 1807 11073 1833
rect 12783 1807 12809 1833
rect 8807 1751 8833 1777
rect 10543 1751 10569 1777
rect 12279 1751 12305 1777
rect 17599 1639 17625 1665
rect 9919 1555 9945 1581
rect 9971 1555 9997 1581
rect 10023 1555 10049 1581
<< metal2 >>
rect 9408 20600 9464 21000
rect 10080 20600 10136 21000
rect 10416 20600 10472 21000
rect 11424 20600 11480 21000
rect 12768 20600 12824 21000
rect 2238 19222 2370 19227
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2238 19189 2370 19194
rect 9422 19081 9450 20600
rect 9422 19055 9423 19081
rect 9449 19055 9450 19081
rect 9422 19049 9450 19055
rect 9030 19025 9058 19031
rect 9030 18999 9031 19025
rect 9057 18999 9058 19025
rect 2238 18438 2370 18443
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2238 18405 2370 18410
rect 2238 17654 2370 17659
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2238 17621 2370 17626
rect 2238 16870 2370 16875
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2238 16837 2370 16842
rect 2238 16086 2370 16091
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2238 16053 2370 16058
rect 9030 15974 9058 18999
rect 9918 18830 10050 18835
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 9918 18797 10050 18802
rect 10094 18746 10122 20600
rect 10430 19138 10458 20600
rect 10430 19105 10458 19110
rect 11046 19138 11074 19143
rect 11046 19091 11074 19110
rect 11438 19138 11466 20600
rect 12782 19306 12810 20600
rect 12782 19273 12810 19278
rect 13398 19306 13426 19311
rect 11438 19105 11466 19110
rect 12782 19138 12810 19143
rect 12782 19091 12810 19110
rect 10094 18713 10122 18718
rect 10654 19025 10682 19031
rect 10654 18999 10655 19025
rect 10681 18999 10682 19025
rect 10374 18633 10402 18639
rect 10374 18607 10375 18633
rect 10401 18607 10402 18633
rect 9918 18046 10050 18051
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 9918 18013 10050 18018
rect 9918 17262 10050 17267
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 9918 17229 10050 17234
rect 9918 16478 10050 16483
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 9918 16445 10050 16450
rect 9030 15946 9226 15974
rect 2238 15302 2370 15307
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2238 15269 2370 15274
rect 2238 14518 2370 14523
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2238 14485 2370 14490
rect 2238 13734 2370 13739
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2238 13701 2370 13706
rect 966 13593 994 13599
rect 966 13567 967 13593
rect 993 13567 994 13593
rect 966 13146 994 13567
rect 2142 13538 2170 13543
rect 2142 13491 2170 13510
rect 6622 13538 6650 13543
rect 966 13113 994 13118
rect 2086 13482 2114 13487
rect 966 13033 994 13039
rect 966 13007 967 13033
rect 993 13007 994 13033
rect 966 12810 994 13007
rect 966 12777 994 12782
rect 966 12025 994 12031
rect 966 11999 967 12025
rect 993 11999 994 12025
rect 966 11802 994 11999
rect 966 11769 994 11774
rect 966 11242 994 11247
rect 966 11195 994 11214
rect 2086 10738 2114 13454
rect 2142 13146 2170 13151
rect 2142 13099 2170 13118
rect 5950 13146 5978 13151
rect 2238 12950 2370 12955
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2238 12917 2370 12922
rect 5950 12362 5978 13118
rect 6622 13090 6650 13510
rect 8974 13537 9002 13543
rect 8974 13511 8975 13537
rect 9001 13511 9002 13537
rect 8750 13482 8778 13487
rect 8974 13482 9002 13511
rect 8750 13481 9002 13482
rect 8750 13455 8751 13481
rect 8777 13455 9002 13481
rect 8750 13454 9002 13455
rect 8750 13449 8778 13454
rect 8022 13145 8050 13151
rect 8022 13119 8023 13145
rect 8049 13119 8050 13145
rect 6622 13043 6650 13062
rect 7630 13090 7658 13095
rect 7294 12810 7322 12815
rect 7574 12810 7602 12815
rect 7294 12809 7602 12810
rect 7294 12783 7295 12809
rect 7321 12783 7575 12809
rect 7601 12783 7602 12809
rect 7294 12782 7602 12783
rect 7294 12777 7322 12782
rect 7574 12777 7602 12782
rect 7630 12753 7658 13062
rect 7630 12727 7631 12753
rect 7657 12727 7658 12753
rect 7630 12721 7658 12727
rect 7686 13089 7714 13095
rect 7686 13063 7687 13089
rect 7713 13063 7714 13089
rect 7686 12754 7714 13063
rect 7686 12721 7714 12726
rect 8022 13090 8050 13119
rect 8022 12753 8050 13062
rect 8302 13090 8330 13095
rect 8302 13043 8330 13062
rect 8974 13090 9002 13454
rect 9198 13202 9226 15946
rect 9918 15694 10050 15699
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 9918 15661 10050 15666
rect 9918 14910 10050 14915
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 9918 14877 10050 14882
rect 9918 14126 10050 14131
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 9918 14093 10050 14098
rect 10374 13593 10402 18607
rect 10374 13567 10375 13593
rect 10401 13567 10402 13593
rect 9310 13481 9338 13487
rect 9310 13455 9311 13481
rect 9337 13455 9338 13481
rect 9310 13426 9338 13455
rect 9310 13393 9338 13398
rect 10094 13482 10122 13487
rect 9918 13342 10050 13347
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 9918 13309 10050 13314
rect 9702 13258 9730 13263
rect 9926 13258 9954 13263
rect 9702 13211 9730 13230
rect 9758 13257 9954 13258
rect 9758 13231 9927 13257
rect 9953 13231 9954 13257
rect 9758 13230 9954 13231
rect 9198 13155 9226 13174
rect 9478 13202 9506 13207
rect 8974 12810 9002 13062
rect 8974 12777 9002 12782
rect 9142 13145 9170 13151
rect 9142 13119 9143 13145
rect 9169 13119 9170 13145
rect 8022 12727 8023 12753
rect 8049 12727 8050 12753
rect 6846 12697 6874 12703
rect 6846 12671 6847 12697
rect 6873 12671 6874 12697
rect 6846 12530 6874 12671
rect 7350 12698 7378 12703
rect 7350 12651 7378 12670
rect 7854 12698 7882 12703
rect 7854 12697 7994 12698
rect 7854 12671 7855 12697
rect 7881 12671 7994 12697
rect 7854 12670 7994 12671
rect 7854 12665 7882 12670
rect 6902 12642 6930 12647
rect 6902 12641 7042 12642
rect 6902 12615 6903 12641
rect 6929 12615 7042 12641
rect 6902 12614 7042 12615
rect 6902 12609 6930 12614
rect 6846 12497 6874 12502
rect 7014 12417 7042 12614
rect 7574 12641 7602 12647
rect 7574 12615 7575 12641
rect 7601 12615 7602 12641
rect 7574 12530 7602 12615
rect 7742 12642 7770 12647
rect 7742 12641 7826 12642
rect 7742 12615 7743 12641
rect 7769 12615 7826 12641
rect 7742 12614 7826 12615
rect 7742 12609 7770 12614
rect 7742 12530 7770 12535
rect 7462 12502 7658 12530
rect 7014 12391 7015 12417
rect 7041 12391 7042 12417
rect 7014 12385 7042 12391
rect 7406 12418 7434 12423
rect 7406 12362 7434 12390
rect 5950 12305 5978 12334
rect 5950 12279 5951 12305
rect 5977 12279 5978 12305
rect 5950 12273 5978 12279
rect 7350 12361 7434 12362
rect 7350 12335 7407 12361
rect 7433 12335 7434 12361
rect 7350 12334 7434 12335
rect 2238 12166 2370 12171
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2238 12133 2370 12138
rect 2142 11970 2170 11975
rect 2142 11923 2170 11942
rect 5670 11970 5698 11975
rect 5670 11521 5698 11942
rect 7294 11858 7322 11863
rect 7070 11857 7322 11858
rect 7070 11831 7295 11857
rect 7321 11831 7322 11857
rect 7070 11830 7322 11831
rect 5670 11495 5671 11521
rect 5697 11495 5698 11521
rect 5670 11489 5698 11495
rect 6734 11521 6762 11527
rect 6734 11495 6735 11521
rect 6761 11495 6762 11521
rect 2238 11382 2370 11387
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2238 11349 2370 11354
rect 2142 11185 2170 11191
rect 2142 11159 2143 11185
rect 2169 11159 2170 11185
rect 2142 10850 2170 11159
rect 6734 11074 6762 11495
rect 6734 11041 6762 11046
rect 6790 11522 6818 11527
rect 2142 10817 2170 10822
rect 5726 10850 5754 10855
rect 2086 10705 2114 10710
rect 5726 10737 5754 10822
rect 6790 10849 6818 11494
rect 7070 11185 7098 11830
rect 7294 11825 7322 11830
rect 7350 11690 7378 12334
rect 7406 12329 7434 12334
rect 7406 11970 7434 11975
rect 7406 11913 7434 11942
rect 7462 11969 7490 12502
rect 7630 12474 7658 12502
rect 7630 12427 7658 12446
rect 7742 12473 7770 12502
rect 7742 12447 7743 12473
rect 7769 12447 7770 12473
rect 7742 12441 7770 12447
rect 7574 12418 7602 12423
rect 7574 12250 7602 12390
rect 7686 12362 7714 12367
rect 7686 12315 7714 12334
rect 7798 12362 7826 12614
rect 7798 12361 7882 12362
rect 7798 12335 7799 12361
rect 7825 12335 7882 12361
rect 7798 12334 7882 12335
rect 7798 12329 7826 12334
rect 7574 12222 7714 12250
rect 7686 12025 7714 12222
rect 7686 11999 7687 12025
rect 7713 11999 7714 12025
rect 7686 11993 7714 11999
rect 7462 11943 7463 11969
rect 7489 11943 7490 11969
rect 7462 11937 7490 11943
rect 7406 11887 7407 11913
rect 7433 11887 7434 11913
rect 7406 11881 7434 11887
rect 7070 11159 7071 11185
rect 7097 11159 7098 11185
rect 7070 11153 7098 11159
rect 7126 11689 7378 11690
rect 7126 11663 7351 11689
rect 7377 11663 7378 11689
rect 7126 11662 7378 11663
rect 7126 11577 7154 11662
rect 7350 11657 7378 11662
rect 7126 11551 7127 11577
rect 7153 11551 7154 11577
rect 6790 10823 6791 10849
rect 6817 10823 6818 10849
rect 6790 10817 6818 10823
rect 7126 10794 7154 11551
rect 7518 11577 7546 11583
rect 7518 11551 7519 11577
rect 7545 11551 7546 11577
rect 7294 11186 7322 11191
rect 7294 11139 7322 11158
rect 7350 11074 7378 11079
rect 7350 11027 7378 11046
rect 7406 11073 7434 11079
rect 7406 11047 7407 11073
rect 7433 11047 7434 11073
rect 7126 10793 7322 10794
rect 7126 10767 7127 10793
rect 7153 10767 7322 10793
rect 7126 10766 7322 10767
rect 7126 10761 7154 10766
rect 5726 10711 5727 10737
rect 5753 10711 5754 10737
rect 5726 10705 5754 10711
rect 2238 10598 2370 10603
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2238 10565 2370 10570
rect 6566 10458 6594 10463
rect 4998 10010 5026 10015
rect 2238 9814 2370 9819
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2238 9781 2370 9786
rect 966 9673 994 9679
rect 966 9647 967 9673
rect 993 9647 994 9673
rect 966 9450 994 9647
rect 4998 9674 5026 9982
rect 4998 9627 5026 9646
rect 6566 9953 6594 10430
rect 7294 10458 7322 10766
rect 7406 10682 7434 11047
rect 7462 10850 7490 10855
rect 7462 10803 7490 10822
rect 7518 10737 7546 11551
rect 7630 11577 7658 11583
rect 7742 11578 7770 11583
rect 7630 11551 7631 11577
rect 7657 11551 7658 11577
rect 7574 11522 7602 11527
rect 7574 11475 7602 11494
rect 7630 11185 7658 11551
rect 7630 11159 7631 11185
rect 7657 11159 7658 11185
rect 7630 11153 7658 11159
rect 7686 11577 7770 11578
rect 7686 11551 7743 11577
rect 7769 11551 7770 11577
rect 7686 11550 7770 11551
rect 7518 10711 7519 10737
rect 7545 10711 7546 10737
rect 7518 10705 7546 10711
rect 7574 10793 7602 10799
rect 7574 10767 7575 10793
rect 7601 10767 7602 10793
rect 7406 10649 7434 10654
rect 7294 10411 7322 10430
rect 7574 10122 7602 10767
rect 7686 10626 7714 11550
rect 7742 11545 7770 11550
rect 7798 11130 7826 11135
rect 7854 11130 7882 12334
rect 7910 12361 7938 12367
rect 7910 12335 7911 12361
rect 7937 12335 7938 12361
rect 7910 11690 7938 12335
rect 7910 11657 7938 11662
rect 7966 11634 7994 12670
rect 8022 12418 8050 12727
rect 8414 12698 8442 12703
rect 8414 12697 9058 12698
rect 8414 12671 8415 12697
rect 8441 12671 9058 12697
rect 8414 12670 9058 12671
rect 8414 12665 8442 12670
rect 9030 12473 9058 12670
rect 9030 12447 9031 12473
rect 9057 12447 9058 12473
rect 9030 12441 9058 12447
rect 9142 12474 9170 13119
rect 9142 12441 9170 12446
rect 9310 13145 9338 13151
rect 9310 13119 9311 13145
rect 9337 13119 9338 13145
rect 8022 12385 8050 12390
rect 8974 12362 9002 12367
rect 8918 12361 9002 12362
rect 8918 12335 8975 12361
rect 9001 12335 9002 12361
rect 8918 12334 9002 12335
rect 8918 11689 8946 12334
rect 8974 12329 9002 12334
rect 9086 12362 9114 12367
rect 9086 12315 9114 12334
rect 9310 12361 9338 13119
rect 9478 12809 9506 13174
rect 9478 12783 9479 12809
rect 9505 12783 9506 12809
rect 9478 12777 9506 12783
rect 9646 13146 9674 13151
rect 9758 13146 9786 13230
rect 9926 13225 9954 13230
rect 10094 13257 10122 13454
rect 10094 13231 10095 13257
rect 10121 13231 10122 13257
rect 10094 13225 10122 13231
rect 10150 13426 10178 13431
rect 9646 13145 9786 13146
rect 9646 13119 9647 13145
rect 9673 13119 9786 13145
rect 9646 13118 9786 13119
rect 9814 13145 9842 13151
rect 9814 13119 9815 13145
rect 9841 13119 9842 13145
rect 9310 12335 9311 12361
rect 9337 12335 9338 12361
rect 9310 12329 9338 12335
rect 9366 12642 9394 12647
rect 8918 11663 8919 11689
rect 8945 11663 8946 11689
rect 8918 11657 8946 11663
rect 7966 11186 7994 11606
rect 8862 11634 8890 11639
rect 8862 11587 8890 11606
rect 8694 11578 8722 11583
rect 7966 11185 8274 11186
rect 7966 11159 7967 11185
rect 7993 11159 8274 11185
rect 7966 11158 8274 11159
rect 7966 11153 7994 11158
rect 7826 11102 7882 11130
rect 7798 11083 7826 11102
rect 7742 11074 7770 11079
rect 7742 11027 7770 11046
rect 7966 11074 7994 11079
rect 7966 10850 7994 11046
rect 8246 10905 8274 11158
rect 8638 11185 8666 11191
rect 8638 11159 8639 11185
rect 8665 11159 8666 11185
rect 8638 11130 8666 11159
rect 8638 11097 8666 11102
rect 8694 11129 8722 11550
rect 9030 11578 9058 11583
rect 9030 11531 9058 11550
rect 9030 11242 9058 11247
rect 9030 11241 9114 11242
rect 9030 11215 9031 11241
rect 9057 11215 9114 11241
rect 9030 11214 9114 11215
rect 9030 11209 9058 11214
rect 8694 11103 8695 11129
rect 8721 11103 8722 11129
rect 8246 10879 8247 10905
rect 8273 10879 8274 10905
rect 8246 10873 8274 10879
rect 8302 10906 8330 10911
rect 8694 10906 8722 11103
rect 8862 11186 8890 11191
rect 8750 10906 8778 10911
rect 7910 10849 7994 10850
rect 7910 10823 7967 10849
rect 7993 10823 7994 10849
rect 7910 10822 7994 10823
rect 7742 10794 7770 10799
rect 7742 10682 7770 10766
rect 7742 10649 7770 10654
rect 7686 10593 7714 10598
rect 7854 10570 7882 10575
rect 7630 10458 7658 10463
rect 7630 10411 7658 10430
rect 7574 10089 7602 10094
rect 7070 10066 7098 10071
rect 7014 10038 7070 10066
rect 6902 10010 6930 10015
rect 6566 9927 6567 9953
rect 6593 9927 6594 9953
rect 2142 9618 2170 9623
rect 2142 9571 2170 9590
rect 6398 9618 6426 9623
rect 6566 9618 6594 9927
rect 6398 9617 6594 9618
rect 6398 9591 6399 9617
rect 6425 9591 6594 9617
rect 6398 9590 6594 9591
rect 6846 10009 6930 10010
rect 6846 9983 6903 10009
rect 6929 9983 6930 10009
rect 6846 9982 6930 9983
rect 6062 9561 6090 9567
rect 6062 9535 6063 9561
rect 6089 9535 6090 9561
rect 6062 9506 6090 9535
rect 6062 9473 6090 9478
rect 966 9417 994 9422
rect 5054 9226 5082 9231
rect 5054 9179 5082 9198
rect 6398 9226 6426 9590
rect 6846 9394 6874 9982
rect 6902 9977 6930 9982
rect 6958 9618 6986 9623
rect 7014 9618 7042 10038
rect 7070 10019 7098 10038
rect 7406 10066 7434 10071
rect 7742 10066 7770 10071
rect 7434 10038 7546 10066
rect 7406 10019 7434 10038
rect 7238 10010 7266 10015
rect 7238 9963 7266 9982
rect 7238 9898 7266 9903
rect 7070 9897 7266 9898
rect 7070 9871 7239 9897
rect 7265 9871 7266 9897
rect 7070 9870 7266 9871
rect 7070 9729 7098 9870
rect 7238 9865 7266 9870
rect 7070 9703 7071 9729
rect 7097 9703 7098 9729
rect 7070 9697 7098 9703
rect 7294 9786 7322 9791
rect 7126 9618 7154 9623
rect 7014 9617 7154 9618
rect 7014 9591 7127 9617
rect 7153 9591 7154 9617
rect 7014 9590 7154 9591
rect 6958 9571 6986 9590
rect 7126 9585 7154 9590
rect 7294 9617 7322 9758
rect 7294 9591 7295 9617
rect 7321 9591 7322 9617
rect 7294 9585 7322 9591
rect 6902 9506 6930 9511
rect 6902 9459 6930 9478
rect 7462 9505 7490 9511
rect 7462 9479 7463 9505
rect 7489 9479 7490 9505
rect 7462 9394 7490 9479
rect 6846 9366 7490 9394
rect 6790 9338 6818 9343
rect 6846 9338 6874 9366
rect 6790 9337 6874 9338
rect 6790 9311 6791 9337
rect 6817 9311 6874 9337
rect 6790 9310 6874 9311
rect 7518 9337 7546 10038
rect 7742 10019 7770 10038
rect 7686 10009 7714 10015
rect 7686 9983 7687 10009
rect 7713 9983 7714 10009
rect 7574 9730 7602 9735
rect 7686 9730 7714 9983
rect 7742 9898 7770 9903
rect 7742 9851 7770 9870
rect 7602 9702 7714 9730
rect 7574 9394 7602 9702
rect 7742 9674 7770 9679
rect 7686 9618 7714 9623
rect 7630 9562 7658 9567
rect 7630 9515 7658 9534
rect 7630 9394 7658 9399
rect 7574 9366 7630 9394
rect 7630 9361 7658 9366
rect 7518 9311 7519 9337
rect 7545 9311 7546 9337
rect 6790 9305 6818 9310
rect 7518 9305 7546 9311
rect 7126 9281 7154 9287
rect 7126 9255 7127 9281
rect 7153 9255 7154 9281
rect 6734 9226 6762 9231
rect 6958 9226 6986 9231
rect 5390 9170 5418 9175
rect 5390 9123 5418 9142
rect 2238 9030 2370 9035
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2238 8997 2370 9002
rect 6398 8722 6426 9198
rect 6454 9225 6986 9226
rect 6454 9199 6735 9225
rect 6761 9199 6959 9225
rect 6985 9199 6986 9225
rect 6454 9198 6986 9199
rect 6454 9169 6482 9198
rect 6734 9193 6762 9198
rect 6958 9193 6986 9198
rect 6454 9143 6455 9169
rect 6481 9143 6482 9169
rect 6454 9137 6482 9143
rect 7126 9114 7154 9255
rect 7630 9282 7658 9287
rect 7406 9226 7434 9231
rect 7126 9081 7154 9086
rect 7182 9225 7434 9226
rect 7182 9199 7407 9225
rect 7433 9199 7434 9225
rect 7182 9198 7434 9199
rect 7126 8946 7154 8951
rect 7182 8946 7210 9198
rect 7406 9193 7434 9198
rect 6790 8945 7210 8946
rect 6790 8919 7127 8945
rect 7153 8919 7210 8945
rect 6790 8918 7210 8919
rect 7462 9169 7490 9175
rect 7462 9143 7463 9169
rect 7489 9143 7490 9169
rect 7462 8946 7490 9143
rect 6790 8833 6818 8918
rect 7126 8913 7154 8918
rect 7462 8913 7490 8918
rect 7630 8889 7658 9254
rect 7686 9225 7714 9590
rect 7686 9199 7687 9225
rect 7713 9199 7714 9225
rect 7686 9193 7714 9199
rect 7630 8863 7631 8889
rect 7657 8863 7658 8889
rect 7630 8857 7658 8863
rect 7686 8890 7714 8895
rect 6790 8807 6791 8833
rect 6817 8807 6818 8833
rect 6790 8801 6818 8807
rect 6902 8806 7098 8834
rect 6846 8778 6874 8783
rect 6902 8778 6930 8806
rect 6846 8777 6930 8778
rect 6846 8751 6847 8777
rect 6873 8751 6930 8777
rect 6846 8750 6930 8751
rect 6846 8745 6874 8750
rect 6454 8722 6482 8727
rect 6398 8694 6454 8722
rect 6454 8675 6482 8694
rect 6790 8722 6818 8727
rect 2238 8246 2370 8251
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2238 8213 2370 8218
rect 5950 7714 5978 7719
rect 5950 7667 5978 7686
rect 5614 7657 5642 7663
rect 5614 7631 5615 7657
rect 5641 7631 5642 7657
rect 5614 7602 5642 7631
rect 5614 7569 5642 7574
rect 6790 7602 6818 8694
rect 2238 7462 2370 7467
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2238 7429 2370 7434
rect 6790 7265 6818 7574
rect 6790 7239 6791 7265
rect 6817 7239 6818 7265
rect 6790 7098 6818 7239
rect 6958 8721 6986 8727
rect 6958 8695 6959 8721
rect 6985 8695 6986 8721
rect 6958 8498 6986 8695
rect 7070 8610 7098 8806
rect 7126 8778 7154 8783
rect 7126 8731 7154 8750
rect 7182 8777 7210 8783
rect 7182 8751 7183 8777
rect 7209 8751 7210 8777
rect 7182 8722 7210 8751
rect 7182 8689 7210 8694
rect 7350 8721 7378 8727
rect 7350 8695 7351 8721
rect 7377 8695 7378 8721
rect 7350 8610 7378 8695
rect 7070 8582 7378 8610
rect 7238 8553 7266 8582
rect 7238 8527 7239 8553
rect 7265 8527 7266 8553
rect 7238 8521 7266 8527
rect 7350 8498 7378 8503
rect 6958 7266 6986 8470
rect 7294 8497 7378 8498
rect 7294 8471 7351 8497
rect 7377 8471 7378 8497
rect 7294 8470 7378 8471
rect 7294 8050 7322 8470
rect 7350 8465 7378 8470
rect 7406 8442 7434 8447
rect 7406 8395 7434 8414
rect 7630 8442 7658 8447
rect 7630 8395 7658 8414
rect 7686 8161 7714 8862
rect 7742 8834 7770 9646
rect 7854 9506 7882 10542
rect 7910 9674 7938 10822
rect 7966 10817 7994 10822
rect 8022 10850 8050 10855
rect 8022 10849 8218 10850
rect 8022 10823 8023 10849
rect 8049 10823 8218 10849
rect 8022 10822 8218 10823
rect 8022 10817 8050 10822
rect 8022 10682 8050 10687
rect 8022 10635 8050 10654
rect 8078 10122 8106 10127
rect 8022 10066 8050 10071
rect 8022 10019 8050 10038
rect 7966 10010 7994 10015
rect 7966 9963 7994 9982
rect 8022 9898 8050 9903
rect 8078 9898 8106 10094
rect 7910 9627 7938 9646
rect 7966 9897 8106 9898
rect 7966 9871 8023 9897
rect 8049 9871 8106 9897
rect 7966 9870 8106 9871
rect 7910 9506 7938 9511
rect 7854 9505 7938 9506
rect 7854 9479 7911 9505
rect 7937 9479 7938 9505
rect 7854 9478 7938 9479
rect 7910 9473 7938 9478
rect 7910 9394 7938 9399
rect 7910 9337 7938 9366
rect 7910 9311 7911 9337
rect 7937 9311 7938 9337
rect 7910 9305 7938 9311
rect 7966 9114 7994 9870
rect 8022 9865 8050 9870
rect 8022 9617 8050 9623
rect 8022 9591 8023 9617
rect 8049 9591 8050 9617
rect 8022 9338 8050 9591
rect 8190 9394 8218 10822
rect 8302 10121 8330 10878
rect 8582 10905 8778 10906
rect 8582 10879 8751 10905
rect 8777 10879 8778 10905
rect 8582 10878 8778 10879
rect 8358 10793 8386 10799
rect 8358 10767 8359 10793
rect 8385 10767 8386 10793
rect 8358 10570 8386 10767
rect 8358 10537 8386 10542
rect 8302 10095 8303 10121
rect 8329 10095 8330 10121
rect 8302 10089 8330 10095
rect 8246 10010 8274 10015
rect 8414 10010 8442 10015
rect 8246 9897 8274 9982
rect 8246 9871 8247 9897
rect 8273 9871 8274 9897
rect 8246 9562 8274 9871
rect 8358 10009 8442 10010
rect 8358 9983 8415 10009
rect 8441 9983 8442 10009
rect 8358 9982 8442 9983
rect 8358 9618 8386 9982
rect 8414 9977 8442 9982
rect 8358 9585 8386 9590
rect 8470 9842 8498 9847
rect 8246 9529 8274 9534
rect 8190 9366 8330 9394
rect 8022 9310 8274 9338
rect 8022 9281 8050 9310
rect 8022 9255 8023 9281
rect 8049 9255 8050 9281
rect 8022 9249 8050 9255
rect 7966 9081 7994 9086
rect 8078 9226 8106 9231
rect 8078 9002 8106 9198
rect 8022 8946 8050 8951
rect 8078 8946 8106 8974
rect 8022 8945 8106 8946
rect 8022 8919 8023 8945
rect 8049 8919 8106 8945
rect 8022 8918 8106 8919
rect 8190 9226 8218 9231
rect 8022 8913 8050 8918
rect 8190 8889 8218 9198
rect 8190 8863 8191 8889
rect 8217 8863 8218 8889
rect 7742 8553 7770 8806
rect 8134 8833 8162 8839
rect 8134 8807 8135 8833
rect 8161 8807 8162 8833
rect 7742 8527 7743 8553
rect 7769 8527 7770 8553
rect 7742 8521 7770 8527
rect 7910 8722 7938 8727
rect 7910 8498 7938 8694
rect 7910 8451 7938 8470
rect 7686 8135 7687 8161
rect 7713 8135 7714 8161
rect 7630 8106 7658 8111
rect 7014 8049 7322 8050
rect 7014 8023 7295 8049
rect 7321 8023 7322 8049
rect 7014 8022 7322 8023
rect 7014 7601 7042 8022
rect 7294 8017 7322 8022
rect 7462 8078 7630 8106
rect 7462 7993 7490 8078
rect 7630 8059 7658 8078
rect 7462 7967 7463 7993
rect 7489 7967 7490 7993
rect 7462 7961 7490 7967
rect 7686 7714 7714 8135
rect 7854 8442 7882 8447
rect 8078 8442 8106 8447
rect 7854 8161 7882 8414
rect 7854 8135 7855 8161
rect 7881 8135 7882 8161
rect 7854 8129 7882 8135
rect 7966 8414 8078 8442
rect 7910 8106 7938 8111
rect 7966 8106 7994 8414
rect 8078 8395 8106 8414
rect 8134 8386 8162 8807
rect 8190 8498 8218 8863
rect 8190 8465 8218 8470
rect 8246 8553 8274 9310
rect 8302 8890 8330 9366
rect 8470 9282 8498 9814
rect 8582 9506 8610 10878
rect 8750 10873 8778 10878
rect 8806 10793 8834 10799
rect 8806 10767 8807 10793
rect 8833 10767 8834 10793
rect 8806 10122 8834 10767
rect 8806 10089 8834 10094
rect 8862 10737 8890 11158
rect 8862 10711 8863 10737
rect 8889 10711 8890 10737
rect 8750 10066 8778 10071
rect 8694 10038 8750 10066
rect 8638 10010 8666 10015
rect 8638 9617 8666 9982
rect 8638 9591 8639 9617
rect 8665 9591 8666 9617
rect 8638 9585 8666 9591
rect 8638 9506 8666 9511
rect 8582 9478 8638 9506
rect 8638 9473 8666 9478
rect 8694 9282 8722 10038
rect 8750 10033 8778 10038
rect 8862 9842 8890 10711
rect 8974 11129 9002 11135
rect 8974 11103 8975 11129
rect 9001 11103 9002 11129
rect 8974 10458 9002 11103
rect 8862 9809 8890 9814
rect 8918 10430 9002 10458
rect 8750 9617 8778 9623
rect 8750 9591 8751 9617
rect 8777 9591 8778 9617
rect 8750 9562 8778 9591
rect 8750 9529 8778 9534
rect 8806 9562 8834 9567
rect 8918 9562 8946 10430
rect 8806 9561 8946 9562
rect 8806 9535 8807 9561
rect 8833 9535 8946 9561
rect 8806 9534 8946 9535
rect 8974 10290 9002 10295
rect 8806 9338 8834 9534
rect 8806 9305 8834 9310
rect 8918 9338 8946 9343
rect 8974 9338 9002 10262
rect 9030 10010 9058 10015
rect 9030 9963 9058 9982
rect 9030 9562 9058 9567
rect 9030 9515 9058 9534
rect 9086 9338 9114 11214
rect 9254 11130 9282 11135
rect 9254 11083 9282 11102
rect 9366 10850 9394 12614
rect 9422 12474 9450 12479
rect 9422 12427 9450 12446
rect 9534 12362 9562 12367
rect 9646 12362 9674 13118
rect 9814 12753 9842 13119
rect 10094 12866 10122 12871
rect 10150 12866 10178 13398
rect 10318 13426 10346 13431
rect 10318 13145 10346 13398
rect 10374 13258 10402 13567
rect 10654 13481 10682 18999
rect 12278 19025 12306 19031
rect 12278 18999 12279 19025
rect 12305 18999 12306 19025
rect 10710 18746 10738 18751
rect 10710 18699 10738 18718
rect 11718 14154 11746 14159
rect 11662 14126 11718 14154
rect 11158 13594 11186 13599
rect 10654 13455 10655 13481
rect 10681 13455 10682 13481
rect 10654 13449 10682 13455
rect 10766 13537 10794 13543
rect 10766 13511 10767 13537
rect 10793 13511 10794 13537
rect 10374 13225 10402 13230
rect 10766 13258 10794 13511
rect 11102 13538 11130 13543
rect 11102 13481 11130 13510
rect 11102 13455 11103 13481
rect 11129 13455 11130 13481
rect 11102 13449 11130 13455
rect 11158 13482 11186 13566
rect 11158 13435 11186 13454
rect 11382 13537 11410 13543
rect 11382 13511 11383 13537
rect 11409 13511 11410 13537
rect 11382 13482 11410 13511
rect 11382 13449 11410 13454
rect 11662 13538 11690 14126
rect 11718 14121 11746 14126
rect 12278 14154 12306 18999
rect 13398 18745 13426 19278
rect 17598 19222 17730 19227
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17598 19189 17730 19194
rect 13398 18719 13399 18745
rect 13425 18719 13426 18745
rect 13398 18713 13426 18719
rect 20118 18689 20146 18695
rect 20118 18663 20119 18689
rect 20145 18663 20146 18689
rect 12278 14121 12306 14126
rect 13006 18633 13034 18639
rect 13006 18607 13007 18633
rect 13033 18607 13034 18633
rect 13006 13986 13034 18607
rect 20118 18522 20146 18663
rect 20118 18489 20146 18494
rect 17598 18438 17730 18443
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17598 18405 17730 18410
rect 17598 17654 17730 17659
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17598 17621 17730 17626
rect 20118 17345 20146 17351
rect 20118 17319 20119 17345
rect 20145 17319 20146 17345
rect 20118 17178 20146 17319
rect 20118 17145 20146 17150
rect 17598 16870 17730 16875
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17598 16837 17730 16842
rect 17598 16086 17730 16091
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17598 16053 17730 16058
rect 17598 15302 17730 15307
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17598 15269 17730 15274
rect 17598 14518 17730 14523
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17598 14485 17730 14490
rect 12782 13958 13034 13986
rect 12782 13593 12810 13958
rect 12782 13567 12783 13593
rect 12809 13567 12810 13593
rect 12782 13561 12810 13567
rect 12950 13873 12978 13879
rect 12950 13847 12951 13873
rect 12977 13847 12978 13873
rect 10766 13225 10794 13230
rect 10990 13425 11018 13431
rect 10990 13399 10991 13425
rect 11017 13399 11018 13425
rect 10318 13119 10319 13145
rect 10345 13119 10346 13145
rect 10318 13113 10346 13119
rect 10654 13090 10682 13095
rect 10654 13089 10906 13090
rect 10654 13063 10655 13089
rect 10681 13063 10906 13089
rect 10654 13062 10906 13063
rect 10654 13057 10682 13062
rect 10094 12865 10178 12866
rect 10094 12839 10095 12865
rect 10121 12839 10178 12865
rect 10094 12838 10178 12839
rect 10094 12833 10122 12838
rect 10374 12810 10402 12815
rect 10374 12763 10402 12782
rect 9814 12727 9815 12753
rect 9841 12727 9842 12753
rect 9814 12721 9842 12727
rect 10150 12754 10178 12759
rect 10150 12707 10178 12726
rect 10318 12754 10346 12759
rect 9926 12642 9954 12647
rect 9534 12361 9674 12362
rect 9534 12335 9535 12361
rect 9561 12335 9674 12361
rect 9534 12334 9674 12335
rect 9758 12641 9954 12642
rect 9758 12615 9927 12641
rect 9953 12615 9954 12641
rect 9758 12614 9954 12615
rect 9366 10817 9394 10822
rect 9422 11073 9450 11079
rect 9422 11047 9423 11073
rect 9449 11047 9450 11073
rect 9422 10794 9450 11047
rect 9534 10906 9562 12334
rect 9758 11969 9786 12614
rect 9926 12609 9954 12614
rect 10038 12642 10066 12661
rect 10038 12609 10066 12614
rect 9918 12558 10050 12563
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 9918 12525 10050 12530
rect 9814 12362 9842 12367
rect 9814 12315 9842 12334
rect 9758 11943 9759 11969
rect 9785 11943 9786 11969
rect 9758 11937 9786 11943
rect 9590 11913 9618 11919
rect 9590 11887 9591 11913
rect 9617 11887 9618 11913
rect 9590 11634 9618 11887
rect 9590 11601 9618 11606
rect 9646 11857 9674 11863
rect 9646 11831 9647 11857
rect 9673 11831 9674 11857
rect 9646 11354 9674 11831
rect 9918 11774 10050 11779
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 9918 11741 10050 11746
rect 10206 11690 10234 11695
rect 10318 11690 10346 12726
rect 10878 12753 10906 13062
rect 10878 12727 10879 12753
rect 10905 12727 10906 12753
rect 10878 12721 10906 12727
rect 10990 12754 11018 13399
rect 11662 13090 11690 13510
rect 11998 13538 12026 13543
rect 11718 13481 11746 13487
rect 11718 13455 11719 13481
rect 11745 13455 11746 13481
rect 11718 13454 11746 13455
rect 11718 13426 11858 13454
rect 11830 13257 11858 13426
rect 11830 13231 11831 13257
rect 11857 13231 11858 13257
rect 11830 13225 11858 13231
rect 11942 13201 11970 13207
rect 11942 13175 11943 13201
rect 11969 13175 11970 13201
rect 11718 13090 11746 13095
rect 11662 13089 11746 13090
rect 11662 13063 11719 13089
rect 11745 13063 11746 13089
rect 11662 13062 11746 13063
rect 11718 13057 11746 13062
rect 11046 12754 11074 12759
rect 10990 12753 11074 12754
rect 10990 12727 11047 12753
rect 11073 12727 11074 12753
rect 10990 12726 11074 12727
rect 11046 12721 11074 12726
rect 11942 12754 11970 13175
rect 11998 13201 12026 13510
rect 12894 13538 12922 13543
rect 12894 13491 12922 13510
rect 11998 13175 11999 13201
rect 12025 13175 12026 13201
rect 11998 13169 12026 13175
rect 12222 13482 12250 13487
rect 12950 13454 12978 13847
rect 12222 13089 12250 13454
rect 12222 13063 12223 13089
rect 12249 13063 12250 13089
rect 11942 12721 11970 12726
rect 12110 12754 12138 12759
rect 12222 12754 12250 13063
rect 12110 12753 12250 12754
rect 12110 12727 12111 12753
rect 12137 12727 12250 12753
rect 12110 12726 12250 12727
rect 12726 13426 12978 13454
rect 13006 13481 13034 13958
rect 18942 13929 18970 13935
rect 18942 13903 18943 13929
rect 18969 13903 18970 13929
rect 17598 13734 17730 13739
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17598 13701 17730 13706
rect 13006 13455 13007 13481
rect 13033 13455 13034 13481
rect 13006 13449 13034 13455
rect 13062 13594 13090 13599
rect 13062 13481 13090 13566
rect 13342 13594 13370 13599
rect 13342 13537 13370 13566
rect 13342 13511 13343 13537
rect 13369 13511 13370 13537
rect 13342 13505 13370 13511
rect 18830 13537 18858 13543
rect 18830 13511 18831 13537
rect 18857 13511 18858 13537
rect 13062 13455 13063 13481
rect 13089 13455 13090 13481
rect 13062 13454 13090 13455
rect 13398 13482 13426 13487
rect 13062 13426 13146 13454
rect 13398 13435 13426 13454
rect 14630 13482 14658 13487
rect 12726 13089 12754 13426
rect 12950 13201 12978 13207
rect 12950 13175 12951 13201
rect 12977 13175 12978 13201
rect 12838 13146 12866 13151
rect 12726 13063 12727 13089
rect 12753 13063 12754 13089
rect 10990 12642 11018 12647
rect 10990 12595 11018 12614
rect 12110 12642 12138 12726
rect 12446 12698 12474 12703
rect 12446 12697 12586 12698
rect 12446 12671 12447 12697
rect 12473 12671 12586 12697
rect 12446 12670 12586 12671
rect 12446 12665 12474 12670
rect 12110 12609 12138 12614
rect 12558 12473 12586 12670
rect 12726 12642 12754 13063
rect 12726 12609 12754 12614
rect 12782 13145 12866 13146
rect 12782 13119 12839 13145
rect 12865 13119 12866 13145
rect 12782 13118 12866 13119
rect 12558 12447 12559 12473
rect 12585 12447 12586 12473
rect 12558 12441 12586 12447
rect 12670 12417 12698 12423
rect 12670 12391 12671 12417
rect 12697 12391 12698 12417
rect 12390 12362 12418 12367
rect 12390 12026 12418 12334
rect 12390 12025 12586 12026
rect 12390 11999 12391 12025
rect 12417 11999 12586 12025
rect 12390 11998 12586 11999
rect 12390 11993 12418 11998
rect 10206 11643 10234 11662
rect 10262 11689 10346 11690
rect 10262 11663 10319 11689
rect 10345 11663 10346 11689
rect 10262 11662 10346 11663
rect 10150 11577 10178 11583
rect 10150 11551 10151 11577
rect 10177 11551 10178 11577
rect 9646 11321 9674 11326
rect 9870 11521 9898 11527
rect 9870 11495 9871 11521
rect 9897 11495 9898 11521
rect 9870 11242 9898 11495
rect 10150 11522 10178 11551
rect 10150 11494 10234 11522
rect 9926 11466 9954 11471
rect 9926 11465 10178 11466
rect 9926 11439 9927 11465
rect 9953 11439 10178 11465
rect 9926 11438 10178 11439
rect 9926 11433 9954 11438
rect 10038 11354 10066 11359
rect 10066 11326 10122 11354
rect 10038 11321 10066 11326
rect 9534 10873 9562 10878
rect 9646 11214 9898 11242
rect 9534 10794 9562 10799
rect 9646 10794 9674 11214
rect 9926 11186 9954 11191
rect 9870 11185 9954 11186
rect 9870 11159 9927 11185
rect 9953 11159 9954 11185
rect 9870 11158 9954 11159
rect 9814 11129 9842 11135
rect 9814 11103 9815 11129
rect 9841 11103 9842 11129
rect 9422 10793 9674 10794
rect 9422 10767 9535 10793
rect 9561 10767 9674 10793
rect 9422 10766 9674 10767
rect 9702 10906 9730 10911
rect 9814 10906 9842 11103
rect 9870 11074 9898 11158
rect 9926 11153 9954 11158
rect 9870 11041 9898 11046
rect 9918 10990 10050 10995
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 9918 10957 10050 10962
rect 9814 10878 9898 10906
rect 9702 10849 9730 10878
rect 9702 10823 9703 10849
rect 9729 10823 9730 10849
rect 9310 10738 9338 10743
rect 9198 10066 9226 10071
rect 9198 10009 9226 10038
rect 9198 9983 9199 10009
rect 9225 9983 9226 10009
rect 9198 9977 9226 9983
rect 9310 10010 9338 10710
rect 9422 10010 9450 10015
rect 9310 10009 9450 10010
rect 9310 9983 9423 10009
rect 9449 9983 9450 10009
rect 9310 9982 9450 9983
rect 9422 9977 9450 9982
rect 8918 9337 9002 9338
rect 8918 9311 8919 9337
rect 8945 9311 9002 9337
rect 8918 9310 9002 9311
rect 9030 9310 9114 9338
rect 9142 9898 9170 9903
rect 8470 9249 8498 9254
rect 8638 9281 8722 9282
rect 8638 9255 8695 9281
rect 8721 9255 8722 9281
rect 8638 9254 8722 9255
rect 8638 9058 8666 9254
rect 8694 9249 8722 9254
rect 8806 9226 8834 9231
rect 8806 9179 8834 9198
rect 8638 9025 8666 9030
rect 8694 9114 8722 9119
rect 8694 8945 8722 9086
rect 8694 8919 8695 8945
rect 8721 8919 8722 8945
rect 8694 8913 8722 8919
rect 8302 8857 8330 8862
rect 8526 8834 8554 8839
rect 8526 8787 8554 8806
rect 8246 8527 8247 8553
rect 8273 8527 8274 8553
rect 8190 8386 8218 8391
rect 8134 8358 8190 8386
rect 8190 8353 8218 8358
rect 7910 8105 7994 8106
rect 7910 8079 7911 8105
rect 7937 8079 7994 8105
rect 7910 8078 7994 8079
rect 7910 8073 7938 8078
rect 7686 7681 7714 7686
rect 7014 7575 7015 7601
rect 7041 7575 7042 7601
rect 7014 7569 7042 7575
rect 7238 7601 7266 7607
rect 7238 7575 7239 7601
rect 7265 7575 7266 7601
rect 6958 7238 7154 7266
rect 7126 7209 7154 7238
rect 7126 7183 7127 7209
rect 7153 7183 7154 7209
rect 7126 7177 7154 7183
rect 7238 7154 7266 7575
rect 7966 7574 7994 8078
rect 8246 8106 8274 8527
rect 8638 8721 8666 8727
rect 8638 8695 8639 8721
rect 8665 8695 8666 8721
rect 8414 8497 8442 8503
rect 8414 8471 8415 8497
rect 8441 8471 8442 8497
rect 8414 8386 8442 8471
rect 8414 8353 8442 8358
rect 8246 8073 8274 8078
rect 7966 7546 8218 7574
rect 8190 7321 8218 7546
rect 8190 7295 8191 7321
rect 8217 7295 8218 7321
rect 8190 7289 8218 7295
rect 8638 7266 8666 8695
rect 8862 8442 8890 8447
rect 8862 8395 8890 8414
rect 8918 8386 8946 9310
rect 8974 9226 9002 9231
rect 8974 9179 9002 9198
rect 8918 8353 8946 8358
rect 8638 7233 8666 7238
rect 7406 7154 7434 7159
rect 7182 7126 7406 7154
rect 7182 7098 7210 7126
rect 7406 7121 7434 7126
rect 7742 7154 7770 7159
rect 6790 7070 7210 7098
rect 2238 6678 2370 6683
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2238 6645 2370 6650
rect 7742 6481 7770 7126
rect 8414 7154 8442 7159
rect 8414 7107 8442 7126
rect 8974 7154 9002 7159
rect 8246 6930 8274 6935
rect 8078 6929 8274 6930
rect 8078 6903 8247 6929
rect 8273 6903 8274 6929
rect 8078 6902 8274 6903
rect 8078 6537 8106 6902
rect 8246 6897 8274 6902
rect 8414 6874 8442 6879
rect 8414 6827 8442 6846
rect 8750 6874 8778 6879
rect 8750 6827 8778 6846
rect 8918 6874 8946 6879
rect 8918 6827 8946 6846
rect 8974 6818 9002 7126
rect 9030 6873 9058 9310
rect 9086 9226 9114 9231
rect 9086 8833 9114 9198
rect 9086 8807 9087 8833
rect 9113 8807 9114 8833
rect 9086 8801 9114 8807
rect 9142 8777 9170 9870
rect 9198 9898 9226 9903
rect 9534 9898 9562 10766
rect 9702 10122 9730 10823
rect 9870 10794 9898 10878
rect 10038 10905 10066 10911
rect 10038 10879 10039 10905
rect 10065 10879 10066 10905
rect 9870 10761 9898 10766
rect 9926 10849 9954 10855
rect 9926 10823 9927 10849
rect 9953 10823 9954 10849
rect 9926 10290 9954 10823
rect 10038 10850 10066 10879
rect 10038 10817 10066 10822
rect 10038 10402 10066 10407
rect 10038 10355 10066 10374
rect 9926 10257 9954 10262
rect 9918 10206 10050 10211
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 9918 10173 10050 10178
rect 9702 10089 9730 10094
rect 9702 10010 9730 10015
rect 9730 9982 9786 10010
rect 9702 9977 9730 9982
rect 9198 9897 9562 9898
rect 9198 9871 9199 9897
rect 9225 9871 9562 9897
rect 9198 9870 9562 9871
rect 9198 9282 9226 9870
rect 9254 9730 9282 9735
rect 9254 9617 9282 9702
rect 9254 9591 9255 9617
rect 9281 9591 9282 9617
rect 9254 9394 9282 9591
rect 9422 9618 9450 9623
rect 9422 9571 9450 9590
rect 9702 9618 9730 9623
rect 9702 9561 9730 9590
rect 9702 9535 9703 9561
rect 9729 9535 9730 9561
rect 9702 9529 9730 9535
rect 9254 9361 9282 9366
rect 9478 9505 9506 9511
rect 9478 9479 9479 9505
rect 9505 9479 9506 9505
rect 9254 9282 9282 9287
rect 9198 9254 9254 9282
rect 9254 9249 9282 9254
rect 9422 9225 9450 9231
rect 9422 9199 9423 9225
rect 9449 9199 9450 9225
rect 9310 9170 9338 9175
rect 9310 9123 9338 9142
rect 9422 9170 9450 9199
rect 9422 9137 9450 9142
rect 9142 8751 9143 8777
rect 9169 8751 9170 8777
rect 9142 8745 9170 8751
rect 9198 9114 9226 9119
rect 9142 8442 9170 8447
rect 9198 8442 9226 9086
rect 9254 9113 9282 9119
rect 9254 9087 9255 9113
rect 9281 9087 9282 9113
rect 9254 8834 9282 9087
rect 9254 8787 9282 8806
rect 9142 8441 9226 8442
rect 9142 8415 9143 8441
rect 9169 8415 9226 8441
rect 9142 8414 9226 8415
rect 9478 8442 9506 9479
rect 9590 9226 9618 9231
rect 9590 9179 9618 9198
rect 9758 9225 9786 9982
rect 9870 9618 9898 9623
rect 9870 9571 9898 9590
rect 9918 9422 10050 9427
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 9918 9389 10050 9394
rect 9982 9338 10010 9343
rect 9982 9281 10010 9310
rect 9982 9255 9983 9281
rect 10009 9255 10010 9281
rect 9982 9249 10010 9255
rect 9758 9199 9759 9225
rect 9785 9199 9786 9225
rect 9758 9193 9786 9199
rect 9702 9169 9730 9175
rect 9702 9143 9703 9169
rect 9729 9143 9730 9169
rect 9142 8409 9170 8414
rect 9478 8409 9506 8414
rect 9646 8442 9674 8447
rect 9534 8386 9562 8391
rect 9478 8274 9506 8279
rect 9422 7937 9450 7943
rect 9422 7911 9423 7937
rect 9449 7911 9450 7937
rect 9422 7574 9450 7911
rect 9478 7769 9506 8246
rect 9534 8049 9562 8358
rect 9534 8023 9535 8049
rect 9561 8023 9562 8049
rect 9534 8017 9562 8023
rect 9478 7743 9479 7769
rect 9505 7743 9506 7769
rect 9478 7737 9506 7743
rect 9646 7769 9674 8414
rect 9702 8386 9730 9143
rect 10094 9170 10122 11326
rect 10150 11297 10178 11438
rect 10150 11271 10151 11297
rect 10177 11271 10178 11297
rect 10150 11265 10178 11271
rect 10206 10794 10234 11494
rect 10262 10906 10290 11662
rect 10318 11657 10346 11662
rect 11998 11578 12026 11583
rect 11942 11577 12026 11578
rect 11942 11551 11999 11577
rect 12025 11551 12026 11577
rect 11942 11550 12026 11551
rect 11494 11242 11522 11247
rect 10822 11185 10850 11191
rect 10822 11159 10823 11185
rect 10849 11159 10850 11185
rect 10318 11074 10346 11079
rect 10318 11027 10346 11046
rect 10822 10962 10850 11159
rect 10822 10929 10850 10934
rect 11158 11129 11186 11135
rect 11158 11103 11159 11129
rect 11185 11103 11186 11129
rect 10262 10873 10290 10878
rect 11158 10905 11186 11103
rect 11158 10879 11159 10905
rect 11185 10879 11186 10905
rect 11158 10873 11186 10879
rect 11494 11074 11522 11214
rect 11494 10905 11522 11046
rect 11494 10879 11495 10905
rect 11521 10879 11522 10905
rect 11494 10873 11522 10879
rect 11886 10906 11914 10911
rect 11886 10859 11914 10878
rect 10318 10850 10346 10855
rect 10318 10849 10458 10850
rect 10318 10823 10319 10849
rect 10345 10823 10458 10849
rect 10318 10822 10458 10823
rect 10318 10817 10346 10822
rect 10262 10794 10290 10799
rect 10206 10793 10290 10794
rect 10206 10767 10263 10793
rect 10289 10767 10290 10793
rect 10206 10766 10290 10767
rect 10206 10514 10234 10519
rect 10206 10066 10234 10486
rect 10206 9617 10234 10038
rect 10206 9591 10207 9617
rect 10233 9591 10234 9617
rect 10206 9585 10234 9591
rect 10262 9338 10290 10766
rect 10318 10738 10346 10743
rect 10318 10681 10346 10710
rect 10318 10655 10319 10681
rect 10345 10655 10346 10681
rect 10318 10649 10346 10655
rect 10430 10570 10458 10822
rect 10598 10849 10626 10855
rect 10598 10823 10599 10849
rect 10625 10823 10626 10849
rect 10430 10537 10458 10542
rect 10542 10793 10570 10799
rect 10542 10767 10543 10793
rect 10569 10767 10570 10793
rect 10542 10514 10570 10767
rect 10542 10481 10570 10486
rect 10486 10458 10514 10463
rect 10374 10430 10486 10458
rect 10374 10401 10402 10430
rect 10486 10425 10514 10430
rect 10374 10375 10375 10401
rect 10401 10375 10402 10401
rect 10374 10369 10402 10375
rect 10318 10290 10346 10295
rect 10598 10290 10626 10823
rect 11046 10849 11074 10855
rect 11046 10823 11047 10849
rect 11073 10823 11074 10849
rect 10710 10794 10738 10799
rect 10710 10747 10738 10766
rect 10990 10793 11018 10799
rect 10990 10767 10991 10793
rect 11017 10767 11018 10793
rect 10822 10738 10850 10743
rect 10822 10514 10850 10710
rect 10822 10481 10850 10486
rect 10934 10570 10962 10575
rect 10878 10458 10906 10463
rect 10318 10289 10626 10290
rect 10318 10263 10319 10289
rect 10345 10263 10626 10289
rect 10318 10262 10626 10263
rect 10654 10401 10682 10407
rect 10654 10375 10655 10401
rect 10681 10375 10682 10401
rect 10318 9618 10346 10262
rect 10654 10010 10682 10375
rect 10878 10401 10906 10430
rect 10878 10375 10879 10401
rect 10905 10375 10906 10401
rect 10878 10369 10906 10375
rect 10654 9977 10682 9982
rect 10654 9786 10682 9791
rect 10318 9585 10346 9590
rect 10598 9758 10654 9786
rect 10374 9505 10402 9511
rect 10374 9479 10375 9505
rect 10401 9479 10402 9505
rect 10374 9394 10402 9479
rect 10374 9361 10402 9366
rect 10486 9506 10514 9511
rect 10262 9305 10290 9310
rect 10374 9282 10402 9287
rect 10094 9137 10122 9142
rect 10150 9225 10178 9231
rect 10150 9199 10151 9225
rect 10177 9199 10178 9225
rect 9870 8946 9898 8951
rect 9870 8833 9898 8918
rect 9870 8807 9871 8833
rect 9897 8807 9898 8833
rect 9870 8801 9898 8807
rect 9982 8834 10010 8839
rect 9982 8787 10010 8806
rect 9926 8722 9954 8727
rect 9702 8353 9730 8358
rect 9758 8721 9954 8722
rect 9758 8695 9927 8721
rect 9953 8695 9954 8721
rect 9758 8694 9954 8695
rect 9646 7743 9647 7769
rect 9673 7743 9674 7769
rect 9646 7574 9674 7743
rect 9758 7714 9786 8694
rect 9926 8689 9954 8694
rect 9918 8638 10050 8643
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 9918 8605 10050 8610
rect 10150 8498 10178 9199
rect 10374 9225 10402 9254
rect 10486 9281 10514 9478
rect 10486 9255 10487 9281
rect 10513 9255 10514 9281
rect 10486 9249 10514 9255
rect 10374 9199 10375 9225
rect 10401 9199 10402 9225
rect 10374 9193 10402 9199
rect 10206 8834 10234 8839
rect 10598 8834 10626 9758
rect 10654 9753 10682 9758
rect 10822 9618 10850 9623
rect 10822 9571 10850 9590
rect 10654 9561 10682 9567
rect 10654 9535 10655 9561
rect 10681 9535 10682 9561
rect 10654 9170 10682 9535
rect 10934 9225 10962 10542
rect 10990 9954 11018 10767
rect 11046 10794 11074 10823
rect 11774 10850 11802 10855
rect 11774 10803 11802 10822
rect 11046 10761 11074 10766
rect 11270 10793 11298 10799
rect 11270 10767 11271 10793
rect 11297 10767 11298 10793
rect 11270 10682 11298 10767
rect 11382 10793 11410 10799
rect 11382 10767 11383 10793
rect 11409 10767 11410 10793
rect 11270 10649 11298 10654
rect 11326 10737 11354 10743
rect 11326 10711 11327 10737
rect 11353 10711 11354 10737
rect 11326 10626 11354 10711
rect 11382 10738 11410 10767
rect 11382 10705 11410 10710
rect 11438 10794 11466 10799
rect 11326 10593 11354 10598
rect 11158 10402 11186 10407
rect 11158 10065 11186 10374
rect 11158 10039 11159 10065
rect 11185 10039 11186 10065
rect 11158 10033 11186 10039
rect 10990 9921 11018 9926
rect 11326 9842 11354 9847
rect 11046 9617 11074 9623
rect 11046 9591 11047 9617
rect 11073 9591 11074 9617
rect 11046 9394 11074 9591
rect 11046 9361 11074 9366
rect 10934 9199 10935 9225
rect 10961 9199 10962 9225
rect 10934 9193 10962 9199
rect 11102 9337 11130 9343
rect 11102 9311 11103 9337
rect 11129 9311 11130 9337
rect 10682 9142 10738 9170
rect 10654 9137 10682 9142
rect 10206 8833 10626 8834
rect 10206 8807 10207 8833
rect 10233 8807 10626 8833
rect 10206 8806 10626 8807
rect 10206 8801 10234 8806
rect 10598 8553 10626 8806
rect 10598 8527 10599 8553
rect 10625 8527 10626 8553
rect 10598 8521 10626 8527
rect 10654 9002 10682 9007
rect 10654 8833 10682 8974
rect 10654 8807 10655 8833
rect 10681 8807 10682 8833
rect 10150 8465 10178 8470
rect 10038 8441 10066 8447
rect 10038 8415 10039 8441
rect 10065 8415 10066 8441
rect 10038 8386 10066 8415
rect 10206 8442 10234 8447
rect 10206 8395 10234 8414
rect 10654 8441 10682 8807
rect 10710 8777 10738 9142
rect 11102 9058 11130 9311
rect 11326 9337 11354 9814
rect 11438 9729 11466 10766
rect 11942 10682 11970 11550
rect 11998 11545 12026 11550
rect 12110 11578 12138 11583
rect 12110 11531 12138 11550
rect 12278 11577 12306 11583
rect 12278 11551 12279 11577
rect 12305 11551 12306 11577
rect 12054 11521 12082 11527
rect 12054 11495 12055 11521
rect 12081 11495 12082 11521
rect 12054 11186 12082 11495
rect 12054 11153 12082 11158
rect 12222 11241 12250 11247
rect 12222 11215 12223 11241
rect 12249 11215 12250 11241
rect 12166 11130 12194 11135
rect 11998 10906 12026 10911
rect 11998 10859 12026 10878
rect 12166 10905 12194 11102
rect 12166 10879 12167 10905
rect 12193 10879 12194 10905
rect 12166 10873 12194 10879
rect 11942 10649 11970 10654
rect 12110 10793 12138 10799
rect 12110 10767 12111 10793
rect 12137 10767 12138 10793
rect 11438 9703 11439 9729
rect 11465 9703 11466 9729
rect 11438 9697 11466 9703
rect 11886 10458 11914 10463
rect 11606 9617 11634 9623
rect 11606 9591 11607 9617
rect 11633 9591 11634 9617
rect 11326 9311 11327 9337
rect 11353 9311 11354 9337
rect 11326 9305 11354 9311
rect 11438 9394 11466 9399
rect 11438 9337 11466 9366
rect 11438 9311 11439 9337
rect 11465 9311 11466 9337
rect 11438 9305 11466 9311
rect 11550 9338 11578 9343
rect 11550 9291 11578 9310
rect 11606 9226 11634 9591
rect 11830 9617 11858 9623
rect 11830 9591 11831 9617
rect 11857 9591 11858 9617
rect 11718 9562 11746 9567
rect 11830 9562 11858 9591
rect 11718 9561 11858 9562
rect 11718 9535 11719 9561
rect 11745 9535 11858 9561
rect 11718 9534 11858 9535
rect 11718 9338 11746 9534
rect 11774 9338 11802 9343
rect 11718 9310 11774 9338
rect 11774 9291 11802 9310
rect 11606 9193 11634 9198
rect 11886 9225 11914 10430
rect 12110 9730 12138 10767
rect 12222 10458 12250 11215
rect 12222 10425 12250 10430
rect 12278 10066 12306 11551
rect 12558 11185 12586 11998
rect 12670 11746 12698 12391
rect 12726 12418 12754 12423
rect 12782 12418 12810 13118
rect 12838 13113 12866 13118
rect 12950 12866 12978 13175
rect 13006 13202 13034 13207
rect 13118 13202 13146 13426
rect 13510 13426 13538 13431
rect 13510 13425 13818 13426
rect 13510 13399 13511 13425
rect 13537 13399 13818 13425
rect 13510 13398 13818 13399
rect 13510 13393 13538 13398
rect 13006 13201 13146 13202
rect 13006 13175 13007 13201
rect 13033 13175 13146 13201
rect 13006 13174 13146 13175
rect 13006 13169 13034 13174
rect 12950 12833 12978 12838
rect 13174 13145 13202 13151
rect 13174 13119 13175 13145
rect 13201 13119 13202 13145
rect 13174 12642 13202 13119
rect 13566 13090 13594 13095
rect 13566 13089 13650 13090
rect 13566 13063 13567 13089
rect 13593 13063 13650 13089
rect 13566 13062 13650 13063
rect 13566 13057 13594 13062
rect 13510 12866 13538 12871
rect 13510 12809 13538 12838
rect 13510 12783 13511 12809
rect 13537 12783 13538 12809
rect 13510 12777 13538 12783
rect 13622 12753 13650 13062
rect 13622 12727 13623 12753
rect 13649 12727 13650 12753
rect 13622 12721 13650 12727
rect 13790 12753 13818 13398
rect 14630 13202 14658 13454
rect 18830 13258 18858 13511
rect 18830 13225 18858 13230
rect 14798 13202 14826 13207
rect 14630 13201 14826 13202
rect 14630 13175 14799 13201
rect 14825 13175 14826 13201
rect 14630 13174 14826 13175
rect 14630 13089 14658 13174
rect 14630 13063 14631 13089
rect 14657 13063 14658 13089
rect 14630 13057 14658 13063
rect 14798 13090 14826 13174
rect 14966 13202 14994 13207
rect 14966 13155 14994 13174
rect 18830 13146 18858 13151
rect 18830 13099 18858 13118
rect 14798 13057 14826 13062
rect 17598 12950 17730 12955
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17598 12917 17730 12922
rect 18942 12866 18970 13903
rect 19950 13873 19978 13879
rect 19950 13847 19951 13873
rect 19977 13847 19978 13873
rect 19950 13482 19978 13847
rect 19950 13449 19978 13454
rect 20006 13593 20034 13599
rect 20006 13567 20007 13593
rect 20033 13567 20034 13593
rect 20006 13146 20034 13567
rect 20006 13113 20034 13118
rect 18942 12833 18970 12838
rect 20006 13033 20034 13039
rect 20006 13007 20007 13033
rect 20033 13007 20034 13033
rect 20006 12810 20034 13007
rect 20006 12777 20034 12782
rect 13790 12727 13791 12753
rect 13817 12727 13818 12753
rect 13790 12721 13818 12727
rect 13174 12609 13202 12614
rect 13398 12642 13426 12647
rect 12726 12417 12810 12418
rect 12726 12391 12727 12417
rect 12753 12391 12810 12417
rect 12726 12390 12810 12391
rect 12726 12385 12754 12390
rect 13230 11802 13258 11807
rect 12670 11718 12978 11746
rect 12726 11634 12754 11639
rect 12726 11587 12754 11606
rect 12558 11159 12559 11185
rect 12585 11159 12586 11185
rect 12334 10962 12362 10967
rect 12334 10794 12362 10934
rect 12334 10747 12362 10766
rect 12390 10626 12418 10631
rect 12334 10178 12362 10183
rect 12334 10066 12362 10150
rect 12278 10065 12362 10066
rect 12278 10039 12279 10065
rect 12305 10039 12362 10065
rect 12278 10038 12362 10039
rect 12278 10033 12306 10038
rect 12222 10009 12250 10015
rect 12222 9983 12223 10009
rect 12249 9983 12250 10009
rect 12222 9730 12250 9983
rect 12278 9954 12306 9959
rect 12278 9897 12306 9926
rect 12278 9871 12279 9897
rect 12305 9871 12306 9897
rect 12278 9865 12306 9871
rect 12110 9729 12194 9730
rect 12110 9703 12111 9729
rect 12137 9703 12194 9729
rect 12110 9702 12194 9703
rect 12110 9697 12138 9702
rect 12110 9338 12138 9343
rect 12110 9291 12138 9310
rect 11886 9199 11887 9225
rect 11913 9199 11914 9225
rect 11886 9193 11914 9199
rect 11382 9170 11410 9175
rect 11102 9025 11130 9030
rect 11326 9169 11410 9170
rect 11326 9143 11383 9169
rect 11409 9143 11410 9169
rect 11326 9142 11410 9143
rect 10710 8751 10711 8777
rect 10737 8751 10738 8777
rect 10710 8497 10738 8751
rect 10710 8471 10711 8497
rect 10737 8471 10738 8497
rect 10710 8465 10738 8471
rect 10822 8721 10850 8727
rect 10822 8695 10823 8721
rect 10849 8695 10850 8721
rect 10654 8415 10655 8441
rect 10681 8415 10682 8441
rect 10654 8409 10682 8415
rect 10038 8353 10066 8358
rect 10766 8330 10794 8335
rect 10374 7938 10402 7943
rect 9918 7854 10050 7859
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 9918 7821 10050 7826
rect 9758 7681 9786 7686
rect 9814 7770 9842 7775
rect 9814 7574 9842 7742
rect 9254 7546 9282 7551
rect 9030 6847 9031 6873
rect 9057 6847 9058 6873
rect 9030 6841 9058 6847
rect 9198 7265 9226 7271
rect 9198 7239 9199 7265
rect 9225 7239 9226 7265
rect 8974 6785 9002 6790
rect 9198 6594 9226 7239
rect 9254 7265 9282 7518
rect 9254 7239 9255 7265
rect 9281 7239 9282 7265
rect 9254 7233 9282 7239
rect 9366 7546 9450 7574
rect 9534 7546 9674 7574
rect 9758 7546 9842 7574
rect 10374 7657 10402 7910
rect 10374 7631 10375 7657
rect 10401 7631 10402 7657
rect 10038 7546 10066 7551
rect 9366 7434 9394 7546
rect 9534 7513 9562 7518
rect 9758 7434 9786 7546
rect 9366 7406 9786 7434
rect 9366 7265 9394 7406
rect 9646 7322 9674 7327
rect 9366 7239 9367 7265
rect 9393 7239 9394 7265
rect 9366 7233 9394 7239
rect 9422 7266 9450 7271
rect 9422 7219 9450 7238
rect 9646 7265 9674 7294
rect 9646 7239 9647 7265
rect 9673 7239 9674 7265
rect 9646 7233 9674 7239
rect 9758 7265 9786 7406
rect 9758 7239 9759 7265
rect 9785 7239 9786 7265
rect 9758 7233 9786 7239
rect 10038 7265 10066 7518
rect 10038 7239 10039 7265
rect 10065 7239 10066 7265
rect 10038 7233 10066 7239
rect 10374 7266 10402 7631
rect 10486 7770 10514 7775
rect 10766 7770 10794 8302
rect 10486 7769 10794 7770
rect 10486 7743 10487 7769
rect 10513 7743 10794 7769
rect 10486 7742 10794 7743
rect 10486 7322 10514 7742
rect 10766 7713 10794 7742
rect 10766 7687 10767 7713
rect 10793 7687 10794 7713
rect 10766 7681 10794 7687
rect 10822 7714 10850 8695
rect 11326 7994 11354 9142
rect 11382 9137 11410 9142
rect 11606 9114 11634 9119
rect 11270 7938 11298 7943
rect 11270 7891 11298 7910
rect 11326 7826 11354 7966
rect 11550 8498 11578 8503
rect 11438 7938 11466 7943
rect 11438 7891 11466 7910
rect 11270 7798 11354 7826
rect 11382 7882 11410 7887
rect 11270 7769 11298 7798
rect 11270 7743 11271 7769
rect 11297 7743 11298 7769
rect 11270 7737 11298 7743
rect 10878 7714 10906 7719
rect 10822 7713 10906 7714
rect 10822 7687 10879 7713
rect 10905 7687 10906 7713
rect 10822 7686 10906 7687
rect 10878 7658 10906 7686
rect 11382 7713 11410 7854
rect 11382 7687 11383 7713
rect 11409 7687 11410 7713
rect 11382 7681 11410 7687
rect 10878 7625 10906 7630
rect 11102 7657 11130 7663
rect 11102 7631 11103 7657
rect 11129 7631 11130 7657
rect 10486 7289 10514 7294
rect 10710 7602 10738 7607
rect 10374 7219 10402 7238
rect 10710 7266 10738 7574
rect 10990 7601 11018 7607
rect 10990 7575 10991 7601
rect 11017 7575 11018 7601
rect 10990 7322 11018 7575
rect 11102 7574 11130 7631
rect 11326 7657 11354 7663
rect 11326 7631 11327 7657
rect 11353 7631 11354 7657
rect 11102 7546 11242 7574
rect 11326 7546 11354 7631
rect 11214 7518 11354 7546
rect 11438 7658 11466 7663
rect 11046 7322 11074 7327
rect 10990 7321 11074 7322
rect 10990 7295 11047 7321
rect 11073 7295 11074 7321
rect 10990 7294 11074 7295
rect 11046 7289 11074 7294
rect 10710 7219 10738 7238
rect 11214 7266 11242 7271
rect 9926 7210 9954 7215
rect 9926 7163 9954 7182
rect 10262 7209 10290 7215
rect 10262 7183 10263 7209
rect 10289 7183 10290 7209
rect 9310 7153 9338 7159
rect 9310 7127 9311 7153
rect 9337 7127 9338 7153
rect 9254 6873 9282 6879
rect 9254 6847 9255 6873
rect 9281 6847 9282 6873
rect 9254 6818 9282 6847
rect 9310 6874 9338 7127
rect 9702 7153 9730 7159
rect 9702 7127 9703 7153
rect 9729 7127 9730 7153
rect 9702 6986 9730 7127
rect 10150 7154 10178 7159
rect 10150 7107 10178 7126
rect 9918 7070 10050 7075
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 9918 7037 10050 7042
rect 9590 6958 9730 6986
rect 9590 6929 9618 6958
rect 9590 6903 9591 6929
rect 9617 6903 9618 6929
rect 9590 6897 9618 6903
rect 9310 6841 9338 6846
rect 9254 6785 9282 6790
rect 9646 6818 9674 6823
rect 10262 6818 10290 7183
rect 10654 6818 10682 6823
rect 10262 6817 10682 6818
rect 10262 6791 10655 6817
rect 10681 6791 10682 6817
rect 10262 6790 10682 6791
rect 9310 6594 9338 6599
rect 9198 6593 9338 6594
rect 9198 6567 9311 6593
rect 9337 6567 9338 6593
rect 9198 6566 9338 6567
rect 9310 6561 9338 6566
rect 8078 6511 8079 6537
rect 8105 6511 8106 6537
rect 8078 6505 8106 6511
rect 8806 6538 8834 6543
rect 7742 6455 7743 6481
rect 7769 6455 7770 6481
rect 7742 6449 7770 6455
rect 2238 5894 2370 5899
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2238 5861 2370 5866
rect 2238 5110 2370 5115
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2238 5077 2370 5082
rect 2238 4326 2370 4331
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2238 4293 2370 4298
rect 2238 3542 2370 3547
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2238 3509 2370 3514
rect 2238 2758 2370 2763
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2238 2725 2370 2730
rect 2238 1974 2370 1979
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2238 1941 2370 1946
rect 8806 1777 8834 6510
rect 9142 6538 9170 6543
rect 9142 6491 9170 6510
rect 9366 6538 9394 6543
rect 9366 6491 9394 6510
rect 9646 6537 9674 6790
rect 9646 6511 9647 6537
rect 9673 6511 9674 6537
rect 9646 6505 9674 6511
rect 9918 6286 10050 6291
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 9918 6253 10050 6258
rect 9918 5502 10050 5507
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 9918 5469 10050 5474
rect 9918 4718 10050 4723
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 9918 4685 10050 4690
rect 10654 4214 10682 6790
rect 11214 6481 11242 7238
rect 11438 6929 11466 7630
rect 11494 7658 11522 7663
rect 11550 7658 11578 8470
rect 11494 7657 11578 7658
rect 11494 7631 11495 7657
rect 11521 7631 11578 7657
rect 11494 7630 11578 7631
rect 11606 7657 11634 9086
rect 12166 8834 12194 9702
rect 12222 9697 12250 9702
rect 12278 9282 12306 9287
rect 12334 9282 12362 10038
rect 12390 10122 12418 10598
rect 12390 9617 12418 10094
rect 12390 9591 12391 9617
rect 12417 9591 12418 9617
rect 12390 9585 12418 9591
rect 12502 10010 12530 10015
rect 12502 9617 12530 9982
rect 12502 9591 12503 9617
rect 12529 9591 12530 9617
rect 12502 9394 12530 9591
rect 12502 9361 12530 9366
rect 12278 9281 12362 9282
rect 12278 9255 12279 9281
rect 12305 9255 12362 9281
rect 12278 9254 12362 9255
rect 12278 9114 12306 9254
rect 12558 9226 12586 11159
rect 12614 11578 12642 11583
rect 12614 10793 12642 11550
rect 12782 11578 12810 11583
rect 12782 11531 12810 11550
rect 12726 11465 12754 11471
rect 12726 11439 12727 11465
rect 12753 11439 12754 11465
rect 12670 11186 12698 11191
rect 12726 11186 12754 11439
rect 12670 11185 12754 11186
rect 12670 11159 12671 11185
rect 12697 11159 12754 11185
rect 12670 11158 12754 11159
rect 12838 11242 12866 11247
rect 12670 11153 12698 11158
rect 12726 11073 12754 11079
rect 12726 11047 12727 11073
rect 12753 11047 12754 11073
rect 12670 11018 12698 11023
rect 12670 10905 12698 10990
rect 12726 10962 12754 11047
rect 12782 11074 12810 11079
rect 12782 11027 12810 11046
rect 12782 10962 12810 10967
rect 12726 10934 12782 10962
rect 12782 10929 12810 10934
rect 12670 10879 12671 10905
rect 12697 10879 12698 10905
rect 12670 10873 12698 10879
rect 12614 10767 12615 10793
rect 12641 10767 12642 10793
rect 12614 10738 12642 10767
rect 12614 10122 12642 10710
rect 12726 10849 12754 10855
rect 12726 10823 12727 10849
rect 12753 10823 12754 10849
rect 12726 10626 12754 10823
rect 12726 10593 12754 10598
rect 12782 10849 12810 10855
rect 12782 10823 12783 10849
rect 12809 10823 12810 10849
rect 12614 10089 12642 10094
rect 12726 10514 12754 10519
rect 12726 10065 12754 10486
rect 12782 10178 12810 10823
rect 12782 10145 12810 10150
rect 12726 10039 12727 10065
rect 12753 10039 12754 10065
rect 12726 10033 12754 10039
rect 12838 10065 12866 11214
rect 12894 11186 12922 11191
rect 12894 11139 12922 11158
rect 12950 10906 12978 11718
rect 12950 10873 12978 10878
rect 13006 11690 13034 11695
rect 13006 11577 13034 11662
rect 13006 11551 13007 11577
rect 13033 11551 13034 11577
rect 12894 10850 12922 10855
rect 12894 10803 12922 10822
rect 12950 10794 12978 10799
rect 13006 10794 13034 11551
rect 13230 11185 13258 11774
rect 13398 11690 13426 12614
rect 13734 12641 13762 12647
rect 13734 12615 13735 12641
rect 13761 12615 13762 12641
rect 13734 11802 13762 12615
rect 14014 12642 14042 12647
rect 14014 12595 14042 12614
rect 17598 12166 17730 12171
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17598 12133 17730 12138
rect 13734 11769 13762 11774
rect 13398 11657 13426 11662
rect 14630 11690 14658 11695
rect 14630 11643 14658 11662
rect 18830 11578 18858 11583
rect 18830 11531 18858 11550
rect 13342 11522 13370 11527
rect 13230 11159 13231 11185
rect 13257 11159 13258 11185
rect 13062 11074 13090 11079
rect 13062 11027 13090 11046
rect 12978 10766 13034 10794
rect 12950 10761 12978 10766
rect 13230 10514 13258 11159
rect 13286 11521 13370 11522
rect 13286 11495 13343 11521
rect 13369 11495 13370 11521
rect 13286 11494 13370 11495
rect 13286 10962 13314 11494
rect 13342 11489 13370 11494
rect 14406 11522 14434 11527
rect 14406 11475 14434 11494
rect 20006 11466 20034 11471
rect 20006 11419 20034 11438
rect 17598 11382 17730 11387
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17598 11349 17730 11354
rect 13342 11242 13370 11247
rect 13342 11195 13370 11214
rect 20006 11241 20034 11247
rect 20006 11215 20007 11241
rect 20033 11215 20034 11241
rect 13790 11186 13818 11191
rect 13790 11139 13818 11158
rect 18830 11185 18858 11191
rect 18830 11159 18831 11185
rect 18857 11159 18858 11185
rect 13286 10929 13314 10934
rect 13510 11129 13538 11135
rect 13510 11103 13511 11129
rect 13537 11103 13538 11129
rect 13230 10481 13258 10486
rect 13342 10794 13370 10799
rect 13342 10346 13370 10766
rect 13398 10346 13426 10351
rect 13342 10345 13426 10346
rect 13342 10319 13399 10345
rect 13425 10319 13426 10345
rect 13342 10318 13426 10319
rect 13006 10122 13034 10127
rect 13006 10075 13034 10094
rect 13398 10094 13426 10318
rect 13510 10122 13538 11103
rect 13622 11129 13650 11135
rect 13622 11103 13623 11129
rect 13649 11103 13650 11129
rect 13622 11018 13650 11103
rect 13622 10985 13650 10990
rect 13678 11073 13706 11079
rect 13678 11047 13679 11073
rect 13705 11047 13706 11073
rect 13678 10849 13706 11047
rect 13678 10823 13679 10849
rect 13705 10823 13706 10849
rect 13678 10817 13706 10823
rect 14742 10794 14770 10799
rect 14742 10737 14770 10766
rect 18830 10794 18858 11159
rect 20006 11130 20034 11215
rect 20006 11097 20034 11102
rect 18830 10761 18858 10766
rect 14742 10711 14743 10737
rect 14769 10711 14770 10737
rect 14742 10705 14770 10711
rect 17598 10598 17730 10603
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17598 10565 17730 10570
rect 12838 10039 12839 10065
rect 12865 10039 12866 10065
rect 12838 10033 12866 10039
rect 13398 10066 13482 10094
rect 13510 10089 13538 10094
rect 12614 10009 12642 10015
rect 12614 9983 12615 10009
rect 12641 9983 12642 10009
rect 12614 9786 12642 9983
rect 13118 10010 13146 10015
rect 13118 9963 13146 9982
rect 13286 10010 13314 10015
rect 12614 9753 12642 9758
rect 12894 9897 12922 9903
rect 12894 9871 12895 9897
rect 12921 9871 12922 9897
rect 12558 9198 12642 9226
rect 12278 9081 12306 9086
rect 12166 8801 12194 8806
rect 12614 8274 12642 9198
rect 12614 8241 12642 8246
rect 12670 8386 12698 8391
rect 12334 8050 12362 8055
rect 11606 7631 11607 7657
rect 11633 7631 11634 7657
rect 11494 7625 11522 7630
rect 11606 7625 11634 7631
rect 11662 7994 11690 7999
rect 11662 7574 11690 7966
rect 11830 7938 11858 7943
rect 11830 7770 11858 7910
rect 12110 7938 12138 7943
rect 11998 7882 12026 7887
rect 12026 7854 12082 7882
rect 11998 7849 12026 7854
rect 11662 7546 11746 7574
rect 11438 6903 11439 6929
rect 11465 6903 11466 6929
rect 11438 6897 11466 6903
rect 11606 6985 11634 6991
rect 11606 6959 11607 6985
rect 11633 6959 11634 6985
rect 11550 6874 11578 6879
rect 11550 6827 11578 6846
rect 11606 6537 11634 6959
rect 11718 6761 11746 7546
rect 11830 6873 11858 7742
rect 11998 7714 12026 7719
rect 11998 7667 12026 7686
rect 12054 7574 12082 7854
rect 12110 7769 12138 7910
rect 12110 7743 12111 7769
rect 12137 7743 12138 7769
rect 12110 7737 12138 7743
rect 12222 7826 12250 7831
rect 12222 7769 12250 7798
rect 12222 7743 12223 7769
rect 12249 7743 12250 7769
rect 12222 7737 12250 7743
rect 12334 7770 12362 8022
rect 12334 7657 12362 7742
rect 12334 7631 12335 7657
rect 12361 7631 12362 7657
rect 12334 7625 12362 7631
rect 12166 7601 12194 7607
rect 12166 7575 12167 7601
rect 12193 7575 12194 7601
rect 12054 7546 12138 7574
rect 11830 6847 11831 6873
rect 11857 6847 11858 6873
rect 11830 6841 11858 6847
rect 12110 7321 12138 7546
rect 12110 7295 12111 7321
rect 12137 7295 12138 7321
rect 11718 6735 11719 6761
rect 11745 6735 11746 6761
rect 11718 6729 11746 6735
rect 11606 6511 11607 6537
rect 11633 6511 11634 6537
rect 11606 6505 11634 6511
rect 11214 6455 11215 6481
rect 11241 6455 11242 6481
rect 11214 6449 11242 6455
rect 10542 4186 10682 4214
rect 12110 4214 12138 7295
rect 12166 7322 12194 7575
rect 12670 7602 12698 8358
rect 12726 8050 12754 8055
rect 12726 8003 12754 8022
rect 12894 8049 12922 9871
rect 13062 9898 13090 9903
rect 13062 9505 13090 9870
rect 13286 9562 13314 9982
rect 13342 9954 13370 9959
rect 13342 9673 13370 9926
rect 13398 9953 13426 10066
rect 13454 10010 13482 10066
rect 13566 10010 13594 10015
rect 13454 10009 13594 10010
rect 13454 9983 13567 10009
rect 13593 9983 13594 10009
rect 13454 9982 13594 9983
rect 13566 9977 13594 9982
rect 13398 9927 13399 9953
rect 13425 9927 13426 9953
rect 13398 9898 13426 9927
rect 13958 9954 13986 9959
rect 13958 9907 13986 9926
rect 14686 9954 14714 9959
rect 13398 9865 13426 9870
rect 13342 9647 13343 9673
rect 13369 9647 13370 9673
rect 13342 9641 13370 9647
rect 13398 9674 13426 9679
rect 13566 9674 13594 9679
rect 13398 9673 13594 9674
rect 13398 9647 13399 9673
rect 13425 9647 13567 9673
rect 13593 9647 13594 9673
rect 13398 9646 13594 9647
rect 13398 9641 13426 9646
rect 13566 9641 13594 9646
rect 13734 9674 13762 9679
rect 13958 9674 13986 9679
rect 13734 9673 13986 9674
rect 13734 9647 13735 9673
rect 13761 9647 13959 9673
rect 13985 9647 13986 9673
rect 13734 9646 13986 9647
rect 13734 9641 13762 9646
rect 13958 9641 13986 9646
rect 14686 9673 14714 9926
rect 15022 9954 15050 9959
rect 15022 9907 15050 9926
rect 18830 9954 18858 9959
rect 17598 9814 17730 9819
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17598 9781 17730 9786
rect 14686 9647 14687 9673
rect 14713 9647 14714 9673
rect 14686 9641 14714 9647
rect 14070 9618 14098 9623
rect 14070 9571 14098 9590
rect 14630 9618 14658 9623
rect 14630 9571 14658 9590
rect 18830 9617 18858 9926
rect 18830 9591 18831 9617
rect 18857 9591 18858 9617
rect 18830 9585 18858 9591
rect 20006 9673 20034 9679
rect 20006 9647 20007 9673
rect 20033 9647 20034 9673
rect 13062 9479 13063 9505
rect 13089 9479 13090 9505
rect 12950 9170 12978 9175
rect 13062 9170 13090 9479
rect 13230 9561 13314 9562
rect 13230 9535 13287 9561
rect 13313 9535 13314 9561
rect 13230 9534 13314 9535
rect 13118 9225 13146 9231
rect 13118 9199 13119 9225
rect 13145 9199 13146 9225
rect 13118 9170 13146 9199
rect 12950 9169 13146 9170
rect 12950 9143 12951 9169
rect 12977 9143 13146 9169
rect 12950 9142 13146 9143
rect 13174 9170 13202 9175
rect 12950 8386 12978 9142
rect 13062 9058 13090 9063
rect 13062 8833 13090 9030
rect 13062 8807 13063 8833
rect 13089 8807 13090 8833
rect 13062 8801 13090 8807
rect 13174 8834 13202 9142
rect 13174 8787 13202 8806
rect 12950 8353 12978 8358
rect 13006 8385 13034 8391
rect 13006 8359 13007 8385
rect 13033 8359 13034 8385
rect 13006 8274 13034 8359
rect 13230 8330 13258 9534
rect 13286 9529 13314 9534
rect 13902 9561 13930 9567
rect 13902 9535 13903 9561
rect 13929 9535 13930 9561
rect 13622 9506 13650 9511
rect 13622 9459 13650 9478
rect 13510 9170 13538 9175
rect 13454 9169 13538 9170
rect 13454 9143 13511 9169
rect 13537 9143 13538 9169
rect 13454 9142 13538 9143
rect 13286 8834 13314 8839
rect 13286 8787 13314 8806
rect 13342 8833 13370 8839
rect 13342 8807 13343 8833
rect 13369 8807 13370 8833
rect 13230 8297 13258 8302
rect 13006 8241 13034 8246
rect 13286 8274 13314 8279
rect 12894 8023 12895 8049
rect 12921 8023 12922 8049
rect 12894 8017 12922 8023
rect 13286 8049 13314 8246
rect 13286 8023 13287 8049
rect 13313 8023 13314 8049
rect 13006 7994 13034 7999
rect 13118 7994 13146 7999
rect 13006 7993 13146 7994
rect 13006 7967 13007 7993
rect 13033 7967 13119 7993
rect 13145 7967 13146 7993
rect 13006 7966 13146 7967
rect 13006 7961 13034 7966
rect 13118 7961 13146 7966
rect 13286 7994 13314 8023
rect 13342 8050 13370 8807
rect 13454 8721 13482 9142
rect 13510 9137 13538 9142
rect 13790 9170 13818 9175
rect 13902 9170 13930 9535
rect 20006 9450 20034 9647
rect 20006 9417 20034 9422
rect 18830 9226 18858 9231
rect 18830 9179 18858 9198
rect 13818 9142 13930 9170
rect 13958 9170 13986 9175
rect 13790 8945 13818 9142
rect 13790 8919 13791 8945
rect 13817 8919 13818 8945
rect 13790 8913 13818 8919
rect 13846 8834 13874 8839
rect 13846 8787 13874 8806
rect 13958 8833 13986 9142
rect 14574 9170 14602 9175
rect 14574 9123 14602 9142
rect 20006 9114 20034 9119
rect 20006 9067 20034 9086
rect 17598 9030 17730 9035
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17598 8997 17730 9002
rect 13958 8807 13959 8833
rect 13985 8807 13986 8833
rect 13958 8801 13986 8807
rect 13454 8695 13455 8721
rect 13481 8695 13482 8721
rect 13454 8689 13482 8695
rect 13342 8017 13370 8022
rect 14462 8386 14490 8391
rect 13286 7961 13314 7966
rect 13566 7994 13594 7999
rect 13566 7947 13594 7966
rect 13790 7994 13818 7999
rect 13790 7947 13818 7966
rect 12782 7937 12810 7943
rect 12782 7911 12783 7937
rect 12809 7911 12810 7937
rect 12782 7826 12810 7911
rect 12782 7793 12810 7798
rect 12838 7937 12866 7943
rect 12838 7911 12839 7937
rect 12865 7911 12866 7937
rect 12838 7770 12866 7911
rect 13230 7937 13258 7943
rect 13230 7911 13231 7937
rect 13257 7911 13258 7937
rect 12838 7742 13202 7770
rect 13174 7713 13202 7742
rect 13174 7687 13175 7713
rect 13201 7687 13202 7713
rect 13174 7681 13202 7687
rect 12670 7569 12698 7574
rect 12782 7657 12810 7663
rect 12782 7631 12783 7657
rect 12809 7631 12810 7657
rect 12166 7289 12194 7294
rect 12334 7266 12362 7271
rect 12334 7219 12362 7238
rect 12614 7266 12642 7271
rect 12782 7266 12810 7631
rect 13230 7602 13258 7911
rect 13398 7938 13426 7943
rect 13398 7891 13426 7910
rect 13510 7937 13538 7943
rect 13510 7911 13511 7937
rect 13537 7911 13538 7937
rect 13510 7882 13538 7911
rect 13510 7849 13538 7854
rect 14070 7882 14098 7887
rect 13230 7569 13258 7574
rect 13006 7322 13034 7327
rect 13006 7275 13034 7294
rect 14070 7321 14098 7854
rect 14238 7602 14266 7607
rect 14238 7555 14266 7574
rect 14462 7601 14490 8358
rect 17598 8246 17730 8251
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17598 8213 17730 8218
rect 20006 8105 20034 8111
rect 20006 8079 20007 8105
rect 20033 8079 20034 8105
rect 18942 8049 18970 8055
rect 18942 8023 18943 8049
rect 18969 8023 18970 8049
rect 18830 7882 18858 7887
rect 18830 7657 18858 7854
rect 18830 7631 18831 7657
rect 18857 7631 18858 7657
rect 18830 7625 18858 7631
rect 14462 7575 14463 7601
rect 14489 7575 14490 7601
rect 14070 7295 14071 7321
rect 14097 7295 14098 7321
rect 14070 7289 14098 7295
rect 14294 7322 14322 7327
rect 14462 7322 14490 7575
rect 18942 7602 18970 8023
rect 20006 7770 20034 8079
rect 20006 7737 20034 7742
rect 18942 7569 18970 7574
rect 20006 7601 20034 7607
rect 20006 7575 20007 7601
rect 20033 7575 20034 7601
rect 17598 7462 17730 7467
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17598 7429 17730 7434
rect 20006 7434 20034 7575
rect 20006 7401 20034 7406
rect 14294 7321 14490 7322
rect 14294 7295 14295 7321
rect 14321 7295 14490 7321
rect 14294 7294 14490 7295
rect 14294 7289 14322 7294
rect 12642 7238 12978 7266
rect 12614 7219 12642 7238
rect 12166 6874 12194 6879
rect 12166 6827 12194 6846
rect 12222 6817 12250 6823
rect 12222 6791 12223 6817
rect 12249 6791 12250 6817
rect 12222 6538 12250 6791
rect 12222 6505 12250 6510
rect 12614 6538 12642 6543
rect 12670 6538 12698 6543
rect 12642 6537 12698 6538
rect 12642 6511 12671 6537
rect 12697 6511 12698 6537
rect 12642 6510 12698 6511
rect 12110 4186 12306 4214
rect 9918 3934 10050 3939
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 9918 3901 10050 3906
rect 9918 3150 10050 3155
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 9918 3117 10050 3122
rect 9918 2366 10050 2371
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 9918 2333 10050 2338
rect 9310 1834 9338 1839
rect 8806 1751 8807 1777
rect 8833 1751 8834 1777
rect 8806 1745 8834 1751
rect 9086 1833 9338 1834
rect 9086 1807 9311 1833
rect 9337 1807 9338 1833
rect 9086 1806 9338 1807
rect 9086 400 9114 1806
rect 9310 1801 9338 1806
rect 10430 1834 10458 1839
rect 9918 1582 10050 1587
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 9918 1549 10050 1554
rect 10430 400 10458 1806
rect 10542 1777 10570 4186
rect 11046 1834 11074 1839
rect 11046 1787 11074 1806
rect 11438 1834 11466 1839
rect 10542 1751 10543 1777
rect 10569 1751 10570 1777
rect 10542 1745 10570 1751
rect 11438 400 11466 1806
rect 12278 1777 12306 4186
rect 12614 2169 12642 6510
rect 12670 6505 12698 6510
rect 12950 6537 12978 7238
rect 17598 6678 17730 6683
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17598 6645 17730 6650
rect 12950 6511 12951 6537
rect 12977 6511 12978 6537
rect 12950 6505 12978 6511
rect 17598 5894 17730 5899
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17598 5861 17730 5866
rect 17598 5110 17730 5115
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17598 5077 17730 5082
rect 17598 4326 17730 4331
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17598 4293 17730 4298
rect 17598 3542 17730 3547
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17598 3509 17730 3514
rect 17598 2758 17730 2763
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17598 2725 17730 2730
rect 12614 2143 12615 2169
rect 12641 2143 12642 2169
rect 12614 2137 12642 2143
rect 12278 1751 12279 1777
rect 12305 1751 12306 1777
rect 12278 1745 12306 1751
rect 12446 2058 12474 2063
rect 12446 400 12474 2030
rect 13118 2058 13146 2063
rect 13118 2011 13146 2030
rect 17598 1974 17730 1979
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17598 1941 17730 1946
rect 12782 1834 12810 1839
rect 12782 1787 12810 1806
rect 17598 1666 17626 1671
rect 17486 1665 17626 1666
rect 17486 1639 17599 1665
rect 17625 1639 17626 1665
rect 17486 1638 17626 1639
rect 17486 400 17514 1638
rect 17598 1633 17626 1638
rect 9072 0 9128 400
rect 10416 0 10472 400
rect 11424 0 11480 400
rect 12432 0 12488 400
rect 17472 0 17528 400
<< via2 >>
rect 2238 19221 2266 19222
rect 2238 19195 2239 19221
rect 2239 19195 2265 19221
rect 2265 19195 2266 19221
rect 2238 19194 2266 19195
rect 2290 19221 2318 19222
rect 2290 19195 2291 19221
rect 2291 19195 2317 19221
rect 2317 19195 2318 19221
rect 2290 19194 2318 19195
rect 2342 19221 2370 19222
rect 2342 19195 2343 19221
rect 2343 19195 2369 19221
rect 2369 19195 2370 19221
rect 2342 19194 2370 19195
rect 2238 18437 2266 18438
rect 2238 18411 2239 18437
rect 2239 18411 2265 18437
rect 2265 18411 2266 18437
rect 2238 18410 2266 18411
rect 2290 18437 2318 18438
rect 2290 18411 2291 18437
rect 2291 18411 2317 18437
rect 2317 18411 2318 18437
rect 2290 18410 2318 18411
rect 2342 18437 2370 18438
rect 2342 18411 2343 18437
rect 2343 18411 2369 18437
rect 2369 18411 2370 18437
rect 2342 18410 2370 18411
rect 2238 17653 2266 17654
rect 2238 17627 2239 17653
rect 2239 17627 2265 17653
rect 2265 17627 2266 17653
rect 2238 17626 2266 17627
rect 2290 17653 2318 17654
rect 2290 17627 2291 17653
rect 2291 17627 2317 17653
rect 2317 17627 2318 17653
rect 2290 17626 2318 17627
rect 2342 17653 2370 17654
rect 2342 17627 2343 17653
rect 2343 17627 2369 17653
rect 2369 17627 2370 17653
rect 2342 17626 2370 17627
rect 2238 16869 2266 16870
rect 2238 16843 2239 16869
rect 2239 16843 2265 16869
rect 2265 16843 2266 16869
rect 2238 16842 2266 16843
rect 2290 16869 2318 16870
rect 2290 16843 2291 16869
rect 2291 16843 2317 16869
rect 2317 16843 2318 16869
rect 2290 16842 2318 16843
rect 2342 16869 2370 16870
rect 2342 16843 2343 16869
rect 2343 16843 2369 16869
rect 2369 16843 2370 16869
rect 2342 16842 2370 16843
rect 2238 16085 2266 16086
rect 2238 16059 2239 16085
rect 2239 16059 2265 16085
rect 2265 16059 2266 16085
rect 2238 16058 2266 16059
rect 2290 16085 2318 16086
rect 2290 16059 2291 16085
rect 2291 16059 2317 16085
rect 2317 16059 2318 16085
rect 2290 16058 2318 16059
rect 2342 16085 2370 16086
rect 2342 16059 2343 16085
rect 2343 16059 2369 16085
rect 2369 16059 2370 16085
rect 2342 16058 2370 16059
rect 9918 18829 9946 18830
rect 9918 18803 9919 18829
rect 9919 18803 9945 18829
rect 9945 18803 9946 18829
rect 9918 18802 9946 18803
rect 9970 18829 9998 18830
rect 9970 18803 9971 18829
rect 9971 18803 9997 18829
rect 9997 18803 9998 18829
rect 9970 18802 9998 18803
rect 10022 18829 10050 18830
rect 10022 18803 10023 18829
rect 10023 18803 10049 18829
rect 10049 18803 10050 18829
rect 10022 18802 10050 18803
rect 10430 19110 10458 19138
rect 11046 19137 11074 19138
rect 11046 19111 11047 19137
rect 11047 19111 11073 19137
rect 11073 19111 11074 19137
rect 11046 19110 11074 19111
rect 12782 19278 12810 19306
rect 13398 19278 13426 19306
rect 11438 19110 11466 19138
rect 12782 19137 12810 19138
rect 12782 19111 12783 19137
rect 12783 19111 12809 19137
rect 12809 19111 12810 19137
rect 12782 19110 12810 19111
rect 10094 18718 10122 18746
rect 9918 18045 9946 18046
rect 9918 18019 9919 18045
rect 9919 18019 9945 18045
rect 9945 18019 9946 18045
rect 9918 18018 9946 18019
rect 9970 18045 9998 18046
rect 9970 18019 9971 18045
rect 9971 18019 9997 18045
rect 9997 18019 9998 18045
rect 9970 18018 9998 18019
rect 10022 18045 10050 18046
rect 10022 18019 10023 18045
rect 10023 18019 10049 18045
rect 10049 18019 10050 18045
rect 10022 18018 10050 18019
rect 9918 17261 9946 17262
rect 9918 17235 9919 17261
rect 9919 17235 9945 17261
rect 9945 17235 9946 17261
rect 9918 17234 9946 17235
rect 9970 17261 9998 17262
rect 9970 17235 9971 17261
rect 9971 17235 9997 17261
rect 9997 17235 9998 17261
rect 9970 17234 9998 17235
rect 10022 17261 10050 17262
rect 10022 17235 10023 17261
rect 10023 17235 10049 17261
rect 10049 17235 10050 17261
rect 10022 17234 10050 17235
rect 9918 16477 9946 16478
rect 9918 16451 9919 16477
rect 9919 16451 9945 16477
rect 9945 16451 9946 16477
rect 9918 16450 9946 16451
rect 9970 16477 9998 16478
rect 9970 16451 9971 16477
rect 9971 16451 9997 16477
rect 9997 16451 9998 16477
rect 9970 16450 9998 16451
rect 10022 16477 10050 16478
rect 10022 16451 10023 16477
rect 10023 16451 10049 16477
rect 10049 16451 10050 16477
rect 10022 16450 10050 16451
rect 2238 15301 2266 15302
rect 2238 15275 2239 15301
rect 2239 15275 2265 15301
rect 2265 15275 2266 15301
rect 2238 15274 2266 15275
rect 2290 15301 2318 15302
rect 2290 15275 2291 15301
rect 2291 15275 2317 15301
rect 2317 15275 2318 15301
rect 2290 15274 2318 15275
rect 2342 15301 2370 15302
rect 2342 15275 2343 15301
rect 2343 15275 2369 15301
rect 2369 15275 2370 15301
rect 2342 15274 2370 15275
rect 2238 14517 2266 14518
rect 2238 14491 2239 14517
rect 2239 14491 2265 14517
rect 2265 14491 2266 14517
rect 2238 14490 2266 14491
rect 2290 14517 2318 14518
rect 2290 14491 2291 14517
rect 2291 14491 2317 14517
rect 2317 14491 2318 14517
rect 2290 14490 2318 14491
rect 2342 14517 2370 14518
rect 2342 14491 2343 14517
rect 2343 14491 2369 14517
rect 2369 14491 2370 14517
rect 2342 14490 2370 14491
rect 2238 13733 2266 13734
rect 2238 13707 2239 13733
rect 2239 13707 2265 13733
rect 2265 13707 2266 13733
rect 2238 13706 2266 13707
rect 2290 13733 2318 13734
rect 2290 13707 2291 13733
rect 2291 13707 2317 13733
rect 2317 13707 2318 13733
rect 2290 13706 2318 13707
rect 2342 13733 2370 13734
rect 2342 13707 2343 13733
rect 2343 13707 2369 13733
rect 2369 13707 2370 13733
rect 2342 13706 2370 13707
rect 2142 13537 2170 13538
rect 2142 13511 2143 13537
rect 2143 13511 2169 13537
rect 2169 13511 2170 13537
rect 2142 13510 2170 13511
rect 6622 13510 6650 13538
rect 966 13118 994 13146
rect 2086 13454 2114 13482
rect 966 12782 994 12810
rect 966 11774 994 11802
rect 966 11241 994 11242
rect 966 11215 967 11241
rect 967 11215 993 11241
rect 993 11215 994 11241
rect 966 11214 994 11215
rect 2142 13145 2170 13146
rect 2142 13119 2143 13145
rect 2143 13119 2169 13145
rect 2169 13119 2170 13145
rect 2142 13118 2170 13119
rect 5950 13118 5978 13146
rect 2238 12949 2266 12950
rect 2238 12923 2239 12949
rect 2239 12923 2265 12949
rect 2265 12923 2266 12949
rect 2238 12922 2266 12923
rect 2290 12949 2318 12950
rect 2290 12923 2291 12949
rect 2291 12923 2317 12949
rect 2317 12923 2318 12949
rect 2290 12922 2318 12923
rect 2342 12949 2370 12950
rect 2342 12923 2343 12949
rect 2343 12923 2369 12949
rect 2369 12923 2370 12949
rect 2342 12922 2370 12923
rect 6622 13089 6650 13090
rect 6622 13063 6623 13089
rect 6623 13063 6649 13089
rect 6649 13063 6650 13089
rect 6622 13062 6650 13063
rect 7630 13062 7658 13090
rect 7686 12726 7714 12754
rect 8022 13062 8050 13090
rect 8302 13089 8330 13090
rect 8302 13063 8303 13089
rect 8303 13063 8329 13089
rect 8329 13063 8330 13089
rect 8302 13062 8330 13063
rect 9918 15693 9946 15694
rect 9918 15667 9919 15693
rect 9919 15667 9945 15693
rect 9945 15667 9946 15693
rect 9918 15666 9946 15667
rect 9970 15693 9998 15694
rect 9970 15667 9971 15693
rect 9971 15667 9997 15693
rect 9997 15667 9998 15693
rect 9970 15666 9998 15667
rect 10022 15693 10050 15694
rect 10022 15667 10023 15693
rect 10023 15667 10049 15693
rect 10049 15667 10050 15693
rect 10022 15666 10050 15667
rect 9918 14909 9946 14910
rect 9918 14883 9919 14909
rect 9919 14883 9945 14909
rect 9945 14883 9946 14909
rect 9918 14882 9946 14883
rect 9970 14909 9998 14910
rect 9970 14883 9971 14909
rect 9971 14883 9997 14909
rect 9997 14883 9998 14909
rect 9970 14882 9998 14883
rect 10022 14909 10050 14910
rect 10022 14883 10023 14909
rect 10023 14883 10049 14909
rect 10049 14883 10050 14909
rect 10022 14882 10050 14883
rect 9918 14125 9946 14126
rect 9918 14099 9919 14125
rect 9919 14099 9945 14125
rect 9945 14099 9946 14125
rect 9918 14098 9946 14099
rect 9970 14125 9998 14126
rect 9970 14099 9971 14125
rect 9971 14099 9997 14125
rect 9997 14099 9998 14125
rect 9970 14098 9998 14099
rect 10022 14125 10050 14126
rect 10022 14099 10023 14125
rect 10023 14099 10049 14125
rect 10049 14099 10050 14125
rect 10022 14098 10050 14099
rect 9310 13398 9338 13426
rect 10094 13454 10122 13482
rect 9918 13341 9946 13342
rect 9918 13315 9919 13341
rect 9919 13315 9945 13341
rect 9945 13315 9946 13341
rect 9918 13314 9946 13315
rect 9970 13341 9998 13342
rect 9970 13315 9971 13341
rect 9971 13315 9997 13341
rect 9997 13315 9998 13341
rect 9970 13314 9998 13315
rect 10022 13341 10050 13342
rect 10022 13315 10023 13341
rect 10023 13315 10049 13341
rect 10049 13315 10050 13341
rect 10022 13314 10050 13315
rect 9702 13257 9730 13258
rect 9702 13231 9703 13257
rect 9703 13231 9729 13257
rect 9729 13231 9730 13257
rect 9702 13230 9730 13231
rect 9198 13201 9226 13202
rect 9198 13175 9199 13201
rect 9199 13175 9225 13201
rect 9225 13175 9226 13201
rect 9198 13174 9226 13175
rect 9478 13174 9506 13202
rect 8974 13062 9002 13090
rect 8974 12782 9002 12810
rect 7350 12697 7378 12698
rect 7350 12671 7351 12697
rect 7351 12671 7377 12697
rect 7377 12671 7378 12697
rect 7350 12670 7378 12671
rect 6846 12502 6874 12530
rect 7406 12390 7434 12418
rect 5950 12334 5978 12362
rect 2238 12165 2266 12166
rect 2238 12139 2239 12165
rect 2239 12139 2265 12165
rect 2265 12139 2266 12165
rect 2238 12138 2266 12139
rect 2290 12165 2318 12166
rect 2290 12139 2291 12165
rect 2291 12139 2317 12165
rect 2317 12139 2318 12165
rect 2290 12138 2318 12139
rect 2342 12165 2370 12166
rect 2342 12139 2343 12165
rect 2343 12139 2369 12165
rect 2369 12139 2370 12165
rect 2342 12138 2370 12139
rect 2142 11969 2170 11970
rect 2142 11943 2143 11969
rect 2143 11943 2169 11969
rect 2169 11943 2170 11969
rect 2142 11942 2170 11943
rect 5670 11942 5698 11970
rect 2238 11381 2266 11382
rect 2238 11355 2239 11381
rect 2239 11355 2265 11381
rect 2265 11355 2266 11381
rect 2238 11354 2266 11355
rect 2290 11381 2318 11382
rect 2290 11355 2291 11381
rect 2291 11355 2317 11381
rect 2317 11355 2318 11381
rect 2290 11354 2318 11355
rect 2342 11381 2370 11382
rect 2342 11355 2343 11381
rect 2343 11355 2369 11381
rect 2369 11355 2370 11381
rect 2342 11354 2370 11355
rect 6734 11046 6762 11074
rect 6790 11494 6818 11522
rect 2142 10822 2170 10850
rect 5726 10822 5754 10850
rect 2086 10710 2114 10738
rect 7406 11942 7434 11970
rect 7630 12473 7658 12474
rect 7630 12447 7631 12473
rect 7631 12447 7657 12473
rect 7657 12447 7658 12473
rect 7630 12446 7658 12447
rect 7742 12502 7770 12530
rect 7574 12390 7602 12418
rect 7686 12361 7714 12362
rect 7686 12335 7687 12361
rect 7687 12335 7713 12361
rect 7713 12335 7714 12361
rect 7686 12334 7714 12335
rect 7294 11185 7322 11186
rect 7294 11159 7295 11185
rect 7295 11159 7321 11185
rect 7321 11159 7322 11185
rect 7294 11158 7322 11159
rect 7350 11073 7378 11074
rect 7350 11047 7351 11073
rect 7351 11047 7377 11073
rect 7377 11047 7378 11073
rect 7350 11046 7378 11047
rect 2238 10597 2266 10598
rect 2238 10571 2239 10597
rect 2239 10571 2265 10597
rect 2265 10571 2266 10597
rect 2238 10570 2266 10571
rect 2290 10597 2318 10598
rect 2290 10571 2291 10597
rect 2291 10571 2317 10597
rect 2317 10571 2318 10597
rect 2290 10570 2318 10571
rect 2342 10597 2370 10598
rect 2342 10571 2343 10597
rect 2343 10571 2369 10597
rect 2369 10571 2370 10597
rect 2342 10570 2370 10571
rect 6566 10430 6594 10458
rect 4998 9982 5026 10010
rect 2238 9813 2266 9814
rect 2238 9787 2239 9813
rect 2239 9787 2265 9813
rect 2265 9787 2266 9813
rect 2238 9786 2266 9787
rect 2290 9813 2318 9814
rect 2290 9787 2291 9813
rect 2291 9787 2317 9813
rect 2317 9787 2318 9813
rect 2290 9786 2318 9787
rect 2342 9813 2370 9814
rect 2342 9787 2343 9813
rect 2343 9787 2369 9813
rect 2369 9787 2370 9813
rect 2342 9786 2370 9787
rect 4998 9673 5026 9674
rect 4998 9647 4999 9673
rect 4999 9647 5025 9673
rect 5025 9647 5026 9673
rect 4998 9646 5026 9647
rect 7462 10849 7490 10850
rect 7462 10823 7463 10849
rect 7463 10823 7489 10849
rect 7489 10823 7490 10849
rect 7462 10822 7490 10823
rect 7574 11521 7602 11522
rect 7574 11495 7575 11521
rect 7575 11495 7601 11521
rect 7601 11495 7602 11521
rect 7574 11494 7602 11495
rect 7406 10654 7434 10682
rect 7294 10457 7322 10458
rect 7294 10431 7295 10457
rect 7295 10431 7321 10457
rect 7321 10431 7322 10457
rect 7294 10430 7322 10431
rect 7910 11662 7938 11690
rect 9142 12446 9170 12474
rect 8022 12390 8050 12418
rect 9086 12361 9114 12362
rect 9086 12335 9087 12361
rect 9087 12335 9113 12361
rect 9113 12335 9114 12361
rect 9086 12334 9114 12335
rect 10150 13398 10178 13426
rect 9366 12614 9394 12642
rect 7966 11606 7994 11634
rect 8862 11633 8890 11634
rect 8862 11607 8863 11633
rect 8863 11607 8889 11633
rect 8889 11607 8890 11633
rect 8862 11606 8890 11607
rect 8694 11550 8722 11578
rect 7798 11129 7826 11130
rect 7798 11103 7799 11129
rect 7799 11103 7825 11129
rect 7825 11103 7826 11129
rect 7798 11102 7826 11103
rect 7742 11073 7770 11074
rect 7742 11047 7743 11073
rect 7743 11047 7769 11073
rect 7769 11047 7770 11073
rect 7742 11046 7770 11047
rect 7966 11046 7994 11074
rect 8638 11102 8666 11130
rect 9030 11577 9058 11578
rect 9030 11551 9031 11577
rect 9031 11551 9057 11577
rect 9057 11551 9058 11577
rect 9030 11550 9058 11551
rect 8862 11185 8890 11186
rect 8862 11159 8863 11185
rect 8863 11159 8889 11185
rect 8889 11159 8890 11185
rect 8862 11158 8890 11159
rect 8302 10878 8330 10906
rect 7742 10793 7770 10794
rect 7742 10767 7743 10793
rect 7743 10767 7769 10793
rect 7769 10767 7770 10793
rect 7742 10766 7770 10767
rect 7742 10654 7770 10682
rect 7686 10598 7714 10626
rect 7854 10542 7882 10570
rect 7630 10457 7658 10458
rect 7630 10431 7631 10457
rect 7631 10431 7657 10457
rect 7657 10431 7658 10457
rect 7630 10430 7658 10431
rect 7574 10094 7602 10122
rect 7070 10065 7098 10066
rect 7070 10039 7071 10065
rect 7071 10039 7097 10065
rect 7097 10039 7098 10065
rect 7070 10038 7098 10039
rect 2142 9617 2170 9618
rect 2142 9591 2143 9617
rect 2143 9591 2169 9617
rect 2169 9591 2170 9617
rect 2142 9590 2170 9591
rect 6062 9478 6090 9506
rect 966 9422 994 9450
rect 5054 9225 5082 9226
rect 5054 9199 5055 9225
rect 5055 9199 5081 9225
rect 5081 9199 5082 9225
rect 5054 9198 5082 9199
rect 6958 9617 6986 9618
rect 6958 9591 6959 9617
rect 6959 9591 6985 9617
rect 6985 9591 6986 9617
rect 6958 9590 6986 9591
rect 7406 10065 7434 10066
rect 7406 10039 7407 10065
rect 7407 10039 7433 10065
rect 7433 10039 7434 10065
rect 7406 10038 7434 10039
rect 7238 10009 7266 10010
rect 7238 9983 7239 10009
rect 7239 9983 7265 10009
rect 7265 9983 7266 10009
rect 7238 9982 7266 9983
rect 7294 9758 7322 9786
rect 6902 9505 6930 9506
rect 6902 9479 6903 9505
rect 6903 9479 6929 9505
rect 6929 9479 6930 9505
rect 6902 9478 6930 9479
rect 7742 10065 7770 10066
rect 7742 10039 7743 10065
rect 7743 10039 7769 10065
rect 7769 10039 7770 10065
rect 7742 10038 7770 10039
rect 7742 9897 7770 9898
rect 7742 9871 7743 9897
rect 7743 9871 7769 9897
rect 7769 9871 7770 9897
rect 7742 9870 7770 9871
rect 7574 9702 7602 9730
rect 7742 9646 7770 9674
rect 7686 9590 7714 9618
rect 7630 9561 7658 9562
rect 7630 9535 7631 9561
rect 7631 9535 7657 9561
rect 7657 9535 7658 9561
rect 7630 9534 7658 9535
rect 7630 9366 7658 9394
rect 6398 9198 6426 9226
rect 5390 9169 5418 9170
rect 5390 9143 5391 9169
rect 5391 9143 5417 9169
rect 5417 9143 5418 9169
rect 5390 9142 5418 9143
rect 2238 9029 2266 9030
rect 2238 9003 2239 9029
rect 2239 9003 2265 9029
rect 2265 9003 2266 9029
rect 2238 9002 2266 9003
rect 2290 9029 2318 9030
rect 2290 9003 2291 9029
rect 2291 9003 2317 9029
rect 2317 9003 2318 9029
rect 2290 9002 2318 9003
rect 2342 9029 2370 9030
rect 2342 9003 2343 9029
rect 2343 9003 2369 9029
rect 2369 9003 2370 9029
rect 2342 9002 2370 9003
rect 7630 9254 7658 9282
rect 7126 9086 7154 9114
rect 7462 8918 7490 8946
rect 7686 8862 7714 8890
rect 6454 8721 6482 8722
rect 6454 8695 6455 8721
rect 6455 8695 6481 8721
rect 6481 8695 6482 8721
rect 6454 8694 6482 8695
rect 6790 8694 6818 8722
rect 2238 8245 2266 8246
rect 2238 8219 2239 8245
rect 2239 8219 2265 8245
rect 2265 8219 2266 8245
rect 2238 8218 2266 8219
rect 2290 8245 2318 8246
rect 2290 8219 2291 8245
rect 2291 8219 2317 8245
rect 2317 8219 2318 8245
rect 2290 8218 2318 8219
rect 2342 8245 2370 8246
rect 2342 8219 2343 8245
rect 2343 8219 2369 8245
rect 2369 8219 2370 8245
rect 2342 8218 2370 8219
rect 5950 7713 5978 7714
rect 5950 7687 5951 7713
rect 5951 7687 5977 7713
rect 5977 7687 5978 7713
rect 5950 7686 5978 7687
rect 5614 7574 5642 7602
rect 6790 7574 6818 7602
rect 2238 7461 2266 7462
rect 2238 7435 2239 7461
rect 2239 7435 2265 7461
rect 2265 7435 2266 7461
rect 2238 7434 2266 7435
rect 2290 7461 2318 7462
rect 2290 7435 2291 7461
rect 2291 7435 2317 7461
rect 2317 7435 2318 7461
rect 2290 7434 2318 7435
rect 2342 7461 2370 7462
rect 2342 7435 2343 7461
rect 2343 7435 2369 7461
rect 2369 7435 2370 7461
rect 2342 7434 2370 7435
rect 7126 8777 7154 8778
rect 7126 8751 7127 8777
rect 7127 8751 7153 8777
rect 7153 8751 7154 8777
rect 7126 8750 7154 8751
rect 7182 8694 7210 8722
rect 6958 8470 6986 8498
rect 7406 8441 7434 8442
rect 7406 8415 7407 8441
rect 7407 8415 7433 8441
rect 7433 8415 7434 8441
rect 7406 8414 7434 8415
rect 7630 8441 7658 8442
rect 7630 8415 7631 8441
rect 7631 8415 7657 8441
rect 7657 8415 7658 8441
rect 7630 8414 7658 8415
rect 8022 10681 8050 10682
rect 8022 10655 8023 10681
rect 8023 10655 8049 10681
rect 8049 10655 8050 10681
rect 8022 10654 8050 10655
rect 8078 10094 8106 10122
rect 8022 10065 8050 10066
rect 8022 10039 8023 10065
rect 8023 10039 8049 10065
rect 8049 10039 8050 10065
rect 8022 10038 8050 10039
rect 7966 10009 7994 10010
rect 7966 9983 7967 10009
rect 7967 9983 7993 10009
rect 7993 9983 7994 10009
rect 7966 9982 7994 9983
rect 7910 9673 7938 9674
rect 7910 9647 7911 9673
rect 7911 9647 7937 9673
rect 7937 9647 7938 9673
rect 7910 9646 7938 9647
rect 7910 9366 7938 9394
rect 8358 10542 8386 10570
rect 8246 9982 8274 10010
rect 8358 9590 8386 9618
rect 8470 9814 8498 9842
rect 8246 9534 8274 9562
rect 7966 9086 7994 9114
rect 8078 9198 8106 9226
rect 8078 8974 8106 9002
rect 8190 9225 8218 9226
rect 8190 9199 8191 9225
rect 8191 9199 8217 9225
rect 8217 9199 8218 9225
rect 8190 9198 8218 9199
rect 7742 8806 7770 8834
rect 7910 8694 7938 8722
rect 7910 8497 7938 8498
rect 7910 8471 7911 8497
rect 7911 8471 7937 8497
rect 7937 8471 7938 8497
rect 7910 8470 7938 8471
rect 7630 8105 7658 8106
rect 7630 8079 7631 8105
rect 7631 8079 7657 8105
rect 7657 8079 7658 8105
rect 7630 8078 7658 8079
rect 7854 8414 7882 8442
rect 8078 8441 8106 8442
rect 8078 8415 8079 8441
rect 8079 8415 8105 8441
rect 8105 8415 8106 8441
rect 8078 8414 8106 8415
rect 8190 8470 8218 8498
rect 8806 10094 8834 10122
rect 8750 10038 8778 10066
rect 8638 9982 8666 10010
rect 8638 9478 8666 9506
rect 8862 9814 8890 9842
rect 8750 9534 8778 9562
rect 8974 10262 9002 10290
rect 8806 9310 8834 9338
rect 9030 10009 9058 10010
rect 9030 9983 9031 10009
rect 9031 9983 9057 10009
rect 9057 9983 9058 10009
rect 9030 9982 9058 9983
rect 9030 9561 9058 9562
rect 9030 9535 9031 9561
rect 9031 9535 9057 9561
rect 9057 9535 9058 9561
rect 9030 9534 9058 9535
rect 9254 11129 9282 11130
rect 9254 11103 9255 11129
rect 9255 11103 9281 11129
rect 9281 11103 9282 11129
rect 9254 11102 9282 11103
rect 9422 12473 9450 12474
rect 9422 12447 9423 12473
rect 9423 12447 9449 12473
rect 9449 12447 9450 12473
rect 9422 12446 9450 12447
rect 10318 13398 10346 13426
rect 10710 18745 10738 18746
rect 10710 18719 10711 18745
rect 10711 18719 10737 18745
rect 10737 18719 10738 18745
rect 10710 18718 10738 18719
rect 11718 14126 11746 14154
rect 11158 13566 11186 13594
rect 10374 13230 10402 13258
rect 11102 13510 11130 13538
rect 11158 13481 11186 13482
rect 11158 13455 11159 13481
rect 11159 13455 11185 13481
rect 11185 13455 11186 13481
rect 11158 13454 11186 13455
rect 11382 13454 11410 13482
rect 17598 19221 17626 19222
rect 17598 19195 17599 19221
rect 17599 19195 17625 19221
rect 17625 19195 17626 19221
rect 17598 19194 17626 19195
rect 17650 19221 17678 19222
rect 17650 19195 17651 19221
rect 17651 19195 17677 19221
rect 17677 19195 17678 19221
rect 17650 19194 17678 19195
rect 17702 19221 17730 19222
rect 17702 19195 17703 19221
rect 17703 19195 17729 19221
rect 17729 19195 17730 19221
rect 17702 19194 17730 19195
rect 12278 14126 12306 14154
rect 20118 18494 20146 18522
rect 17598 18437 17626 18438
rect 17598 18411 17599 18437
rect 17599 18411 17625 18437
rect 17625 18411 17626 18437
rect 17598 18410 17626 18411
rect 17650 18437 17678 18438
rect 17650 18411 17651 18437
rect 17651 18411 17677 18437
rect 17677 18411 17678 18437
rect 17650 18410 17678 18411
rect 17702 18437 17730 18438
rect 17702 18411 17703 18437
rect 17703 18411 17729 18437
rect 17729 18411 17730 18437
rect 17702 18410 17730 18411
rect 17598 17653 17626 17654
rect 17598 17627 17599 17653
rect 17599 17627 17625 17653
rect 17625 17627 17626 17653
rect 17598 17626 17626 17627
rect 17650 17653 17678 17654
rect 17650 17627 17651 17653
rect 17651 17627 17677 17653
rect 17677 17627 17678 17653
rect 17650 17626 17678 17627
rect 17702 17653 17730 17654
rect 17702 17627 17703 17653
rect 17703 17627 17729 17653
rect 17729 17627 17730 17653
rect 17702 17626 17730 17627
rect 20118 17150 20146 17178
rect 17598 16869 17626 16870
rect 17598 16843 17599 16869
rect 17599 16843 17625 16869
rect 17625 16843 17626 16869
rect 17598 16842 17626 16843
rect 17650 16869 17678 16870
rect 17650 16843 17651 16869
rect 17651 16843 17677 16869
rect 17677 16843 17678 16869
rect 17650 16842 17678 16843
rect 17702 16869 17730 16870
rect 17702 16843 17703 16869
rect 17703 16843 17729 16869
rect 17729 16843 17730 16869
rect 17702 16842 17730 16843
rect 17598 16085 17626 16086
rect 17598 16059 17599 16085
rect 17599 16059 17625 16085
rect 17625 16059 17626 16085
rect 17598 16058 17626 16059
rect 17650 16085 17678 16086
rect 17650 16059 17651 16085
rect 17651 16059 17677 16085
rect 17677 16059 17678 16085
rect 17650 16058 17678 16059
rect 17702 16085 17730 16086
rect 17702 16059 17703 16085
rect 17703 16059 17729 16085
rect 17729 16059 17730 16085
rect 17702 16058 17730 16059
rect 17598 15301 17626 15302
rect 17598 15275 17599 15301
rect 17599 15275 17625 15301
rect 17625 15275 17626 15301
rect 17598 15274 17626 15275
rect 17650 15301 17678 15302
rect 17650 15275 17651 15301
rect 17651 15275 17677 15301
rect 17677 15275 17678 15301
rect 17650 15274 17678 15275
rect 17702 15301 17730 15302
rect 17702 15275 17703 15301
rect 17703 15275 17729 15301
rect 17729 15275 17730 15301
rect 17702 15274 17730 15275
rect 17598 14517 17626 14518
rect 17598 14491 17599 14517
rect 17599 14491 17625 14517
rect 17625 14491 17626 14517
rect 17598 14490 17626 14491
rect 17650 14517 17678 14518
rect 17650 14491 17651 14517
rect 17651 14491 17677 14517
rect 17677 14491 17678 14517
rect 17650 14490 17678 14491
rect 17702 14517 17730 14518
rect 17702 14491 17703 14517
rect 17703 14491 17729 14517
rect 17729 14491 17730 14517
rect 17702 14490 17730 14491
rect 11662 13510 11690 13538
rect 10766 13230 10794 13258
rect 10374 12809 10402 12810
rect 10374 12783 10375 12809
rect 10375 12783 10401 12809
rect 10401 12783 10402 12809
rect 10374 12782 10402 12783
rect 10150 12753 10178 12754
rect 10150 12727 10151 12753
rect 10151 12727 10177 12753
rect 10177 12727 10178 12753
rect 10150 12726 10178 12727
rect 10318 12726 10346 12754
rect 9366 10822 9394 10850
rect 10038 12641 10066 12642
rect 10038 12615 10039 12641
rect 10039 12615 10065 12641
rect 10065 12615 10066 12641
rect 10038 12614 10066 12615
rect 9918 12557 9946 12558
rect 9918 12531 9919 12557
rect 9919 12531 9945 12557
rect 9945 12531 9946 12557
rect 9918 12530 9946 12531
rect 9970 12557 9998 12558
rect 9970 12531 9971 12557
rect 9971 12531 9997 12557
rect 9997 12531 9998 12557
rect 9970 12530 9998 12531
rect 10022 12557 10050 12558
rect 10022 12531 10023 12557
rect 10023 12531 10049 12557
rect 10049 12531 10050 12557
rect 10022 12530 10050 12531
rect 9814 12361 9842 12362
rect 9814 12335 9815 12361
rect 9815 12335 9841 12361
rect 9841 12335 9842 12361
rect 9814 12334 9842 12335
rect 9590 11606 9618 11634
rect 9918 11773 9946 11774
rect 9918 11747 9919 11773
rect 9919 11747 9945 11773
rect 9945 11747 9946 11773
rect 9918 11746 9946 11747
rect 9970 11773 9998 11774
rect 9970 11747 9971 11773
rect 9971 11747 9997 11773
rect 9997 11747 9998 11773
rect 9970 11746 9998 11747
rect 10022 11773 10050 11774
rect 10022 11747 10023 11773
rect 10023 11747 10049 11773
rect 10049 11747 10050 11773
rect 10022 11746 10050 11747
rect 11998 13510 12026 13538
rect 12894 13537 12922 13538
rect 12894 13511 12895 13537
rect 12895 13511 12921 13537
rect 12921 13511 12922 13537
rect 12894 13510 12922 13511
rect 12222 13454 12250 13482
rect 11942 12726 11970 12754
rect 17598 13733 17626 13734
rect 17598 13707 17599 13733
rect 17599 13707 17625 13733
rect 17625 13707 17626 13733
rect 17598 13706 17626 13707
rect 17650 13733 17678 13734
rect 17650 13707 17651 13733
rect 17651 13707 17677 13733
rect 17677 13707 17678 13733
rect 17650 13706 17678 13707
rect 17702 13733 17730 13734
rect 17702 13707 17703 13733
rect 17703 13707 17729 13733
rect 17729 13707 17730 13733
rect 17702 13706 17730 13707
rect 13062 13566 13090 13594
rect 13342 13566 13370 13594
rect 13398 13481 13426 13482
rect 13398 13455 13399 13481
rect 13399 13455 13425 13481
rect 13425 13455 13426 13481
rect 13398 13454 13426 13455
rect 14630 13454 14658 13482
rect 10990 12641 11018 12642
rect 10990 12615 10991 12641
rect 10991 12615 11017 12641
rect 11017 12615 11018 12641
rect 10990 12614 11018 12615
rect 12110 12614 12138 12642
rect 12726 12614 12754 12642
rect 12390 12334 12418 12362
rect 10206 11689 10234 11690
rect 10206 11663 10207 11689
rect 10207 11663 10233 11689
rect 10233 11663 10234 11689
rect 10206 11662 10234 11663
rect 9646 11326 9674 11354
rect 10038 11326 10066 11354
rect 9534 10878 9562 10906
rect 9702 10878 9730 10906
rect 9870 11046 9898 11074
rect 9918 10989 9946 10990
rect 9918 10963 9919 10989
rect 9919 10963 9945 10989
rect 9945 10963 9946 10989
rect 9918 10962 9946 10963
rect 9970 10989 9998 10990
rect 9970 10963 9971 10989
rect 9971 10963 9997 10989
rect 9997 10963 9998 10989
rect 9970 10962 9998 10963
rect 10022 10989 10050 10990
rect 10022 10963 10023 10989
rect 10023 10963 10049 10989
rect 10049 10963 10050 10989
rect 10022 10962 10050 10963
rect 9310 10737 9338 10738
rect 9310 10711 9311 10737
rect 9311 10711 9337 10737
rect 9337 10711 9338 10737
rect 9310 10710 9338 10711
rect 9198 10038 9226 10066
rect 9142 9870 9170 9898
rect 8470 9254 8498 9282
rect 8806 9225 8834 9226
rect 8806 9199 8807 9225
rect 8807 9199 8833 9225
rect 8833 9199 8834 9225
rect 8806 9198 8834 9199
rect 8638 9030 8666 9058
rect 8694 9086 8722 9114
rect 8302 8862 8330 8890
rect 8526 8833 8554 8834
rect 8526 8807 8527 8833
rect 8527 8807 8553 8833
rect 8553 8807 8554 8833
rect 8526 8806 8554 8807
rect 8190 8358 8218 8386
rect 7686 7686 7714 7714
rect 8414 8358 8442 8386
rect 8246 8078 8274 8106
rect 8862 8441 8890 8442
rect 8862 8415 8863 8441
rect 8863 8415 8889 8441
rect 8889 8415 8890 8441
rect 8862 8414 8890 8415
rect 8974 9225 9002 9226
rect 8974 9199 8975 9225
rect 8975 9199 9001 9225
rect 9001 9199 9002 9225
rect 8974 9198 9002 9199
rect 8918 8358 8946 8386
rect 8638 7238 8666 7266
rect 7406 7126 7434 7154
rect 7742 7126 7770 7154
rect 2238 6677 2266 6678
rect 2238 6651 2239 6677
rect 2239 6651 2265 6677
rect 2265 6651 2266 6677
rect 2238 6650 2266 6651
rect 2290 6677 2318 6678
rect 2290 6651 2291 6677
rect 2291 6651 2317 6677
rect 2317 6651 2318 6677
rect 2290 6650 2318 6651
rect 2342 6677 2370 6678
rect 2342 6651 2343 6677
rect 2343 6651 2369 6677
rect 2369 6651 2370 6677
rect 2342 6650 2370 6651
rect 8414 7153 8442 7154
rect 8414 7127 8415 7153
rect 8415 7127 8441 7153
rect 8441 7127 8442 7153
rect 8414 7126 8442 7127
rect 8974 7153 9002 7154
rect 8974 7127 8975 7153
rect 8975 7127 9001 7153
rect 9001 7127 9002 7153
rect 8974 7126 9002 7127
rect 8414 6873 8442 6874
rect 8414 6847 8415 6873
rect 8415 6847 8441 6873
rect 8441 6847 8442 6873
rect 8414 6846 8442 6847
rect 8750 6873 8778 6874
rect 8750 6847 8751 6873
rect 8751 6847 8777 6873
rect 8777 6847 8778 6873
rect 8750 6846 8778 6847
rect 8918 6873 8946 6874
rect 8918 6847 8919 6873
rect 8919 6847 8945 6873
rect 8945 6847 8946 6873
rect 8918 6846 8946 6847
rect 9086 9198 9114 9226
rect 9870 10766 9898 10794
rect 10038 10822 10066 10850
rect 10038 10401 10066 10402
rect 10038 10375 10039 10401
rect 10039 10375 10065 10401
rect 10065 10375 10066 10401
rect 10038 10374 10066 10375
rect 9926 10262 9954 10290
rect 9918 10205 9946 10206
rect 9918 10179 9919 10205
rect 9919 10179 9945 10205
rect 9945 10179 9946 10205
rect 9918 10178 9946 10179
rect 9970 10205 9998 10206
rect 9970 10179 9971 10205
rect 9971 10179 9997 10205
rect 9997 10179 9998 10205
rect 9970 10178 9998 10179
rect 10022 10205 10050 10206
rect 10022 10179 10023 10205
rect 10023 10179 10049 10205
rect 10049 10179 10050 10205
rect 10022 10178 10050 10179
rect 9702 10094 9730 10122
rect 9702 9982 9730 10010
rect 9254 9702 9282 9730
rect 9422 9617 9450 9618
rect 9422 9591 9423 9617
rect 9423 9591 9449 9617
rect 9449 9591 9450 9617
rect 9422 9590 9450 9591
rect 9702 9590 9730 9618
rect 9254 9366 9282 9394
rect 9254 9254 9282 9282
rect 9310 9169 9338 9170
rect 9310 9143 9311 9169
rect 9311 9143 9337 9169
rect 9337 9143 9338 9169
rect 9310 9142 9338 9143
rect 9422 9142 9450 9170
rect 9198 9086 9226 9114
rect 9254 8833 9282 8834
rect 9254 8807 9255 8833
rect 9255 8807 9281 8833
rect 9281 8807 9282 8833
rect 9254 8806 9282 8807
rect 9590 9225 9618 9226
rect 9590 9199 9591 9225
rect 9591 9199 9617 9225
rect 9617 9199 9618 9225
rect 9590 9198 9618 9199
rect 9870 9617 9898 9618
rect 9870 9591 9871 9617
rect 9871 9591 9897 9617
rect 9897 9591 9898 9617
rect 9870 9590 9898 9591
rect 9918 9421 9946 9422
rect 9918 9395 9919 9421
rect 9919 9395 9945 9421
rect 9945 9395 9946 9421
rect 9918 9394 9946 9395
rect 9970 9421 9998 9422
rect 9970 9395 9971 9421
rect 9971 9395 9997 9421
rect 9997 9395 9998 9421
rect 9970 9394 9998 9395
rect 10022 9421 10050 9422
rect 10022 9395 10023 9421
rect 10023 9395 10049 9421
rect 10049 9395 10050 9421
rect 10022 9394 10050 9395
rect 9982 9310 10010 9338
rect 9478 8414 9506 8442
rect 9646 8414 9674 8442
rect 9534 8358 9562 8386
rect 9478 8246 9506 8274
rect 11494 11214 11522 11242
rect 10318 11073 10346 11074
rect 10318 11047 10319 11073
rect 10319 11047 10345 11073
rect 10345 11047 10346 11073
rect 10318 11046 10346 11047
rect 10822 10934 10850 10962
rect 10262 10878 10290 10906
rect 11494 11046 11522 11074
rect 11886 10905 11914 10906
rect 11886 10879 11887 10905
rect 11887 10879 11913 10905
rect 11913 10879 11914 10905
rect 11886 10878 11914 10879
rect 10206 10486 10234 10514
rect 10206 10038 10234 10066
rect 10318 10710 10346 10738
rect 10430 10542 10458 10570
rect 10542 10486 10570 10514
rect 10486 10430 10514 10458
rect 10710 10793 10738 10794
rect 10710 10767 10711 10793
rect 10711 10767 10737 10793
rect 10737 10767 10738 10793
rect 10710 10766 10738 10767
rect 10822 10710 10850 10738
rect 10822 10486 10850 10514
rect 10934 10542 10962 10570
rect 10878 10430 10906 10458
rect 10654 9982 10682 10010
rect 10318 9590 10346 9618
rect 10654 9758 10682 9786
rect 10374 9366 10402 9394
rect 10486 9478 10514 9506
rect 10262 9310 10290 9338
rect 10374 9254 10402 9282
rect 10094 9142 10122 9170
rect 9870 8918 9898 8946
rect 9982 8833 10010 8834
rect 9982 8807 9983 8833
rect 9983 8807 10009 8833
rect 10009 8807 10010 8833
rect 9982 8806 10010 8807
rect 9702 8358 9730 8386
rect 9918 8637 9946 8638
rect 9918 8611 9919 8637
rect 9919 8611 9945 8637
rect 9945 8611 9946 8637
rect 9918 8610 9946 8611
rect 9970 8637 9998 8638
rect 9970 8611 9971 8637
rect 9971 8611 9997 8637
rect 9997 8611 9998 8637
rect 9970 8610 9998 8611
rect 10022 8637 10050 8638
rect 10022 8611 10023 8637
rect 10023 8611 10049 8637
rect 10049 8611 10050 8637
rect 10022 8610 10050 8611
rect 10822 9617 10850 9618
rect 10822 9591 10823 9617
rect 10823 9591 10849 9617
rect 10849 9591 10850 9617
rect 10822 9590 10850 9591
rect 11774 10849 11802 10850
rect 11774 10823 11775 10849
rect 11775 10823 11801 10849
rect 11801 10823 11802 10849
rect 11774 10822 11802 10823
rect 11046 10766 11074 10794
rect 11270 10654 11298 10682
rect 11382 10710 11410 10738
rect 11438 10766 11466 10794
rect 11326 10598 11354 10626
rect 11158 10401 11186 10402
rect 11158 10375 11159 10401
rect 11159 10375 11185 10401
rect 11185 10375 11186 10401
rect 11158 10374 11186 10375
rect 10990 9926 11018 9954
rect 11326 9814 11354 9842
rect 11046 9366 11074 9394
rect 10654 9142 10682 9170
rect 10654 8974 10682 9002
rect 10150 8470 10178 8498
rect 10206 8441 10234 8442
rect 10206 8415 10207 8441
rect 10207 8415 10233 8441
rect 10233 8415 10234 8441
rect 10206 8414 10234 8415
rect 12110 11577 12138 11578
rect 12110 11551 12111 11577
rect 12111 11551 12137 11577
rect 12137 11551 12138 11577
rect 12110 11550 12138 11551
rect 12054 11158 12082 11186
rect 12166 11102 12194 11130
rect 11998 10905 12026 10906
rect 11998 10879 11999 10905
rect 11999 10879 12025 10905
rect 12025 10879 12026 10905
rect 11998 10878 12026 10879
rect 11942 10654 11970 10682
rect 11886 10430 11914 10458
rect 11438 9366 11466 9394
rect 11550 9337 11578 9338
rect 11550 9311 11551 9337
rect 11551 9311 11577 9337
rect 11577 9311 11578 9337
rect 11550 9310 11578 9311
rect 11774 9337 11802 9338
rect 11774 9311 11775 9337
rect 11775 9311 11801 9337
rect 11801 9311 11802 9337
rect 11774 9310 11802 9311
rect 11606 9198 11634 9226
rect 12222 10430 12250 10458
rect 12950 12838 12978 12866
rect 13510 12838 13538 12866
rect 18830 13230 18858 13258
rect 14966 13201 14994 13202
rect 14966 13175 14967 13201
rect 14967 13175 14993 13201
rect 14993 13175 14994 13201
rect 14966 13174 14994 13175
rect 18830 13145 18858 13146
rect 18830 13119 18831 13145
rect 18831 13119 18857 13145
rect 18857 13119 18858 13145
rect 18830 13118 18858 13119
rect 14798 13062 14826 13090
rect 17598 12949 17626 12950
rect 17598 12923 17599 12949
rect 17599 12923 17625 12949
rect 17625 12923 17626 12949
rect 17598 12922 17626 12923
rect 17650 12949 17678 12950
rect 17650 12923 17651 12949
rect 17651 12923 17677 12949
rect 17677 12923 17678 12949
rect 17650 12922 17678 12923
rect 17702 12949 17730 12950
rect 17702 12923 17703 12949
rect 17703 12923 17729 12949
rect 17729 12923 17730 12949
rect 17702 12922 17730 12923
rect 19950 13454 19978 13482
rect 20006 13118 20034 13146
rect 18942 12838 18970 12866
rect 20006 12782 20034 12810
rect 13174 12614 13202 12642
rect 13398 12614 13426 12642
rect 13230 11774 13258 11802
rect 12726 11633 12754 11634
rect 12726 11607 12727 11633
rect 12727 11607 12753 11633
rect 12753 11607 12754 11633
rect 12726 11606 12754 11607
rect 12334 10934 12362 10962
rect 12334 10793 12362 10794
rect 12334 10767 12335 10793
rect 12335 10767 12361 10793
rect 12361 10767 12362 10793
rect 12334 10766 12362 10767
rect 12390 10598 12418 10626
rect 12334 10150 12362 10178
rect 12278 9926 12306 9954
rect 12110 9337 12138 9338
rect 12110 9311 12111 9337
rect 12111 9311 12137 9337
rect 12137 9311 12138 9337
rect 12110 9310 12138 9311
rect 11102 9030 11130 9058
rect 10038 8358 10066 8386
rect 10766 8302 10794 8330
rect 10374 7910 10402 7938
rect 9918 7853 9946 7854
rect 9918 7827 9919 7853
rect 9919 7827 9945 7853
rect 9945 7827 9946 7853
rect 9918 7826 9946 7827
rect 9970 7853 9998 7854
rect 9970 7827 9971 7853
rect 9971 7827 9997 7853
rect 9997 7827 9998 7853
rect 9970 7826 9998 7827
rect 10022 7853 10050 7854
rect 10022 7827 10023 7853
rect 10023 7827 10049 7853
rect 10049 7827 10050 7853
rect 10022 7826 10050 7827
rect 9758 7686 9786 7714
rect 9814 7742 9842 7770
rect 9254 7518 9282 7546
rect 8974 6790 9002 6818
rect 9534 7518 9562 7546
rect 9646 7294 9674 7322
rect 9422 7265 9450 7266
rect 9422 7239 9423 7265
rect 9423 7239 9449 7265
rect 9449 7239 9450 7265
rect 9422 7238 9450 7239
rect 10038 7518 10066 7546
rect 11606 9086 11634 9114
rect 11326 7966 11354 7994
rect 11270 7937 11298 7938
rect 11270 7911 11271 7937
rect 11271 7911 11297 7937
rect 11297 7911 11298 7937
rect 11270 7910 11298 7911
rect 11550 8470 11578 8498
rect 11438 7937 11466 7938
rect 11438 7911 11439 7937
rect 11439 7911 11465 7937
rect 11465 7911 11466 7937
rect 11438 7910 11466 7911
rect 11382 7854 11410 7882
rect 10878 7630 10906 7658
rect 10486 7294 10514 7322
rect 10710 7574 10738 7602
rect 10374 7265 10402 7266
rect 10374 7239 10375 7265
rect 10375 7239 10401 7265
rect 10401 7239 10402 7265
rect 10374 7238 10402 7239
rect 11438 7630 11466 7658
rect 10710 7265 10738 7266
rect 10710 7239 10711 7265
rect 10711 7239 10737 7265
rect 10737 7239 10738 7265
rect 10710 7238 10738 7239
rect 11214 7238 11242 7266
rect 9926 7209 9954 7210
rect 9926 7183 9927 7209
rect 9927 7183 9953 7209
rect 9953 7183 9954 7209
rect 9926 7182 9954 7183
rect 10150 7153 10178 7154
rect 10150 7127 10151 7153
rect 10151 7127 10177 7153
rect 10177 7127 10178 7153
rect 10150 7126 10178 7127
rect 9918 7069 9946 7070
rect 9918 7043 9919 7069
rect 9919 7043 9945 7069
rect 9945 7043 9946 7069
rect 9918 7042 9946 7043
rect 9970 7069 9998 7070
rect 9970 7043 9971 7069
rect 9971 7043 9997 7069
rect 9997 7043 9998 7069
rect 9970 7042 9998 7043
rect 10022 7069 10050 7070
rect 10022 7043 10023 7069
rect 10023 7043 10049 7069
rect 10049 7043 10050 7069
rect 10022 7042 10050 7043
rect 9310 6846 9338 6874
rect 9254 6790 9282 6818
rect 9646 6790 9674 6818
rect 8806 6510 8834 6538
rect 2238 5893 2266 5894
rect 2238 5867 2239 5893
rect 2239 5867 2265 5893
rect 2265 5867 2266 5893
rect 2238 5866 2266 5867
rect 2290 5893 2318 5894
rect 2290 5867 2291 5893
rect 2291 5867 2317 5893
rect 2317 5867 2318 5893
rect 2290 5866 2318 5867
rect 2342 5893 2370 5894
rect 2342 5867 2343 5893
rect 2343 5867 2369 5893
rect 2369 5867 2370 5893
rect 2342 5866 2370 5867
rect 2238 5109 2266 5110
rect 2238 5083 2239 5109
rect 2239 5083 2265 5109
rect 2265 5083 2266 5109
rect 2238 5082 2266 5083
rect 2290 5109 2318 5110
rect 2290 5083 2291 5109
rect 2291 5083 2317 5109
rect 2317 5083 2318 5109
rect 2290 5082 2318 5083
rect 2342 5109 2370 5110
rect 2342 5083 2343 5109
rect 2343 5083 2369 5109
rect 2369 5083 2370 5109
rect 2342 5082 2370 5083
rect 2238 4325 2266 4326
rect 2238 4299 2239 4325
rect 2239 4299 2265 4325
rect 2265 4299 2266 4325
rect 2238 4298 2266 4299
rect 2290 4325 2318 4326
rect 2290 4299 2291 4325
rect 2291 4299 2317 4325
rect 2317 4299 2318 4325
rect 2290 4298 2318 4299
rect 2342 4325 2370 4326
rect 2342 4299 2343 4325
rect 2343 4299 2369 4325
rect 2369 4299 2370 4325
rect 2342 4298 2370 4299
rect 2238 3541 2266 3542
rect 2238 3515 2239 3541
rect 2239 3515 2265 3541
rect 2265 3515 2266 3541
rect 2238 3514 2266 3515
rect 2290 3541 2318 3542
rect 2290 3515 2291 3541
rect 2291 3515 2317 3541
rect 2317 3515 2318 3541
rect 2290 3514 2318 3515
rect 2342 3541 2370 3542
rect 2342 3515 2343 3541
rect 2343 3515 2369 3541
rect 2369 3515 2370 3541
rect 2342 3514 2370 3515
rect 2238 2757 2266 2758
rect 2238 2731 2239 2757
rect 2239 2731 2265 2757
rect 2265 2731 2266 2757
rect 2238 2730 2266 2731
rect 2290 2757 2318 2758
rect 2290 2731 2291 2757
rect 2291 2731 2317 2757
rect 2317 2731 2318 2757
rect 2290 2730 2318 2731
rect 2342 2757 2370 2758
rect 2342 2731 2343 2757
rect 2343 2731 2369 2757
rect 2369 2731 2370 2757
rect 2342 2730 2370 2731
rect 2238 1973 2266 1974
rect 2238 1947 2239 1973
rect 2239 1947 2265 1973
rect 2265 1947 2266 1973
rect 2238 1946 2266 1947
rect 2290 1973 2318 1974
rect 2290 1947 2291 1973
rect 2291 1947 2317 1973
rect 2317 1947 2318 1973
rect 2290 1946 2318 1947
rect 2342 1973 2370 1974
rect 2342 1947 2343 1973
rect 2343 1947 2369 1973
rect 2369 1947 2370 1973
rect 2342 1946 2370 1947
rect 9142 6537 9170 6538
rect 9142 6511 9143 6537
rect 9143 6511 9169 6537
rect 9169 6511 9170 6537
rect 9142 6510 9170 6511
rect 9366 6537 9394 6538
rect 9366 6511 9367 6537
rect 9367 6511 9393 6537
rect 9393 6511 9394 6537
rect 9366 6510 9394 6511
rect 9918 6285 9946 6286
rect 9918 6259 9919 6285
rect 9919 6259 9945 6285
rect 9945 6259 9946 6285
rect 9918 6258 9946 6259
rect 9970 6285 9998 6286
rect 9970 6259 9971 6285
rect 9971 6259 9997 6285
rect 9997 6259 9998 6285
rect 9970 6258 9998 6259
rect 10022 6285 10050 6286
rect 10022 6259 10023 6285
rect 10023 6259 10049 6285
rect 10049 6259 10050 6285
rect 10022 6258 10050 6259
rect 9918 5501 9946 5502
rect 9918 5475 9919 5501
rect 9919 5475 9945 5501
rect 9945 5475 9946 5501
rect 9918 5474 9946 5475
rect 9970 5501 9998 5502
rect 9970 5475 9971 5501
rect 9971 5475 9997 5501
rect 9997 5475 9998 5501
rect 9970 5474 9998 5475
rect 10022 5501 10050 5502
rect 10022 5475 10023 5501
rect 10023 5475 10049 5501
rect 10049 5475 10050 5501
rect 10022 5474 10050 5475
rect 9918 4717 9946 4718
rect 9918 4691 9919 4717
rect 9919 4691 9945 4717
rect 9945 4691 9946 4717
rect 9918 4690 9946 4691
rect 9970 4717 9998 4718
rect 9970 4691 9971 4717
rect 9971 4691 9997 4717
rect 9997 4691 9998 4717
rect 9970 4690 9998 4691
rect 10022 4717 10050 4718
rect 10022 4691 10023 4717
rect 10023 4691 10049 4717
rect 10049 4691 10050 4717
rect 10022 4690 10050 4691
rect 12222 9702 12250 9730
rect 12390 10094 12418 10122
rect 12502 9982 12530 10010
rect 12502 9366 12530 9394
rect 12614 11550 12642 11578
rect 12782 11577 12810 11578
rect 12782 11551 12783 11577
rect 12783 11551 12809 11577
rect 12809 11551 12810 11577
rect 12782 11550 12810 11551
rect 12838 11214 12866 11242
rect 12670 10990 12698 11018
rect 12782 11073 12810 11074
rect 12782 11047 12783 11073
rect 12783 11047 12809 11073
rect 12809 11047 12810 11073
rect 12782 11046 12810 11047
rect 12782 10934 12810 10962
rect 12614 10710 12642 10738
rect 12726 10598 12754 10626
rect 12614 10094 12642 10122
rect 12726 10486 12754 10514
rect 12782 10150 12810 10178
rect 12894 11185 12922 11186
rect 12894 11159 12895 11185
rect 12895 11159 12921 11185
rect 12921 11159 12922 11185
rect 12894 11158 12922 11159
rect 12950 10878 12978 10906
rect 13006 11662 13034 11690
rect 12894 10849 12922 10850
rect 12894 10823 12895 10849
rect 12895 10823 12921 10849
rect 12921 10823 12922 10849
rect 12894 10822 12922 10823
rect 14014 12641 14042 12642
rect 14014 12615 14015 12641
rect 14015 12615 14041 12641
rect 14041 12615 14042 12641
rect 14014 12614 14042 12615
rect 17598 12165 17626 12166
rect 17598 12139 17599 12165
rect 17599 12139 17625 12165
rect 17625 12139 17626 12165
rect 17598 12138 17626 12139
rect 17650 12165 17678 12166
rect 17650 12139 17651 12165
rect 17651 12139 17677 12165
rect 17677 12139 17678 12165
rect 17650 12138 17678 12139
rect 17702 12165 17730 12166
rect 17702 12139 17703 12165
rect 17703 12139 17729 12165
rect 17729 12139 17730 12165
rect 17702 12138 17730 12139
rect 13734 11774 13762 11802
rect 13398 11662 13426 11690
rect 14630 11689 14658 11690
rect 14630 11663 14631 11689
rect 14631 11663 14657 11689
rect 14657 11663 14658 11689
rect 14630 11662 14658 11663
rect 18830 11577 18858 11578
rect 18830 11551 18831 11577
rect 18831 11551 18857 11577
rect 18857 11551 18858 11577
rect 18830 11550 18858 11551
rect 13062 11073 13090 11074
rect 13062 11047 13063 11073
rect 13063 11047 13089 11073
rect 13089 11047 13090 11073
rect 13062 11046 13090 11047
rect 12950 10766 12978 10794
rect 14406 11521 14434 11522
rect 14406 11495 14407 11521
rect 14407 11495 14433 11521
rect 14433 11495 14434 11521
rect 14406 11494 14434 11495
rect 20006 11465 20034 11466
rect 20006 11439 20007 11465
rect 20007 11439 20033 11465
rect 20033 11439 20034 11465
rect 20006 11438 20034 11439
rect 17598 11381 17626 11382
rect 17598 11355 17599 11381
rect 17599 11355 17625 11381
rect 17625 11355 17626 11381
rect 17598 11354 17626 11355
rect 17650 11381 17678 11382
rect 17650 11355 17651 11381
rect 17651 11355 17677 11381
rect 17677 11355 17678 11381
rect 17650 11354 17678 11355
rect 17702 11381 17730 11382
rect 17702 11355 17703 11381
rect 17703 11355 17729 11381
rect 17729 11355 17730 11381
rect 17702 11354 17730 11355
rect 13342 11241 13370 11242
rect 13342 11215 13343 11241
rect 13343 11215 13369 11241
rect 13369 11215 13370 11241
rect 13342 11214 13370 11215
rect 13790 11185 13818 11186
rect 13790 11159 13791 11185
rect 13791 11159 13817 11185
rect 13817 11159 13818 11185
rect 13790 11158 13818 11159
rect 13286 10934 13314 10962
rect 13230 10486 13258 10514
rect 13342 10793 13370 10794
rect 13342 10767 13343 10793
rect 13343 10767 13369 10793
rect 13369 10767 13370 10793
rect 13342 10766 13370 10767
rect 13006 10121 13034 10122
rect 13006 10095 13007 10121
rect 13007 10095 13033 10121
rect 13033 10095 13034 10121
rect 13006 10094 13034 10095
rect 13622 10990 13650 11018
rect 14742 10766 14770 10794
rect 20006 11102 20034 11130
rect 18830 10766 18858 10794
rect 17598 10597 17626 10598
rect 17598 10571 17599 10597
rect 17599 10571 17625 10597
rect 17625 10571 17626 10597
rect 17598 10570 17626 10571
rect 17650 10597 17678 10598
rect 17650 10571 17651 10597
rect 17651 10571 17677 10597
rect 17677 10571 17678 10597
rect 17650 10570 17678 10571
rect 17702 10597 17730 10598
rect 17702 10571 17703 10597
rect 17703 10571 17729 10597
rect 17729 10571 17730 10597
rect 17702 10570 17730 10571
rect 13510 10094 13538 10122
rect 13118 10009 13146 10010
rect 13118 9983 13119 10009
rect 13119 9983 13145 10009
rect 13145 9983 13146 10009
rect 13118 9982 13146 9983
rect 13286 9982 13314 10010
rect 12614 9758 12642 9786
rect 12278 9086 12306 9114
rect 12166 8806 12194 8834
rect 12614 8246 12642 8274
rect 12670 8358 12698 8386
rect 12334 8022 12362 8050
rect 11662 7966 11690 7994
rect 11830 7910 11858 7938
rect 12110 7910 12138 7938
rect 11998 7854 12026 7882
rect 11830 7742 11858 7770
rect 11550 6873 11578 6874
rect 11550 6847 11551 6873
rect 11551 6847 11577 6873
rect 11577 6847 11578 6873
rect 11550 6846 11578 6847
rect 11998 7713 12026 7714
rect 11998 7687 11999 7713
rect 11999 7687 12025 7713
rect 12025 7687 12026 7713
rect 11998 7686 12026 7687
rect 12222 7798 12250 7826
rect 12334 7742 12362 7770
rect 12726 8049 12754 8050
rect 12726 8023 12727 8049
rect 12727 8023 12753 8049
rect 12753 8023 12754 8049
rect 12726 8022 12754 8023
rect 13062 9870 13090 9898
rect 13342 9926 13370 9954
rect 13958 9953 13986 9954
rect 13958 9927 13959 9953
rect 13959 9927 13985 9953
rect 13985 9927 13986 9953
rect 13958 9926 13986 9927
rect 14686 9926 14714 9954
rect 13398 9870 13426 9898
rect 15022 9953 15050 9954
rect 15022 9927 15023 9953
rect 15023 9927 15049 9953
rect 15049 9927 15050 9953
rect 15022 9926 15050 9927
rect 18830 9926 18858 9954
rect 17598 9813 17626 9814
rect 17598 9787 17599 9813
rect 17599 9787 17625 9813
rect 17625 9787 17626 9813
rect 17598 9786 17626 9787
rect 17650 9813 17678 9814
rect 17650 9787 17651 9813
rect 17651 9787 17677 9813
rect 17677 9787 17678 9813
rect 17650 9786 17678 9787
rect 17702 9813 17730 9814
rect 17702 9787 17703 9813
rect 17703 9787 17729 9813
rect 17729 9787 17730 9813
rect 17702 9786 17730 9787
rect 14070 9617 14098 9618
rect 14070 9591 14071 9617
rect 14071 9591 14097 9617
rect 14097 9591 14098 9617
rect 14070 9590 14098 9591
rect 14630 9617 14658 9618
rect 14630 9591 14631 9617
rect 14631 9591 14657 9617
rect 14657 9591 14658 9617
rect 14630 9590 14658 9591
rect 13174 9142 13202 9170
rect 13062 9030 13090 9058
rect 13174 8833 13202 8834
rect 13174 8807 13175 8833
rect 13175 8807 13201 8833
rect 13201 8807 13202 8833
rect 13174 8806 13202 8807
rect 12950 8358 12978 8386
rect 13622 9505 13650 9506
rect 13622 9479 13623 9505
rect 13623 9479 13649 9505
rect 13649 9479 13650 9505
rect 13622 9478 13650 9479
rect 13286 8833 13314 8834
rect 13286 8807 13287 8833
rect 13287 8807 13313 8833
rect 13313 8807 13314 8833
rect 13286 8806 13314 8807
rect 13230 8302 13258 8330
rect 13006 8246 13034 8274
rect 13286 8246 13314 8274
rect 20006 9422 20034 9450
rect 18830 9225 18858 9226
rect 18830 9199 18831 9225
rect 18831 9199 18857 9225
rect 18857 9199 18858 9225
rect 18830 9198 18858 9199
rect 13790 9142 13818 9170
rect 13958 9142 13986 9170
rect 13846 8833 13874 8834
rect 13846 8807 13847 8833
rect 13847 8807 13873 8833
rect 13873 8807 13874 8833
rect 13846 8806 13874 8807
rect 14574 9169 14602 9170
rect 14574 9143 14575 9169
rect 14575 9143 14601 9169
rect 14601 9143 14602 9169
rect 14574 9142 14602 9143
rect 20006 9113 20034 9114
rect 20006 9087 20007 9113
rect 20007 9087 20033 9113
rect 20033 9087 20034 9113
rect 20006 9086 20034 9087
rect 17598 9029 17626 9030
rect 17598 9003 17599 9029
rect 17599 9003 17625 9029
rect 17625 9003 17626 9029
rect 17598 9002 17626 9003
rect 17650 9029 17678 9030
rect 17650 9003 17651 9029
rect 17651 9003 17677 9029
rect 17677 9003 17678 9029
rect 17650 9002 17678 9003
rect 17702 9029 17730 9030
rect 17702 9003 17703 9029
rect 17703 9003 17729 9029
rect 17729 9003 17730 9029
rect 17702 9002 17730 9003
rect 13342 8022 13370 8050
rect 14462 8358 14490 8386
rect 13286 7966 13314 7994
rect 13566 7993 13594 7994
rect 13566 7967 13567 7993
rect 13567 7967 13593 7993
rect 13593 7967 13594 7993
rect 13566 7966 13594 7967
rect 13790 7993 13818 7994
rect 13790 7967 13791 7993
rect 13791 7967 13817 7993
rect 13817 7967 13818 7993
rect 13790 7966 13818 7967
rect 12782 7798 12810 7826
rect 12670 7574 12698 7602
rect 12166 7294 12194 7322
rect 12334 7265 12362 7266
rect 12334 7239 12335 7265
rect 12335 7239 12361 7265
rect 12361 7239 12362 7265
rect 12334 7238 12362 7239
rect 13398 7937 13426 7938
rect 13398 7911 13399 7937
rect 13399 7911 13425 7937
rect 13425 7911 13426 7937
rect 13398 7910 13426 7911
rect 13510 7854 13538 7882
rect 14070 7854 14098 7882
rect 13230 7574 13258 7602
rect 13006 7321 13034 7322
rect 13006 7295 13007 7321
rect 13007 7295 13033 7321
rect 13033 7295 13034 7321
rect 13006 7294 13034 7295
rect 14238 7601 14266 7602
rect 14238 7575 14239 7601
rect 14239 7575 14265 7601
rect 14265 7575 14266 7601
rect 14238 7574 14266 7575
rect 17598 8245 17626 8246
rect 17598 8219 17599 8245
rect 17599 8219 17625 8245
rect 17625 8219 17626 8245
rect 17598 8218 17626 8219
rect 17650 8245 17678 8246
rect 17650 8219 17651 8245
rect 17651 8219 17677 8245
rect 17677 8219 17678 8245
rect 17650 8218 17678 8219
rect 17702 8245 17730 8246
rect 17702 8219 17703 8245
rect 17703 8219 17729 8245
rect 17729 8219 17730 8245
rect 17702 8218 17730 8219
rect 18830 7854 18858 7882
rect 20006 7742 20034 7770
rect 18942 7574 18970 7602
rect 17598 7461 17626 7462
rect 17598 7435 17599 7461
rect 17599 7435 17625 7461
rect 17625 7435 17626 7461
rect 17598 7434 17626 7435
rect 17650 7461 17678 7462
rect 17650 7435 17651 7461
rect 17651 7435 17677 7461
rect 17677 7435 17678 7461
rect 17650 7434 17678 7435
rect 17702 7461 17730 7462
rect 17702 7435 17703 7461
rect 17703 7435 17729 7461
rect 17729 7435 17730 7461
rect 17702 7434 17730 7435
rect 20006 7406 20034 7434
rect 12614 7265 12642 7266
rect 12614 7239 12615 7265
rect 12615 7239 12641 7265
rect 12641 7239 12642 7265
rect 12614 7238 12642 7239
rect 12166 6873 12194 6874
rect 12166 6847 12167 6873
rect 12167 6847 12193 6873
rect 12193 6847 12194 6873
rect 12166 6846 12194 6847
rect 12222 6510 12250 6538
rect 12614 6510 12642 6538
rect 9918 3933 9946 3934
rect 9918 3907 9919 3933
rect 9919 3907 9945 3933
rect 9945 3907 9946 3933
rect 9918 3906 9946 3907
rect 9970 3933 9998 3934
rect 9970 3907 9971 3933
rect 9971 3907 9997 3933
rect 9997 3907 9998 3933
rect 9970 3906 9998 3907
rect 10022 3933 10050 3934
rect 10022 3907 10023 3933
rect 10023 3907 10049 3933
rect 10049 3907 10050 3933
rect 10022 3906 10050 3907
rect 9918 3149 9946 3150
rect 9918 3123 9919 3149
rect 9919 3123 9945 3149
rect 9945 3123 9946 3149
rect 9918 3122 9946 3123
rect 9970 3149 9998 3150
rect 9970 3123 9971 3149
rect 9971 3123 9997 3149
rect 9997 3123 9998 3149
rect 9970 3122 9998 3123
rect 10022 3149 10050 3150
rect 10022 3123 10023 3149
rect 10023 3123 10049 3149
rect 10049 3123 10050 3149
rect 10022 3122 10050 3123
rect 9918 2365 9946 2366
rect 9918 2339 9919 2365
rect 9919 2339 9945 2365
rect 9945 2339 9946 2365
rect 9918 2338 9946 2339
rect 9970 2365 9998 2366
rect 9970 2339 9971 2365
rect 9971 2339 9997 2365
rect 9997 2339 9998 2365
rect 9970 2338 9998 2339
rect 10022 2365 10050 2366
rect 10022 2339 10023 2365
rect 10023 2339 10049 2365
rect 10049 2339 10050 2365
rect 10022 2338 10050 2339
rect 10430 1806 10458 1834
rect 9918 1581 9946 1582
rect 9918 1555 9919 1581
rect 9919 1555 9945 1581
rect 9945 1555 9946 1581
rect 9918 1554 9946 1555
rect 9970 1581 9998 1582
rect 9970 1555 9971 1581
rect 9971 1555 9997 1581
rect 9997 1555 9998 1581
rect 9970 1554 9998 1555
rect 10022 1581 10050 1582
rect 10022 1555 10023 1581
rect 10023 1555 10049 1581
rect 10049 1555 10050 1581
rect 10022 1554 10050 1555
rect 11046 1833 11074 1834
rect 11046 1807 11047 1833
rect 11047 1807 11073 1833
rect 11073 1807 11074 1833
rect 11046 1806 11074 1807
rect 11438 1806 11466 1834
rect 17598 6677 17626 6678
rect 17598 6651 17599 6677
rect 17599 6651 17625 6677
rect 17625 6651 17626 6677
rect 17598 6650 17626 6651
rect 17650 6677 17678 6678
rect 17650 6651 17651 6677
rect 17651 6651 17677 6677
rect 17677 6651 17678 6677
rect 17650 6650 17678 6651
rect 17702 6677 17730 6678
rect 17702 6651 17703 6677
rect 17703 6651 17729 6677
rect 17729 6651 17730 6677
rect 17702 6650 17730 6651
rect 17598 5893 17626 5894
rect 17598 5867 17599 5893
rect 17599 5867 17625 5893
rect 17625 5867 17626 5893
rect 17598 5866 17626 5867
rect 17650 5893 17678 5894
rect 17650 5867 17651 5893
rect 17651 5867 17677 5893
rect 17677 5867 17678 5893
rect 17650 5866 17678 5867
rect 17702 5893 17730 5894
rect 17702 5867 17703 5893
rect 17703 5867 17729 5893
rect 17729 5867 17730 5893
rect 17702 5866 17730 5867
rect 17598 5109 17626 5110
rect 17598 5083 17599 5109
rect 17599 5083 17625 5109
rect 17625 5083 17626 5109
rect 17598 5082 17626 5083
rect 17650 5109 17678 5110
rect 17650 5083 17651 5109
rect 17651 5083 17677 5109
rect 17677 5083 17678 5109
rect 17650 5082 17678 5083
rect 17702 5109 17730 5110
rect 17702 5083 17703 5109
rect 17703 5083 17729 5109
rect 17729 5083 17730 5109
rect 17702 5082 17730 5083
rect 17598 4325 17626 4326
rect 17598 4299 17599 4325
rect 17599 4299 17625 4325
rect 17625 4299 17626 4325
rect 17598 4298 17626 4299
rect 17650 4325 17678 4326
rect 17650 4299 17651 4325
rect 17651 4299 17677 4325
rect 17677 4299 17678 4325
rect 17650 4298 17678 4299
rect 17702 4325 17730 4326
rect 17702 4299 17703 4325
rect 17703 4299 17729 4325
rect 17729 4299 17730 4325
rect 17702 4298 17730 4299
rect 17598 3541 17626 3542
rect 17598 3515 17599 3541
rect 17599 3515 17625 3541
rect 17625 3515 17626 3541
rect 17598 3514 17626 3515
rect 17650 3541 17678 3542
rect 17650 3515 17651 3541
rect 17651 3515 17677 3541
rect 17677 3515 17678 3541
rect 17650 3514 17678 3515
rect 17702 3541 17730 3542
rect 17702 3515 17703 3541
rect 17703 3515 17729 3541
rect 17729 3515 17730 3541
rect 17702 3514 17730 3515
rect 17598 2757 17626 2758
rect 17598 2731 17599 2757
rect 17599 2731 17625 2757
rect 17625 2731 17626 2757
rect 17598 2730 17626 2731
rect 17650 2757 17678 2758
rect 17650 2731 17651 2757
rect 17651 2731 17677 2757
rect 17677 2731 17678 2757
rect 17650 2730 17678 2731
rect 17702 2757 17730 2758
rect 17702 2731 17703 2757
rect 17703 2731 17729 2757
rect 17729 2731 17730 2757
rect 17702 2730 17730 2731
rect 12446 2030 12474 2058
rect 13118 2057 13146 2058
rect 13118 2031 13119 2057
rect 13119 2031 13145 2057
rect 13145 2031 13146 2057
rect 13118 2030 13146 2031
rect 17598 1973 17626 1974
rect 17598 1947 17599 1973
rect 17599 1947 17625 1973
rect 17625 1947 17626 1973
rect 17598 1946 17626 1947
rect 17650 1973 17678 1974
rect 17650 1947 17651 1973
rect 17651 1947 17677 1973
rect 17677 1947 17678 1973
rect 17650 1946 17678 1947
rect 17702 1973 17730 1974
rect 17702 1947 17703 1973
rect 17703 1947 17729 1973
rect 17729 1947 17730 1973
rect 17702 1946 17730 1947
rect 12782 1833 12810 1834
rect 12782 1807 12783 1833
rect 12783 1807 12809 1833
rect 12809 1807 12810 1833
rect 12782 1806 12810 1807
<< metal3 >>
rect 12777 19278 12782 19306
rect 12810 19278 13398 19306
rect 13426 19278 13431 19306
rect 2233 19194 2238 19222
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2370 19194 2375 19222
rect 17593 19194 17598 19222
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17730 19194 17735 19222
rect 10425 19110 10430 19138
rect 10458 19110 11046 19138
rect 11074 19110 11079 19138
rect 11433 19110 11438 19138
rect 11466 19110 12782 19138
rect 12810 19110 12815 19138
rect 9913 18802 9918 18830
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 10050 18802 10055 18830
rect 10089 18718 10094 18746
rect 10122 18718 10710 18746
rect 10738 18718 10743 18746
rect 20600 18522 21000 18536
rect 20113 18494 20118 18522
rect 20146 18494 21000 18522
rect 20600 18480 21000 18494
rect 2233 18410 2238 18438
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2370 18410 2375 18438
rect 17593 18410 17598 18438
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17730 18410 17735 18438
rect 9913 18018 9918 18046
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 10050 18018 10055 18046
rect 2233 17626 2238 17654
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2370 17626 2375 17654
rect 17593 17626 17598 17654
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17730 17626 17735 17654
rect 9913 17234 9918 17262
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 10050 17234 10055 17262
rect 20600 17178 21000 17192
rect 20113 17150 20118 17178
rect 20146 17150 21000 17178
rect 20600 17136 21000 17150
rect 2233 16842 2238 16870
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2370 16842 2375 16870
rect 17593 16842 17598 16870
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17730 16842 17735 16870
rect 9913 16450 9918 16478
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 10050 16450 10055 16478
rect 2233 16058 2238 16086
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2370 16058 2375 16086
rect 17593 16058 17598 16086
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17730 16058 17735 16086
rect 9913 15666 9918 15694
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 10050 15666 10055 15694
rect 2233 15274 2238 15302
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2370 15274 2375 15302
rect 17593 15274 17598 15302
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17730 15274 17735 15302
rect 9913 14882 9918 14910
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 10050 14882 10055 14910
rect 2233 14490 2238 14518
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2370 14490 2375 14518
rect 17593 14490 17598 14518
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17730 14490 17735 14518
rect 11713 14126 11718 14154
rect 11746 14126 12278 14154
rect 12306 14126 12311 14154
rect 9913 14098 9918 14126
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 10050 14098 10055 14126
rect 2233 13706 2238 13734
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2370 13706 2375 13734
rect 17593 13706 17598 13734
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17730 13706 17735 13734
rect 11153 13566 11158 13594
rect 11186 13566 13062 13594
rect 13090 13566 13342 13594
rect 13370 13566 13375 13594
rect 2137 13510 2142 13538
rect 2170 13510 6622 13538
rect 6650 13510 6655 13538
rect 11097 13510 11102 13538
rect 11130 13510 11662 13538
rect 11690 13510 11695 13538
rect 11993 13510 11998 13538
rect 12026 13510 12894 13538
rect 12922 13510 12927 13538
rect 0 13482 400 13496
rect 20600 13482 21000 13496
rect 0 13454 2086 13482
rect 2114 13454 2119 13482
rect 10089 13454 10094 13482
rect 10122 13454 11158 13482
rect 11186 13454 11191 13482
rect 11377 13454 11382 13482
rect 11410 13454 12222 13482
rect 12250 13454 12255 13482
rect 13393 13454 13398 13482
rect 13426 13454 14630 13482
rect 14658 13454 14663 13482
rect 19945 13454 19950 13482
rect 19978 13454 21000 13482
rect 0 13440 400 13454
rect 11382 13426 11410 13454
rect 20600 13440 21000 13454
rect 9305 13398 9310 13426
rect 9338 13398 10150 13426
rect 10178 13398 10183 13426
rect 10313 13398 10318 13426
rect 10346 13398 11410 13426
rect 9913 13314 9918 13342
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 10050 13314 10055 13342
rect 9697 13230 9702 13258
rect 9730 13230 10374 13258
rect 10402 13230 10766 13258
rect 10794 13230 10799 13258
rect 15946 13230 18830 13258
rect 18858 13230 18863 13258
rect 15946 13202 15974 13230
rect 9193 13174 9198 13202
rect 9226 13174 9478 13202
rect 9506 13174 9511 13202
rect 14961 13174 14966 13202
rect 14994 13174 15974 13202
rect 0 13146 400 13160
rect 20600 13146 21000 13160
rect 0 13118 966 13146
rect 994 13118 999 13146
rect 2137 13118 2142 13146
rect 2170 13118 5950 13146
rect 5978 13118 5983 13146
rect 15946 13118 18830 13146
rect 18858 13118 18863 13146
rect 20001 13118 20006 13146
rect 20034 13118 21000 13146
rect 0 13104 400 13118
rect 15946 13090 15974 13118
rect 20600 13104 21000 13118
rect 6617 13062 6622 13090
rect 6650 13062 7630 13090
rect 7658 13062 7663 13090
rect 8017 13062 8022 13090
rect 8050 13062 8302 13090
rect 8330 13062 8974 13090
rect 9002 13062 9007 13090
rect 14793 13062 14798 13090
rect 14826 13062 15974 13090
rect 2233 12922 2238 12950
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2370 12922 2375 12950
rect 17593 12922 17598 12950
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17730 12922 17735 12950
rect 12945 12838 12950 12866
rect 12978 12838 13510 12866
rect 13538 12838 18942 12866
rect 18970 12838 18975 12866
rect 0 12810 400 12824
rect 20600 12810 21000 12824
rect 0 12782 966 12810
rect 994 12782 999 12810
rect 8969 12782 8974 12810
rect 9002 12782 10374 12810
rect 10402 12782 10407 12810
rect 20001 12782 20006 12810
rect 20034 12782 21000 12810
rect 0 12768 400 12782
rect 20600 12768 21000 12782
rect 7546 12726 7686 12754
rect 7714 12726 7719 12754
rect 10145 12726 10150 12754
rect 10178 12726 10318 12754
rect 10346 12726 11942 12754
rect 11970 12726 11975 12754
rect 7546 12698 7574 12726
rect 7345 12670 7350 12698
rect 7378 12670 7574 12698
rect 9361 12614 9366 12642
rect 9394 12614 10038 12642
rect 10066 12614 10990 12642
rect 11018 12614 11023 12642
rect 12105 12614 12110 12642
rect 12138 12614 12726 12642
rect 12754 12614 13174 12642
rect 13202 12614 13398 12642
rect 13426 12614 14014 12642
rect 14042 12614 14047 12642
rect 9913 12530 9918 12558
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 10050 12530 10055 12558
rect 6841 12502 6846 12530
rect 6874 12502 7742 12530
rect 7770 12502 7775 12530
rect 7625 12446 7630 12474
rect 7658 12446 9142 12474
rect 9170 12446 9422 12474
rect 9450 12446 9455 12474
rect 7401 12390 7406 12418
rect 7434 12390 7574 12418
rect 7602 12390 8022 12418
rect 8050 12390 8055 12418
rect 5945 12334 5950 12362
rect 5978 12334 7686 12362
rect 7714 12334 7719 12362
rect 9081 12334 9086 12362
rect 9114 12334 9814 12362
rect 9842 12334 12390 12362
rect 12418 12334 12423 12362
rect 2233 12138 2238 12166
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2370 12138 2375 12166
rect 17593 12138 17598 12166
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17730 12138 17735 12166
rect 2137 11942 2142 11970
rect 2170 11942 5670 11970
rect 5698 11942 7406 11970
rect 7434 11942 7439 11970
rect 0 11802 400 11816
rect 0 11774 966 11802
rect 994 11774 999 11802
rect 13225 11774 13230 11802
rect 13258 11774 13734 11802
rect 13762 11774 13767 11802
rect 0 11760 400 11774
rect 9913 11746 9918 11774
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 10050 11746 10055 11774
rect 7905 11662 7910 11690
rect 7938 11662 8078 11690
rect 8106 11662 10206 11690
rect 10234 11662 10239 11690
rect 13001 11662 13006 11690
rect 13034 11662 13398 11690
rect 13426 11662 14630 11690
rect 14658 11662 14663 11690
rect 7961 11606 7966 11634
rect 7994 11606 8862 11634
rect 8890 11606 9590 11634
rect 9618 11606 9623 11634
rect 12721 11606 12726 11634
rect 12754 11606 13454 11634
rect 8689 11550 8694 11578
rect 8722 11550 9030 11578
rect 9058 11550 9063 11578
rect 12105 11550 12110 11578
rect 12138 11550 12614 11578
rect 12642 11550 12782 11578
rect 12810 11550 12815 11578
rect 13426 11522 13454 11606
rect 15946 11550 18830 11578
rect 18858 11550 18863 11578
rect 15946 11522 15974 11550
rect 6785 11494 6790 11522
rect 6818 11494 7574 11522
rect 7602 11494 7607 11522
rect 13426 11494 14406 11522
rect 14434 11494 15974 11522
rect 20600 11466 21000 11480
rect 20001 11438 20006 11466
rect 20034 11438 21000 11466
rect 20600 11424 21000 11438
rect 2233 11354 2238 11382
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2370 11354 2375 11382
rect 17593 11354 17598 11382
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17730 11354 17735 11382
rect 9641 11326 9646 11354
rect 9674 11326 10038 11354
rect 10066 11326 10071 11354
rect 961 11214 966 11242
rect 994 11214 999 11242
rect 11489 11214 11494 11242
rect 11522 11214 12838 11242
rect 12866 11214 13342 11242
rect 13370 11214 13375 11242
rect 0 11130 400 11144
rect 966 11130 994 11214
rect 7289 11158 7294 11186
rect 7322 11158 8862 11186
rect 8890 11158 8895 11186
rect 12049 11158 12054 11186
rect 12082 11158 12894 11186
rect 12922 11158 12927 11186
rect 13426 11158 13790 11186
rect 13818 11158 13823 11186
rect 13426 11130 13454 11158
rect 20600 11130 21000 11144
rect 0 11102 994 11130
rect 7793 11102 7798 11130
rect 7826 11102 8638 11130
rect 8666 11102 9254 11130
rect 9282 11102 9287 11130
rect 12161 11102 12166 11130
rect 12194 11102 13454 11130
rect 20001 11102 20006 11130
rect 20034 11102 21000 11130
rect 0 11088 400 11102
rect 20600 11088 21000 11102
rect 6729 11046 6734 11074
rect 6762 11046 7350 11074
rect 7378 11046 7383 11074
rect 7737 11046 7742 11074
rect 7770 11046 7966 11074
rect 7994 11046 7999 11074
rect 9814 11046 9870 11074
rect 9898 11046 9903 11074
rect 10313 11046 10318 11074
rect 10346 11046 11494 11074
rect 11522 11046 11527 11074
rect 12777 11046 12782 11074
rect 12810 11046 13062 11074
rect 13090 11046 13095 11074
rect 9814 10906 9842 11046
rect 12665 10990 12670 11018
rect 12698 10990 13622 11018
rect 13650 10990 13655 11018
rect 9913 10962 9918 10990
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 10050 10962 10055 10990
rect 10817 10934 10822 10962
rect 10850 10934 12334 10962
rect 12362 10934 12367 10962
rect 12777 10934 12782 10962
rect 12810 10934 13286 10962
rect 13314 10934 13319 10962
rect 8297 10878 8302 10906
rect 8330 10878 9534 10906
rect 9562 10878 9567 10906
rect 9697 10878 9702 10906
rect 9730 10878 9842 10906
rect 10257 10878 10262 10906
rect 10290 10878 11886 10906
rect 11914 10878 11919 10906
rect 11993 10878 11998 10906
rect 12026 10878 12950 10906
rect 12978 10878 12983 10906
rect 2137 10822 2142 10850
rect 2170 10822 5726 10850
rect 5754 10822 7462 10850
rect 7490 10822 7495 10850
rect 9361 10822 9366 10850
rect 9394 10822 10038 10850
rect 10066 10822 11774 10850
rect 11802 10822 11807 10850
rect 11998 10794 12026 10878
rect 12889 10822 12894 10850
rect 12922 10822 13454 10850
rect 13426 10794 13454 10822
rect 7737 10766 7742 10794
rect 7770 10766 9870 10794
rect 9898 10766 10710 10794
rect 10738 10766 10743 10794
rect 11041 10766 11046 10794
rect 11074 10766 11438 10794
rect 11466 10766 12026 10794
rect 12329 10766 12334 10794
rect 12362 10766 12950 10794
rect 12978 10766 13342 10794
rect 13370 10766 13375 10794
rect 13426 10766 14742 10794
rect 14770 10766 18830 10794
rect 18858 10766 18863 10794
rect 2081 10710 2086 10738
rect 2114 10710 9310 10738
rect 9338 10710 9343 10738
rect 10313 10710 10318 10738
rect 10346 10710 10822 10738
rect 10850 10710 10855 10738
rect 11377 10710 11382 10738
rect 11410 10710 12614 10738
rect 12642 10710 12647 10738
rect 7401 10654 7406 10682
rect 7434 10654 7742 10682
rect 7770 10654 7775 10682
rect 8017 10654 8022 10682
rect 8050 10654 11270 10682
rect 11298 10654 11942 10682
rect 11970 10654 11975 10682
rect 7681 10598 7686 10626
rect 7714 10598 11326 10626
rect 11354 10598 11359 10626
rect 12385 10598 12390 10626
rect 12418 10598 12726 10626
rect 12754 10598 12759 10626
rect 2233 10570 2238 10598
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2370 10570 2375 10598
rect 17593 10570 17598 10598
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17730 10570 17735 10598
rect 7849 10542 7854 10570
rect 7882 10542 8358 10570
rect 8386 10542 10430 10570
rect 10458 10542 10934 10570
rect 10962 10542 10967 10570
rect 10201 10486 10206 10514
rect 10234 10486 10542 10514
rect 10570 10486 10575 10514
rect 10817 10486 10822 10514
rect 10850 10486 12726 10514
rect 12754 10486 13230 10514
rect 13258 10486 13263 10514
rect 6561 10430 6566 10458
rect 6594 10430 7294 10458
rect 7322 10430 7630 10458
rect 7658 10430 7663 10458
rect 10481 10430 10486 10458
rect 10514 10430 10878 10458
rect 10906 10430 11886 10458
rect 11914 10430 12222 10458
rect 12250 10430 12255 10458
rect 10033 10374 10038 10402
rect 10066 10374 11158 10402
rect 11186 10374 11191 10402
rect 8969 10262 8974 10290
rect 9002 10262 9926 10290
rect 9954 10262 9959 10290
rect 9913 10178 9918 10206
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 10050 10178 10055 10206
rect 12329 10150 12334 10178
rect 12362 10150 12782 10178
rect 12810 10150 12815 10178
rect 7569 10094 7574 10122
rect 7602 10094 8078 10122
rect 8106 10094 8806 10122
rect 8834 10094 8839 10122
rect 9193 10094 9198 10122
rect 9226 10094 9702 10122
rect 9730 10094 12390 10122
rect 12418 10094 12423 10122
rect 12609 10094 12614 10122
rect 12642 10094 13006 10122
rect 13034 10094 13039 10122
rect 13505 10094 13510 10122
rect 13538 10094 13543 10122
rect 7065 10038 7070 10066
rect 7098 10038 7406 10066
rect 7434 10038 7742 10066
rect 7770 10038 7775 10066
rect 8017 10038 8022 10066
rect 8050 10038 8666 10066
rect 8745 10038 8750 10066
rect 8778 10038 9198 10066
rect 9226 10038 10206 10066
rect 10234 10038 10239 10066
rect 8638 10010 8666 10038
rect 13510 10010 13538 10094
rect 4993 9982 4998 10010
rect 5026 9982 7238 10010
rect 7266 9982 7271 10010
rect 7961 9982 7966 10010
rect 7994 9982 8246 10010
rect 8274 9982 8279 10010
rect 8633 9982 8638 10010
rect 8666 9982 9030 10010
rect 9058 9982 9702 10010
rect 9730 9982 10654 10010
rect 10682 9982 10687 10010
rect 12497 9982 12502 10010
rect 12530 9982 13118 10010
rect 13146 9982 13151 10010
rect 13281 9982 13286 10010
rect 13314 9982 13538 10010
rect 10985 9926 10990 9954
rect 11018 9926 12278 9954
rect 12306 9926 12311 9954
rect 13337 9926 13342 9954
rect 13370 9926 13958 9954
rect 13986 9926 13991 9954
rect 14681 9926 14686 9954
rect 14714 9926 15022 9954
rect 15050 9926 18830 9954
rect 18858 9926 18863 9954
rect 7737 9870 7742 9898
rect 7770 9870 9142 9898
rect 9170 9870 9175 9898
rect 13057 9870 13062 9898
rect 13090 9870 13398 9898
rect 13426 9870 13431 9898
rect 8465 9814 8470 9842
rect 8498 9814 8862 9842
rect 8890 9814 11326 9842
rect 11354 9814 11359 9842
rect 2233 9786 2238 9814
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2370 9786 2375 9814
rect 17593 9786 17598 9814
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17730 9786 17735 9814
rect 7289 9758 7294 9786
rect 7322 9758 7574 9786
rect 10649 9758 10654 9786
rect 10682 9758 12614 9786
rect 12642 9758 12647 9786
rect 7546 9702 7574 9758
rect 7602 9702 7607 9730
rect 9249 9702 9254 9730
rect 9282 9702 12222 9730
rect 12250 9702 12255 9730
rect 4186 9646 4998 9674
rect 5026 9646 5031 9674
rect 7737 9646 7742 9674
rect 7770 9646 7910 9674
rect 7938 9646 7943 9674
rect 4186 9618 4214 9646
rect 2137 9590 2142 9618
rect 2170 9590 4214 9618
rect 6953 9590 6958 9618
rect 6986 9590 7686 9618
rect 7714 9590 8358 9618
rect 8386 9590 9422 9618
rect 9450 9590 9702 9618
rect 9730 9590 9735 9618
rect 9865 9590 9870 9618
rect 9898 9590 10318 9618
rect 10346 9590 10822 9618
rect 10850 9590 10855 9618
rect 14065 9590 14070 9618
rect 14098 9590 14630 9618
rect 14658 9590 14663 9618
rect 7625 9534 7630 9562
rect 7658 9534 8246 9562
rect 8274 9534 8750 9562
rect 8778 9534 9030 9562
rect 9058 9534 9063 9562
rect 6057 9478 6062 9506
rect 6090 9478 6902 9506
rect 6930 9478 6935 9506
rect 8633 9478 8638 9506
rect 8666 9478 10486 9506
rect 10514 9478 13622 9506
rect 13650 9478 13655 9506
rect 0 9450 400 9464
rect 20600 9450 21000 9464
rect 0 9422 966 9450
rect 994 9422 999 9450
rect 20001 9422 20006 9450
rect 20034 9422 21000 9450
rect 0 9408 400 9422
rect 9913 9394 9918 9422
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 10050 9394 10055 9422
rect 20600 9408 21000 9422
rect 7625 9366 7630 9394
rect 7658 9366 7910 9394
rect 7938 9366 9254 9394
rect 9282 9366 9287 9394
rect 10369 9366 10374 9394
rect 10402 9366 11046 9394
rect 11074 9366 11438 9394
rect 11466 9366 12502 9394
rect 12530 9366 12535 9394
rect 8801 9310 8806 9338
rect 8834 9310 9982 9338
rect 10010 9310 10262 9338
rect 10290 9310 10295 9338
rect 11545 9310 11550 9338
rect 11578 9310 11774 9338
rect 11802 9310 12110 9338
rect 12138 9310 12143 9338
rect 7625 9254 7630 9282
rect 7658 9254 8470 9282
rect 8498 9254 8503 9282
rect 9249 9254 9254 9282
rect 9282 9254 10374 9282
rect 10402 9254 10407 9282
rect 5049 9198 5054 9226
rect 5082 9198 6398 9226
rect 6426 9198 6431 9226
rect 8059 9198 8078 9226
rect 8106 9198 8111 9226
rect 8185 9198 8190 9226
rect 8218 9198 8806 9226
rect 8834 9198 8839 9226
rect 8969 9198 8974 9226
rect 9002 9198 9086 9226
rect 9114 9198 9590 9226
rect 9618 9198 11606 9226
rect 11634 9198 11639 9226
rect 15946 9198 18830 9226
rect 18858 9198 18863 9226
rect 15946 9170 15974 9198
rect 5385 9142 5390 9170
rect 5418 9142 9310 9170
rect 9338 9142 9343 9170
rect 9417 9142 9422 9170
rect 9450 9142 10094 9170
rect 10122 9142 10654 9170
rect 10682 9142 10687 9170
rect 13169 9142 13174 9170
rect 13202 9142 13790 9170
rect 13818 9142 13823 9170
rect 13953 9142 13958 9170
rect 13986 9142 14574 9170
rect 14602 9142 15974 9170
rect 20600 9114 21000 9128
rect 7121 9086 7126 9114
rect 7154 9086 7574 9114
rect 7961 9086 7966 9114
rect 7994 9086 8694 9114
rect 8722 9086 8727 9114
rect 9179 9086 9198 9114
rect 9226 9086 9231 9114
rect 11601 9086 11606 9114
rect 11634 9086 12278 9114
rect 12306 9086 12311 9114
rect 20001 9086 20006 9114
rect 20034 9086 21000 9114
rect 7546 9058 7574 9086
rect 20600 9072 21000 9086
rect 7546 9030 8638 9058
rect 8666 9030 8671 9058
rect 11097 9030 11102 9058
rect 11130 9030 13062 9058
rect 13090 9030 13095 9058
rect 2233 9002 2238 9030
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2370 9002 2375 9030
rect 17593 9002 17598 9030
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17730 9002 17735 9030
rect 8073 8974 8078 9002
rect 8106 8974 10654 9002
rect 10682 8974 10687 9002
rect 7457 8918 7462 8946
rect 7490 8918 9870 8946
rect 9898 8918 9903 8946
rect 7546 8862 7686 8890
rect 7714 8862 8302 8890
rect 8330 8862 8335 8890
rect 7546 8778 7574 8862
rect 7737 8806 7742 8834
rect 7770 8806 8526 8834
rect 8554 8806 8559 8834
rect 9249 8806 9254 8834
rect 9282 8806 9982 8834
rect 10010 8806 10015 8834
rect 12161 8806 12166 8834
rect 12194 8806 13174 8834
rect 13202 8806 13207 8834
rect 13281 8806 13286 8834
rect 13314 8806 13846 8834
rect 13874 8806 13879 8834
rect 7121 8750 7126 8778
rect 7154 8750 7574 8778
rect 6449 8694 6454 8722
rect 6482 8694 6790 8722
rect 6818 8694 6823 8722
rect 7177 8694 7182 8722
rect 7210 8694 7910 8722
rect 7938 8694 7943 8722
rect 9913 8610 9918 8638
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 10050 8610 10055 8638
rect 7546 8526 10178 8554
rect 7546 8498 7574 8526
rect 10150 8498 10178 8526
rect 6953 8470 6958 8498
rect 6986 8470 7574 8498
rect 7905 8470 7910 8498
rect 7938 8470 8190 8498
rect 8218 8470 8223 8498
rect 10145 8470 10150 8498
rect 10178 8470 11550 8498
rect 11578 8470 11583 8498
rect 7401 8414 7406 8442
rect 7434 8414 7630 8442
rect 7658 8414 7854 8442
rect 7882 8414 7887 8442
rect 8073 8414 8078 8442
rect 8106 8414 8862 8442
rect 8890 8414 8895 8442
rect 9473 8414 9478 8442
rect 9506 8414 9646 8442
rect 9674 8414 10206 8442
rect 10234 8414 10239 8442
rect 8185 8358 8190 8386
rect 8218 8358 8414 8386
rect 8442 8358 8918 8386
rect 8946 8358 9534 8386
rect 9562 8358 9567 8386
rect 9697 8358 9702 8386
rect 9730 8358 10038 8386
rect 10066 8358 10071 8386
rect 12665 8358 12670 8386
rect 12698 8358 12950 8386
rect 12978 8358 14462 8386
rect 14490 8358 14495 8386
rect 10761 8302 10766 8330
rect 10794 8302 13230 8330
rect 13258 8302 13263 8330
rect 9473 8246 9478 8274
rect 9506 8246 12614 8274
rect 12642 8246 13006 8274
rect 13034 8246 13286 8274
rect 13314 8246 13319 8274
rect 2233 8218 2238 8246
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2370 8218 2375 8246
rect 17593 8218 17598 8246
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17730 8218 17735 8246
rect 7625 8078 7630 8106
rect 7658 8078 8246 8106
rect 8274 8078 8279 8106
rect 12329 8022 12334 8050
rect 12362 8022 12726 8050
rect 12754 8022 13342 8050
rect 13370 8022 13375 8050
rect 11321 7966 11326 7994
rect 11354 7966 11662 7994
rect 11690 7966 11695 7994
rect 13281 7966 13286 7994
rect 13314 7966 13566 7994
rect 13594 7966 13790 7994
rect 13818 7966 13823 7994
rect 10369 7910 10374 7938
rect 10402 7910 11270 7938
rect 11298 7910 11303 7938
rect 11433 7910 11438 7938
rect 11466 7910 11830 7938
rect 11858 7910 11863 7938
rect 12105 7910 12110 7938
rect 12138 7910 13398 7938
rect 13426 7910 13431 7938
rect 11377 7854 11382 7882
rect 11410 7854 11998 7882
rect 12026 7854 12031 7882
rect 13505 7854 13510 7882
rect 13538 7854 14070 7882
rect 14098 7854 18830 7882
rect 18858 7854 18863 7882
rect 9913 7826 9918 7854
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 10050 7826 10055 7854
rect 11550 7798 12222 7826
rect 12250 7798 12782 7826
rect 12810 7798 12815 7826
rect 11550 7770 11578 7798
rect 20600 7770 21000 7784
rect 9809 7742 9814 7770
rect 9842 7742 11578 7770
rect 11825 7742 11830 7770
rect 11858 7742 12334 7770
rect 12362 7742 12367 7770
rect 20001 7742 20006 7770
rect 20034 7742 21000 7770
rect 20600 7728 21000 7742
rect 5945 7686 5950 7714
rect 5978 7686 7686 7714
rect 7714 7686 7719 7714
rect 9753 7686 9758 7714
rect 9786 7686 11998 7714
rect 12026 7686 12031 7714
rect 10873 7630 10878 7658
rect 10906 7630 11438 7658
rect 11466 7630 11471 7658
rect 5609 7574 5614 7602
rect 5642 7574 6790 7602
rect 6818 7574 6823 7602
rect 10705 7574 10710 7602
rect 10738 7574 12670 7602
rect 12698 7574 12703 7602
rect 13225 7574 13230 7602
rect 13258 7574 14238 7602
rect 14266 7574 18942 7602
rect 18970 7574 18975 7602
rect 9249 7518 9254 7546
rect 9282 7518 9534 7546
rect 9562 7518 10038 7546
rect 10066 7518 10071 7546
rect 2233 7434 2238 7462
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2370 7434 2375 7462
rect 17593 7434 17598 7462
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17730 7434 17735 7462
rect 20600 7434 21000 7448
rect 20001 7406 20006 7434
rect 20034 7406 21000 7434
rect 20600 7392 21000 7406
rect 9641 7294 9646 7322
rect 9674 7294 10486 7322
rect 10514 7294 10519 7322
rect 12161 7294 12166 7322
rect 12194 7294 13006 7322
rect 13034 7294 13039 7322
rect 8633 7238 8638 7266
rect 8666 7238 9422 7266
rect 9450 7238 10094 7266
rect 10369 7238 10374 7266
rect 10402 7238 10407 7266
rect 10705 7238 10710 7266
rect 10738 7238 11214 7266
rect 11242 7238 12334 7266
rect 12362 7238 12614 7266
rect 12642 7238 12647 7266
rect 10066 7210 10094 7238
rect 10374 7210 10402 7238
rect 9921 7182 9926 7210
rect 9954 7182 9959 7210
rect 10066 7182 10402 7210
rect 9926 7154 9954 7182
rect 7401 7126 7406 7154
rect 7434 7126 7742 7154
rect 7770 7126 8414 7154
rect 8442 7126 8974 7154
rect 9002 7126 9007 7154
rect 9926 7126 10150 7154
rect 10178 7126 10183 7154
rect 9913 7042 9918 7070
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 10050 7042 10055 7070
rect 8409 6846 8414 6874
rect 8442 6846 8750 6874
rect 8778 6846 8783 6874
rect 8913 6846 8918 6874
rect 8946 6846 9310 6874
rect 9338 6846 9343 6874
rect 11545 6846 11550 6874
rect 11578 6846 12166 6874
rect 12194 6846 12199 6874
rect 8969 6790 8974 6818
rect 9002 6790 9254 6818
rect 9282 6790 9646 6818
rect 9674 6790 9679 6818
rect 2233 6650 2238 6678
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2370 6650 2375 6678
rect 17593 6650 17598 6678
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17730 6650 17735 6678
rect 8801 6510 8806 6538
rect 8834 6510 9142 6538
rect 9170 6510 9366 6538
rect 9394 6510 9399 6538
rect 12217 6510 12222 6538
rect 12250 6510 12614 6538
rect 12642 6510 12647 6538
rect 9913 6258 9918 6286
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 10050 6258 10055 6286
rect 2233 5866 2238 5894
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2370 5866 2375 5894
rect 17593 5866 17598 5894
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17730 5866 17735 5894
rect 9913 5474 9918 5502
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 10050 5474 10055 5502
rect 2233 5082 2238 5110
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2370 5082 2375 5110
rect 17593 5082 17598 5110
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17730 5082 17735 5110
rect 9913 4690 9918 4718
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 10050 4690 10055 4718
rect 2233 4298 2238 4326
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2370 4298 2375 4326
rect 17593 4298 17598 4326
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17730 4298 17735 4326
rect 9913 3906 9918 3934
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 10050 3906 10055 3934
rect 2233 3514 2238 3542
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2370 3514 2375 3542
rect 17593 3514 17598 3542
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17730 3514 17735 3542
rect 9913 3122 9918 3150
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 10050 3122 10055 3150
rect 2233 2730 2238 2758
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2370 2730 2375 2758
rect 17593 2730 17598 2758
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17730 2730 17735 2758
rect 9913 2338 9918 2366
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 10050 2338 10055 2366
rect 12441 2030 12446 2058
rect 12474 2030 13118 2058
rect 13146 2030 13151 2058
rect 2233 1946 2238 1974
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2370 1946 2375 1974
rect 17593 1946 17598 1974
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17730 1946 17735 1974
rect 10425 1806 10430 1834
rect 10458 1806 11046 1834
rect 11074 1806 11079 1834
rect 11433 1806 11438 1834
rect 11466 1806 12782 1834
rect 12810 1806 12815 1834
rect 9913 1554 9918 1582
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 10050 1554 10055 1582
<< via3 >>
rect 2238 19194 2266 19222
rect 2290 19194 2318 19222
rect 2342 19194 2370 19222
rect 17598 19194 17626 19222
rect 17650 19194 17678 19222
rect 17702 19194 17730 19222
rect 9918 18802 9946 18830
rect 9970 18802 9998 18830
rect 10022 18802 10050 18830
rect 2238 18410 2266 18438
rect 2290 18410 2318 18438
rect 2342 18410 2370 18438
rect 17598 18410 17626 18438
rect 17650 18410 17678 18438
rect 17702 18410 17730 18438
rect 9918 18018 9946 18046
rect 9970 18018 9998 18046
rect 10022 18018 10050 18046
rect 2238 17626 2266 17654
rect 2290 17626 2318 17654
rect 2342 17626 2370 17654
rect 17598 17626 17626 17654
rect 17650 17626 17678 17654
rect 17702 17626 17730 17654
rect 9918 17234 9946 17262
rect 9970 17234 9998 17262
rect 10022 17234 10050 17262
rect 2238 16842 2266 16870
rect 2290 16842 2318 16870
rect 2342 16842 2370 16870
rect 17598 16842 17626 16870
rect 17650 16842 17678 16870
rect 17702 16842 17730 16870
rect 9918 16450 9946 16478
rect 9970 16450 9998 16478
rect 10022 16450 10050 16478
rect 2238 16058 2266 16086
rect 2290 16058 2318 16086
rect 2342 16058 2370 16086
rect 17598 16058 17626 16086
rect 17650 16058 17678 16086
rect 17702 16058 17730 16086
rect 9918 15666 9946 15694
rect 9970 15666 9998 15694
rect 10022 15666 10050 15694
rect 2238 15274 2266 15302
rect 2290 15274 2318 15302
rect 2342 15274 2370 15302
rect 17598 15274 17626 15302
rect 17650 15274 17678 15302
rect 17702 15274 17730 15302
rect 9918 14882 9946 14910
rect 9970 14882 9998 14910
rect 10022 14882 10050 14910
rect 2238 14490 2266 14518
rect 2290 14490 2318 14518
rect 2342 14490 2370 14518
rect 17598 14490 17626 14518
rect 17650 14490 17678 14518
rect 17702 14490 17730 14518
rect 9918 14098 9946 14126
rect 9970 14098 9998 14126
rect 10022 14098 10050 14126
rect 2238 13706 2266 13734
rect 2290 13706 2318 13734
rect 2342 13706 2370 13734
rect 17598 13706 17626 13734
rect 17650 13706 17678 13734
rect 17702 13706 17730 13734
rect 9918 13314 9946 13342
rect 9970 13314 9998 13342
rect 10022 13314 10050 13342
rect 2238 12922 2266 12950
rect 2290 12922 2318 12950
rect 2342 12922 2370 12950
rect 17598 12922 17626 12950
rect 17650 12922 17678 12950
rect 17702 12922 17730 12950
rect 9918 12530 9946 12558
rect 9970 12530 9998 12558
rect 10022 12530 10050 12558
rect 2238 12138 2266 12166
rect 2290 12138 2318 12166
rect 2342 12138 2370 12166
rect 17598 12138 17626 12166
rect 17650 12138 17678 12166
rect 17702 12138 17730 12166
rect 9918 11746 9946 11774
rect 9970 11746 9998 11774
rect 10022 11746 10050 11774
rect 8078 11662 8106 11690
rect 2238 11354 2266 11382
rect 2290 11354 2318 11382
rect 2342 11354 2370 11382
rect 17598 11354 17626 11382
rect 17650 11354 17678 11382
rect 17702 11354 17730 11382
rect 9918 10962 9946 10990
rect 9970 10962 9998 10990
rect 10022 10962 10050 10990
rect 2238 10570 2266 10598
rect 2290 10570 2318 10598
rect 2342 10570 2370 10598
rect 17598 10570 17626 10598
rect 17650 10570 17678 10598
rect 17702 10570 17730 10598
rect 9918 10178 9946 10206
rect 9970 10178 9998 10206
rect 10022 10178 10050 10206
rect 9198 10094 9226 10122
rect 2238 9786 2266 9814
rect 2290 9786 2318 9814
rect 2342 9786 2370 9814
rect 17598 9786 17626 9814
rect 17650 9786 17678 9814
rect 17702 9786 17730 9814
rect 9918 9394 9946 9422
rect 9970 9394 9998 9422
rect 10022 9394 10050 9422
rect 8078 9198 8106 9226
rect 9198 9086 9226 9114
rect 2238 9002 2266 9030
rect 2290 9002 2318 9030
rect 2342 9002 2370 9030
rect 17598 9002 17626 9030
rect 17650 9002 17678 9030
rect 17702 9002 17730 9030
rect 9918 8610 9946 8638
rect 9970 8610 9998 8638
rect 10022 8610 10050 8638
rect 2238 8218 2266 8246
rect 2290 8218 2318 8246
rect 2342 8218 2370 8246
rect 17598 8218 17626 8246
rect 17650 8218 17678 8246
rect 17702 8218 17730 8246
rect 9918 7826 9946 7854
rect 9970 7826 9998 7854
rect 10022 7826 10050 7854
rect 2238 7434 2266 7462
rect 2290 7434 2318 7462
rect 2342 7434 2370 7462
rect 17598 7434 17626 7462
rect 17650 7434 17678 7462
rect 17702 7434 17730 7462
rect 9918 7042 9946 7070
rect 9970 7042 9998 7070
rect 10022 7042 10050 7070
rect 2238 6650 2266 6678
rect 2290 6650 2318 6678
rect 2342 6650 2370 6678
rect 17598 6650 17626 6678
rect 17650 6650 17678 6678
rect 17702 6650 17730 6678
rect 9918 6258 9946 6286
rect 9970 6258 9998 6286
rect 10022 6258 10050 6286
rect 2238 5866 2266 5894
rect 2290 5866 2318 5894
rect 2342 5866 2370 5894
rect 17598 5866 17626 5894
rect 17650 5866 17678 5894
rect 17702 5866 17730 5894
rect 9918 5474 9946 5502
rect 9970 5474 9998 5502
rect 10022 5474 10050 5502
rect 2238 5082 2266 5110
rect 2290 5082 2318 5110
rect 2342 5082 2370 5110
rect 17598 5082 17626 5110
rect 17650 5082 17678 5110
rect 17702 5082 17730 5110
rect 9918 4690 9946 4718
rect 9970 4690 9998 4718
rect 10022 4690 10050 4718
rect 2238 4298 2266 4326
rect 2290 4298 2318 4326
rect 2342 4298 2370 4326
rect 17598 4298 17626 4326
rect 17650 4298 17678 4326
rect 17702 4298 17730 4326
rect 9918 3906 9946 3934
rect 9970 3906 9998 3934
rect 10022 3906 10050 3934
rect 2238 3514 2266 3542
rect 2290 3514 2318 3542
rect 2342 3514 2370 3542
rect 17598 3514 17626 3542
rect 17650 3514 17678 3542
rect 17702 3514 17730 3542
rect 9918 3122 9946 3150
rect 9970 3122 9998 3150
rect 10022 3122 10050 3150
rect 2238 2730 2266 2758
rect 2290 2730 2318 2758
rect 2342 2730 2370 2758
rect 17598 2730 17626 2758
rect 17650 2730 17678 2758
rect 17702 2730 17730 2758
rect 9918 2338 9946 2366
rect 9970 2338 9998 2366
rect 10022 2338 10050 2366
rect 2238 1946 2266 1974
rect 2290 1946 2318 1974
rect 2342 1946 2370 1974
rect 17598 1946 17626 1974
rect 17650 1946 17678 1974
rect 17702 1946 17730 1974
rect 9918 1554 9946 1582
rect 9970 1554 9998 1582
rect 10022 1554 10050 1582
<< metal4 >>
rect 2224 19222 2384 19238
rect 2224 19194 2238 19222
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2370 19194 2384 19222
rect 2224 18438 2384 19194
rect 2224 18410 2238 18438
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2370 18410 2384 18438
rect 2224 17654 2384 18410
rect 2224 17626 2238 17654
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2370 17626 2384 17654
rect 2224 16870 2384 17626
rect 2224 16842 2238 16870
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2370 16842 2384 16870
rect 2224 16086 2384 16842
rect 2224 16058 2238 16086
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2370 16058 2384 16086
rect 2224 15302 2384 16058
rect 2224 15274 2238 15302
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2370 15274 2384 15302
rect 2224 14518 2384 15274
rect 2224 14490 2238 14518
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2370 14490 2384 14518
rect 2224 13734 2384 14490
rect 2224 13706 2238 13734
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2370 13706 2384 13734
rect 2224 12950 2384 13706
rect 2224 12922 2238 12950
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2370 12922 2384 12950
rect 2224 12166 2384 12922
rect 2224 12138 2238 12166
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2370 12138 2384 12166
rect 2224 11382 2384 12138
rect 9904 18830 10064 19238
rect 9904 18802 9918 18830
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 10050 18802 10064 18830
rect 9904 18046 10064 18802
rect 9904 18018 9918 18046
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 10050 18018 10064 18046
rect 9904 17262 10064 18018
rect 9904 17234 9918 17262
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 10050 17234 10064 17262
rect 9904 16478 10064 17234
rect 9904 16450 9918 16478
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 10050 16450 10064 16478
rect 9904 15694 10064 16450
rect 9904 15666 9918 15694
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 10050 15666 10064 15694
rect 9904 14910 10064 15666
rect 9904 14882 9918 14910
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 10050 14882 10064 14910
rect 9904 14126 10064 14882
rect 9904 14098 9918 14126
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 10050 14098 10064 14126
rect 9904 13342 10064 14098
rect 9904 13314 9918 13342
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 10050 13314 10064 13342
rect 9904 12558 10064 13314
rect 9904 12530 9918 12558
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 10050 12530 10064 12558
rect 9904 11774 10064 12530
rect 9904 11746 9918 11774
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 10050 11746 10064 11774
rect 2224 11354 2238 11382
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2370 11354 2384 11382
rect 2224 10598 2384 11354
rect 2224 10570 2238 10598
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2370 10570 2384 10598
rect 2224 9814 2384 10570
rect 2224 9786 2238 9814
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2370 9786 2384 9814
rect 2224 9030 2384 9786
rect 8078 11690 8106 11695
rect 8078 9226 8106 11662
rect 9904 10990 10064 11746
rect 9904 10962 9918 10990
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 10050 10962 10064 10990
rect 9904 10206 10064 10962
rect 9904 10178 9918 10206
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 10050 10178 10064 10206
rect 8078 9193 8106 9198
rect 9198 10122 9226 10127
rect 9198 9114 9226 10094
rect 9198 9081 9226 9086
rect 9904 9422 10064 10178
rect 9904 9394 9918 9422
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 10050 9394 10064 9422
rect 2224 9002 2238 9030
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2370 9002 2384 9030
rect 2224 8246 2384 9002
rect 2224 8218 2238 8246
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2370 8218 2384 8246
rect 2224 7462 2384 8218
rect 2224 7434 2238 7462
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2370 7434 2384 7462
rect 2224 6678 2384 7434
rect 2224 6650 2238 6678
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2370 6650 2384 6678
rect 2224 5894 2384 6650
rect 2224 5866 2238 5894
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2370 5866 2384 5894
rect 2224 5110 2384 5866
rect 2224 5082 2238 5110
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2370 5082 2384 5110
rect 2224 4326 2384 5082
rect 2224 4298 2238 4326
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2370 4298 2384 4326
rect 2224 3542 2384 4298
rect 2224 3514 2238 3542
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2370 3514 2384 3542
rect 2224 2758 2384 3514
rect 2224 2730 2238 2758
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2370 2730 2384 2758
rect 2224 1974 2384 2730
rect 2224 1946 2238 1974
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2370 1946 2384 1974
rect 2224 1538 2384 1946
rect 9904 8638 10064 9394
rect 9904 8610 9918 8638
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 10050 8610 10064 8638
rect 9904 7854 10064 8610
rect 9904 7826 9918 7854
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 10050 7826 10064 7854
rect 9904 7070 10064 7826
rect 9904 7042 9918 7070
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 10050 7042 10064 7070
rect 9904 6286 10064 7042
rect 9904 6258 9918 6286
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 10050 6258 10064 6286
rect 9904 5502 10064 6258
rect 9904 5474 9918 5502
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 10050 5474 10064 5502
rect 9904 4718 10064 5474
rect 9904 4690 9918 4718
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 10050 4690 10064 4718
rect 9904 3934 10064 4690
rect 9904 3906 9918 3934
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 10050 3906 10064 3934
rect 9904 3150 10064 3906
rect 9904 3122 9918 3150
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 10050 3122 10064 3150
rect 9904 2366 10064 3122
rect 9904 2338 9918 2366
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 10050 2338 10064 2366
rect 9904 1582 10064 2338
rect 9904 1554 9918 1582
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 10050 1554 10064 1582
rect 9904 1538 10064 1554
rect 17584 19222 17744 19238
rect 17584 19194 17598 19222
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17730 19194 17744 19222
rect 17584 18438 17744 19194
rect 17584 18410 17598 18438
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17730 18410 17744 18438
rect 17584 17654 17744 18410
rect 17584 17626 17598 17654
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17730 17626 17744 17654
rect 17584 16870 17744 17626
rect 17584 16842 17598 16870
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17730 16842 17744 16870
rect 17584 16086 17744 16842
rect 17584 16058 17598 16086
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17730 16058 17744 16086
rect 17584 15302 17744 16058
rect 17584 15274 17598 15302
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17730 15274 17744 15302
rect 17584 14518 17744 15274
rect 17584 14490 17598 14518
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17730 14490 17744 14518
rect 17584 13734 17744 14490
rect 17584 13706 17598 13734
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17730 13706 17744 13734
rect 17584 12950 17744 13706
rect 17584 12922 17598 12950
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17730 12922 17744 12950
rect 17584 12166 17744 12922
rect 17584 12138 17598 12166
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17730 12138 17744 12166
rect 17584 11382 17744 12138
rect 17584 11354 17598 11382
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17730 11354 17744 11382
rect 17584 10598 17744 11354
rect 17584 10570 17598 10598
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17730 10570 17744 10598
rect 17584 9814 17744 10570
rect 17584 9786 17598 9814
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17730 9786 17744 9814
rect 17584 9030 17744 9786
rect 17584 9002 17598 9030
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17730 9002 17744 9030
rect 17584 8246 17744 9002
rect 17584 8218 17598 8246
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17730 8218 17744 8246
rect 17584 7462 17744 8218
rect 17584 7434 17598 7462
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17730 7434 17744 7462
rect 17584 6678 17744 7434
rect 17584 6650 17598 6678
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17730 6650 17744 6678
rect 17584 5894 17744 6650
rect 17584 5866 17598 5894
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17730 5866 17744 5894
rect 17584 5110 17744 5866
rect 17584 5082 17598 5110
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17730 5082 17744 5110
rect 17584 4326 17744 5082
rect 17584 4298 17598 4326
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17730 4298 17744 4326
rect 17584 3542 17744 4298
rect 17584 3514 17598 3542
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17730 3514 17744 3542
rect 17584 2758 17744 3514
rect 17584 2730 17598 2758
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17730 2730 17744 2758
rect 17584 1974 17744 2730
rect 17584 1946 17598 1974
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17730 1946 17744 1974
rect 17584 1538 17744 1946
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _118_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 8008 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _119_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 7504 0 -1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _120_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 11032 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _121_
timestamp 1698175906
transform 1 0 6664 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _122_
timestamp 1698175906
transform 1 0 7392 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _123_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 7896 0 -1 10192
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _124_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 8792 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _125_
timestamp 1698175906
transform 1 0 10248 0 -1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _126_
timestamp 1698175906
transform -1 0 7504 0 -1 8624
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _127_
timestamp 1698175906
transform 1 0 7280 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _128_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8624 0 -1 10976
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _129_
timestamp 1698175906
transform -1 0 14784 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _130_
timestamp 1698175906
transform 1 0 8792 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _131_
timestamp 1698175906
transform 1 0 6888 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _132_
timestamp 1698175906
transform 1 0 10136 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _133_
timestamp 1698175906
transform -1 0 12040 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _134_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 11816 0 1 9408
box -43 -43 883 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _135_
timestamp 1698175906
transform 1 0 13832 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _136_
timestamp 1698175906
transform -1 0 13832 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _137_
timestamp 1698175906
transform -1 0 13496 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _138_
timestamp 1698175906
transform 1 0 7224 0 1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _139_
timestamp 1698175906
transform 1 0 7560 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _140_
timestamp 1698175906
transform -1 0 8176 0 -1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _141_
timestamp 1698175906
transform -1 0 7280 0 1 8624
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _142_
timestamp 1698175906
transform 1 0 6720 0 1 8624
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _143_
timestamp 1698175906
transform -1 0 10472 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _144_
timestamp 1698175906
transform -1 0 11144 0 1 9408
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _145_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 6832 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _146_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 8288 0 -1 9408
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _147_
timestamp 1698175906
transform 1 0 7616 0 -1 10192
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _148_
timestamp 1698175906
transform 1 0 8176 0 -1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _149_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8624 0 -1 9408
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _150_
timestamp 1698175906
transform 1 0 9016 0 1 8624
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _151_
timestamp 1698175906
transform 1 0 9184 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _152_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 11816 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _153_
timestamp 1698175906
transform 1 0 12040 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _154_
timestamp 1698175906
transform 1 0 12152 0 -1 10192
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _155_
timestamp 1698175906
transform 1 0 10920 0 -1 10976
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _156_
timestamp 1698175906
transform -1 0 9968 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _157_
timestamp 1698175906
transform 1 0 8176 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _158_
timestamp 1698175906
transform 1 0 9856 0 -1 13328
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _159_
timestamp 1698175906
transform -1 0 13104 0 -1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _160_
timestamp 1698175906
transform -1 0 12824 0 -1 12544
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _161_
timestamp 1698175906
transform 1 0 10472 0 -1 10976
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _162_
timestamp 1698175906
transform -1 0 9688 0 -1 12544
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _163_
timestamp 1698175906
transform -1 0 7560 0 1 11760
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _164_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 7504 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _165_
timestamp 1698175906
transform -1 0 8456 0 1 8624
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _166_
timestamp 1698175906
transform 1 0 8344 0 1 9408
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _167_
timestamp 1698175906
transform 1 0 10080 0 -1 11760
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _168_
timestamp 1698175906
transform -1 0 13160 0 1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _169_
timestamp 1698175906
transform -1 0 12096 0 -1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _170_
timestamp 1698175906
transform 1 0 8792 0 -1 10192
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _171_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 10192 0 -1 10976
box -43 -43 771 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _172_
timestamp 1698175906
transform -1 0 11256 0 1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _173_
timestamp 1698175906
transform -1 0 11144 0 1 12544
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _174_
timestamp 1698175906
transform -1 0 9520 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _175_
timestamp 1698175906
transform 1 0 7784 0 1 9408
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _176_
timestamp 1698175906
transform -1 0 8512 0 -1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _177_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 7952 0 1 12544
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _178_
timestamp 1698175906
transform 1 0 7224 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _179_
timestamp 1698175906
transform -1 0 7896 0 1 10976
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _180_
timestamp 1698175906
transform -1 0 7784 0 -1 10976
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _181_
timestamp 1698175906
transform -1 0 13272 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _182_
timestamp 1698175906
transform 1 0 7896 0 -1 10976
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _183_
timestamp 1698175906
transform 1 0 9800 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _184_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 10472 0 1 10976
box -43 -43 883 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _185_
timestamp 1698175906
transform 1 0 11200 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _186_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 7448 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _187_
timestamp 1698175906
transform -1 0 8008 0 -1 12544
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _188_
timestamp 1698175906
transform 1 0 6776 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _189_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 11144 0 -1 9408
box -43 -43 1331 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _190_
timestamp 1698175906
transform 1 0 13720 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _191_
timestamp 1698175906
transform 1 0 11200 0 1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _192_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 12992 0 1 8624
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _193_
timestamp 1698175906
transform 1 0 10584 0 1 8624
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _194_
timestamp 1698175906
transform 1 0 11256 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _195_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 11704 0 -1 7840
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _196_
timestamp 1698175906
transform -1 0 11144 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _197_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 12544 0 -1 10976
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _198_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 11704 0 -1 10976
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _199_
timestamp 1698175906
transform -1 0 13888 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _200_
timestamp 1698175906
transform 1 0 10192 0 -1 10976
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _201_
timestamp 1698175906
transform 1 0 13272 0 1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _202_
timestamp 1698175906
transform -1 0 13888 0 1 12544
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _203_
timestamp 1698175906
transform -1 0 12320 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _204_
timestamp 1698175906
transform 1 0 11368 0 -1 7056
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _205_
timestamp 1698175906
transform -1 0 9688 0 1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _206_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 9632 0 1 9408
box -43 -43 771 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _207_
timestamp 1698175906
transform 1 0 10024 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _208_
timestamp 1698175906
transform 1 0 9576 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _209_
timestamp 1698175906
transform -1 0 7504 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _210_
timestamp 1698175906
transform -1 0 7392 0 1 9408
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _211_
timestamp 1698175906
transform 1 0 9520 0 1 11760
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _212_
timestamp 1698175906
transform 1 0 9576 0 -1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _213_
timestamp 1698175906
transform 1 0 9744 0 1 12544
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _214_
timestamp 1698175906
transform -1 0 9744 0 -1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _215_
timestamp 1698175906
transform 1 0 8792 0 -1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _216_
timestamp 1698175906
transform 1 0 9072 0 -1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _217_
timestamp 1698175906
transform 1 0 8904 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _218_
timestamp 1698175906
transform 1 0 7896 0 1 10976
box -43 -43 1331 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _219_
timestamp 1698175906
transform -1 0 9464 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _220_
timestamp 1698175906
transform 1 0 9072 0 1 7056
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _221_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 9128 0 -1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _222_
timestamp 1698175906
transform -1 0 8512 0 -1 7056
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _223_
timestamp 1698175906
transform 1 0 9520 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _224_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 10920 0 -1 8624
box -43 -43 995 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _225_
timestamp 1698175906
transform 1 0 12544 0 -1 10192
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _226_
timestamp 1698175906
transform -1 0 13384 0 1 7840
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _227_
timestamp 1698175906
transform -1 0 13104 0 1 7840
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _228_
timestamp 1698175906
transform -1 0 13664 0 1 7840
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _229_
timestamp 1698175906
transform 1 0 7336 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _230_
timestamp 1698175906
transform 1 0 9800 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _231_
timestamp 1698175906
transform 1 0 11928 0 -1 7840
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _232_
timestamp 1698175906
transform -1 0 13440 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _233_
timestamp 1698175906
transform 1 0 11928 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _234_
timestamp 1698175906
transform -1 0 12880 0 -1 11760
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _235_
timestamp 1698175906
transform 1 0 12488 0 1 10976
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _236_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 13496 0 -1 10192
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _237_
timestamp 1698175906
transform 1 0 5488 0 -1 7840
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _238_
timestamp 1698175906
transform 1 0 6664 0 1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _239_
timestamp 1698175906
transform 1 0 4928 0 -1 9408
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _240_
timestamp 1698175906
transform 1 0 10696 0 1 10976
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _241_
timestamp 1698175906
transform 1 0 11984 0 1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _242_
timestamp 1698175906
transform -1 0 7224 0 -1 11760
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _243_
timestamp 1698175906
transform 1 0 11256 0 1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _244_
timestamp 1698175906
transform 1 0 10192 0 -1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _245_
timestamp 1698175906
transform -1 0 8176 0 -1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _246_
timestamp 1698175906
transform -1 0 7280 0 -1 10976
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _247_
timestamp 1698175906
transform -1 0 7504 0 -1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _248_
timestamp 1698175906
transform 1 0 13048 0 -1 9408
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _249_
timestamp 1698175906
transform 1 0 10584 0 1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _250_
timestamp 1698175906
transform 1 0 13216 0 -1 10976
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _251_
timestamp 1698175906
transform 1 0 13104 0 -1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _252_
timestamp 1698175906
transform 1 0 11144 0 1 6272
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _253_
timestamp 1698175906
transform 1 0 9128 0 -1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _254_
timestamp 1698175906
transform -1 0 6552 0 1 9408
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _255_
timestamp 1698175906
transform 1 0 8848 0 1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _256_
timestamp 1698175906
transform 1 0 7952 0 1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _257_
timestamp 1698175906
transform 1 0 7616 0 1 6272
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _258_
timestamp 1698175906
transform 1 0 12712 0 -1 7840
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _259_
timestamp 1698175906
transform 1 0 12544 0 1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _260_
timestamp 1698175906
transform 1 0 12880 0 -1 11760
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _264_
timestamp 1698175906
transform -1 0 10920 0 1 13328
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _265_
timestamp 1698175906
transform 1 0 14728 0 -1 13328
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__217__A1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9800 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__226__A2
timestamp 1698175906
transform 1 0 12992 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__228__A2
timestamp 1698175906
transform 1 0 13776 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__235__B2
timestamp 1698175906
transform 1 0 12376 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__236__CLK
timestamp 1698175906
transform 1 0 13048 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__237__CLK
timestamp 1698175906
transform 1 0 7224 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__238__CLK
timestamp 1698175906
transform 1 0 8400 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__239__CLK
timestamp 1698175906
transform 1 0 6440 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__240__CLK
timestamp 1698175906
transform 1 0 12320 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__241__CLK
timestamp 1698175906
transform 1 0 14000 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__242__CLK
timestamp 1698175906
transform 1 0 7336 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__243__CLK
timestamp 1698175906
transform -1 0 12992 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__244__CLK
timestamp 1698175906
transform 1 0 12208 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__245__CLK
timestamp 1698175906
transform 1 0 8288 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__246__CLK
timestamp 1698175906
transform 1 0 7280 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__247__CLK
timestamp 1698175906
transform 1 0 7672 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__248__CLK
timestamp 1698175906
transform 1 0 12936 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__249__CLK
timestamp 1698175906
transform 1 0 12320 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__250__CLK
timestamp 1698175906
transform 1 0 13384 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__251__CLK
timestamp 1698175906
transform 1 0 12712 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__252__CLK
timestamp 1698175906
transform -1 0 12992 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__253__CLK
timestamp 1698175906
transform 1 0 8960 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__254__CLK
timestamp 1698175906
transform 1 0 6552 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__255__CLK
timestamp 1698175906
transform 1 0 8736 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__256__CLK
timestamp 1698175906
transform 1 0 10360 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__257__CLK
timestamp 1698175906
transform -1 0 9688 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__258__CLK
timestamp 1698175906
transform 1 0 14448 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__259__CLK
timestamp 1698175906
transform 1 0 14280 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__260__CLK
timestamp 1698175906
transform 1 0 14616 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1698175906
transform 1 0 9296 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9352 0 -1 10192
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1698175906
transform -1 0 10248 0 1 10192
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1698175906
transform 1 0 11088 0 1 10192
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 784 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698175906
transform 1 0 2688 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698175906
transform 1 0 4592 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698175906
transform 1 0 6496 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_138 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8400 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_142 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8624 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_172
timestamp 1698175906
transform 1 0 10304 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_174 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10416 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_201
timestamp 1698175906
transform 1 0 11928 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_203
timestamp 1698175906
transform 1 0 12040 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_232
timestamp 1698175906
transform 1 0 13664 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_236
timestamp 1698175906
transform 1 0 13888 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_240
timestamp 1698175906
transform 1 0 14112 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_274 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 16016 0 1 1568
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_290 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 16912 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_298
timestamp 1698175906
transform 1 0 17360 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_300
timestamp 1698175906
transform 1 0 17472 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_305
timestamp 1698175906
transform 1 0 17752 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_308
timestamp 1698175906
transform 1 0 17920 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_342
timestamp 1698175906
transform 1 0 19824 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_346
timestamp 1698175906
transform 1 0 20048 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_348
timestamp 1698175906
transform 1 0 20160 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 784 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698175906
transform 1 0 4368 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698175906
transform 1 0 4704 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698175906
transform 1 0 8288 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_142
timestamp 1698175906
transform 1 0 8624 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_206
timestamp 1698175906
transform 1 0 12208 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_238
timestamp 1698175906
transform 1 0 14000 0 -1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_270
timestamp 1698175906
transform 1 0 15792 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_278
timestamp 1698175906
transform 1 0 16240 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_282
timestamp 1698175906
transform 1 0 16464 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_346
timestamp 1698175906
transform 1 0 20048 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_348
timestamp 1698175906
transform 1 0 20160 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698175906
transform 1 0 784 0 1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698175906
transform 1 0 2576 0 1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698175906
transform 1 0 2744 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698175906
transform 1 0 6328 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_107
timestamp 1698175906
transform 1 0 6664 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_171
timestamp 1698175906
transform 1 0 10248 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_177
timestamp 1698175906
transform 1 0 10584 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_241
timestamp 1698175906
transform 1 0 14168 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698175906
transform 1 0 14504 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698175906
transform 1 0 18088 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_317
timestamp 1698175906
transform 1 0 18424 0 1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698175906
transform 1 0 784 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698175906
transform 1 0 4368 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698175906
transform 1 0 4704 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698175906
transform 1 0 8288 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_142
timestamp 1698175906
transform 1 0 8624 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_206
timestamp 1698175906
transform 1 0 12208 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_212
timestamp 1698175906
transform 1 0 12544 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_276
timestamp 1698175906
transform 1 0 16128 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_282
timestamp 1698175906
transform 1 0 16464 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_346
timestamp 1698175906
transform 1 0 20048 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_348
timestamp 1698175906
transform 1 0 20160 0 -1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698175906
transform 1 0 784 0 1 3136
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698175906
transform 1 0 2576 0 1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698175906
transform 1 0 2744 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698175906
transform 1 0 6328 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_107
timestamp 1698175906
transform 1 0 6664 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698175906
transform 1 0 10248 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_177
timestamp 1698175906
transform 1 0 10584 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_241
timestamp 1698175906
transform 1 0 14168 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698175906
transform 1 0 14504 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698175906
transform 1 0 18088 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_317
timestamp 1698175906
transform 1 0 18424 0 1 3136
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698175906
transform 1 0 784 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698175906
transform 1 0 4368 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698175906
transform 1 0 4704 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698175906
transform 1 0 8288 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_142
timestamp 1698175906
transform 1 0 8624 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_206
timestamp 1698175906
transform 1 0 12208 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_212
timestamp 1698175906
transform 1 0 12544 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698175906
transform 1 0 16128 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_282
timestamp 1698175906
transform 1 0 16464 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_346
timestamp 1698175906
transform 1 0 20048 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_348
timestamp 1698175906
transform 1 0 20160 0 -1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698175906
transform 1 0 784 0 1 3920
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698175906
transform 1 0 2576 0 1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698175906
transform 1 0 2744 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698175906
transform 1 0 6328 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_107
timestamp 1698175906
transform 1 0 6664 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_171
timestamp 1698175906
transform 1 0 10248 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_177
timestamp 1698175906
transform 1 0 10584 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_241
timestamp 1698175906
transform 1 0 14168 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_247
timestamp 1698175906
transform 1 0 14504 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_311
timestamp 1698175906
transform 1 0 18088 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_317
timestamp 1698175906
transform 1 0 18424 0 1 3920
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698175906
transform 1 0 784 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698175906
transform 1 0 4368 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_72
timestamp 1698175906
transform 1 0 4704 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698175906
transform 1 0 8288 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_142
timestamp 1698175906
transform 1 0 8624 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_206
timestamp 1698175906
transform 1 0 12208 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_212
timestamp 1698175906
transform 1 0 12544 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_276
timestamp 1698175906
transform 1 0 16128 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_282
timestamp 1698175906
transform 1 0 16464 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_346
timestamp 1698175906
transform 1 0 20048 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_348
timestamp 1698175906
transform 1 0 20160 0 -1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698175906
transform 1 0 784 0 1 4704
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698175906
transform 1 0 2576 0 1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_37
timestamp 1698175906
transform 1 0 2744 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_101
timestamp 1698175906
transform 1 0 6328 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_107
timestamp 1698175906
transform 1 0 6664 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_171
timestamp 1698175906
transform 1 0 10248 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_177
timestamp 1698175906
transform 1 0 10584 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_241
timestamp 1698175906
transform 1 0 14168 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_247
timestamp 1698175906
transform 1 0 14504 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_311
timestamp 1698175906
transform 1 0 18088 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_317
timestamp 1698175906
transform 1 0 18424 0 1 4704
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698175906
transform 1 0 784 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698175906
transform 1 0 4368 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_72
timestamp 1698175906
transform 1 0 4704 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_136
timestamp 1698175906
transform 1 0 8288 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_142
timestamp 1698175906
transform 1 0 8624 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_206
timestamp 1698175906
transform 1 0 12208 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_212
timestamp 1698175906
transform 1 0 12544 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_276
timestamp 1698175906
transform 1 0 16128 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_282
timestamp 1698175906
transform 1 0 16464 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_346
timestamp 1698175906
transform 1 0 20048 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_348
timestamp 1698175906
transform 1 0 20160 0 -1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698175906
transform 1 0 784 0 1 5488
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698175906
transform 1 0 2576 0 1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_37
timestamp 1698175906
transform 1 0 2744 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698175906
transform 1 0 6328 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_107
timestamp 1698175906
transform 1 0 6664 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_171
timestamp 1698175906
transform 1 0 10248 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_177
timestamp 1698175906
transform 1 0 10584 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_241
timestamp 1698175906
transform 1 0 14168 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_247
timestamp 1698175906
transform 1 0 14504 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_311
timestamp 1698175906
transform 1 0 18088 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_317
timestamp 1698175906
transform 1 0 18424 0 1 5488
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2
timestamp 1698175906
transform 1 0 784 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698175906
transform 1 0 4368 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_72
timestamp 1698175906
transform 1 0 4704 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698175906
transform 1 0 8288 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_142
timestamp 1698175906
transform 1 0 8624 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_206
timestamp 1698175906
transform 1 0 12208 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_212
timestamp 1698175906
transform 1 0 12544 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_276
timestamp 1698175906
transform 1 0 16128 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_282
timestamp 1698175906
transform 1 0 16464 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_346
timestamp 1698175906
transform 1 0 20048 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_348
timestamp 1698175906
transform 1 0 20160 0 -1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698175906
transform 1 0 784 0 1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698175906
transform 1 0 2576 0 1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_37
timestamp 1698175906
transform 1 0 2744 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698175906
transform 1 0 6328 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_107
timestamp 1698175906
transform 1 0 6664 0 1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_123
timestamp 1698175906
transform 1 0 7560 0 1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_157
timestamp 1698175906
transform 1 0 9464 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_161
timestamp 1698175906
transform 1 0 9688 0 1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_169
timestamp 1698175906
transform 1 0 10136 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_173
timestamp 1698175906
transform 1 0 10360 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_177
timestamp 1698175906
transform 1 0 10584 0 1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_185
timestamp 1698175906
transform 1 0 11032 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_216
timestamp 1698175906
transform 1 0 12768 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_220
timestamp 1698175906
transform 1 0 12992 0 1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_236
timestamp 1698175906
transform 1 0 13888 0 1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_244
timestamp 1698175906
transform 1 0 14336 0 1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_247
timestamp 1698175906
transform 1 0 14504 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_311
timestamp 1698175906
transform 1 0 18088 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_317
timestamp 1698175906
transform 1 0 18424 0 1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_2
timestamp 1698175906
transform 1 0 784 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_66
timestamp 1698175906
transform 1 0 4368 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_72
timestamp 1698175906
transform 1 0 4704 0 -1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_104
timestamp 1698175906
transform 1 0 6496 0 -1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_120
timestamp 1698175906
transform 1 0 7392 0 -1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_128
timestamp 1698175906
transform 1 0 7840 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_132
timestamp 1698175906
transform 1 0 8064 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_142
timestamp 1698175906
transform 1 0 8624 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_180
timestamp 1698175906
transform 1 0 10752 0 -1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_188
timestamp 1698175906
transform 1 0 11200 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_190
timestamp 1698175906
transform 1 0 11312 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_201
timestamp 1698175906
transform 1 0 11928 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_203
timestamp 1698175906
transform 1 0 12040 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_208
timestamp 1698175906
transform 1 0 12320 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_212
timestamp 1698175906
transform 1 0 12544 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_276
timestamp 1698175906
transform 1 0 16128 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_282
timestamp 1698175906
transform 1 0 16464 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_346
timestamp 1698175906
transform 1 0 20048 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_348
timestamp 1698175906
transform 1 0 20160 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698175906
transform 1 0 784 0 1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698175906
transform 1 0 2576 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_37
timestamp 1698175906
transform 1 0 2744 0 1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_101
timestamp 1698175906
transform 1 0 6328 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_136
timestamp 1698175906
transform 1 0 8288 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_140
timestamp 1698175906
transform 1 0 8512 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_206
timestamp 1698175906
transform 1 0 12208 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_210
timestamp 1698175906
transform 1 0 12432 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_241
timestamp 1698175906
transform 1 0 14168 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_247
timestamp 1698175906
transform 1 0 14504 0 1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_311
timestamp 1698175906
transform 1 0 18088 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_317
timestamp 1698175906
transform 1 0 18424 0 1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_2
timestamp 1698175906
transform 1 0 784 0 -1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_66
timestamp 1698175906
transform 1 0 4368 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_72
timestamp 1698175906
transform 1 0 4704 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_80
timestamp 1698175906
transform 1 0 5152 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_84
timestamp 1698175906
transform 1 0 5376 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_115
timestamp 1698175906
transform 1 0 7112 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_119
timestamp 1698175906
transform 1 0 7336 0 -1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_135
timestamp 1698175906
transform 1 0 8232 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_139
timestamp 1698175906
transform 1 0 8456 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_142
timestamp 1698175906
transform 1 0 8624 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_150
timestamp 1698175906
transform 1 0 9072 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_154
timestamp 1698175906
transform 1 0 9296 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_162
timestamp 1698175906
transform 1 0 9744 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_170
timestamp 1698175906
transform 1 0 10192 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_177
timestamp 1698175906
transform 1 0 10584 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_197
timestamp 1698175906
transform 1 0 11704 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_212
timestamp 1698175906
transform 1 0 12544 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_214
timestamp 1698175906
transform 1 0 12656 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_244
timestamp 1698175906
transform 1 0 14336 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_248
timestamp 1698175906
transform 1 0 14560 0 -1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_282
timestamp 1698175906
transform 1 0 16464 0 -1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_314
timestamp 1698175906
transform 1 0 18256 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_322
timestamp 1698175906
transform 1 0 18704 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_2
timestamp 1698175906
transform 1 0 784 0 1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698175906
transform 1 0 2576 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_37
timestamp 1698175906
transform 1 0 2744 0 1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_101
timestamp 1698175906
transform 1 0 6328 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_107
timestamp 1698175906
transform 1 0 6664 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_115
timestamp 1698175906
transform 1 0 7112 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_131
timestamp 1698175906
transform 1 0 8008 0 1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_147
timestamp 1698175906
transform 1 0 8904 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_161
timestamp 1698175906
transform 1 0 9688 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_169
timestamp 1698175906
transform 1 0 10136 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_173
timestamp 1698175906
transform 1 0 10360 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_177
timestamp 1698175906
transform 1 0 10584 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_185
timestamp 1698175906
transform 1 0 11032 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_187
timestamp 1698175906
transform 1 0 11144 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_194
timestamp 1698175906
transform 1 0 11536 0 1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_210
timestamp 1698175906
transform 1 0 12432 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_212
timestamp 1698175906
transform 1 0 12544 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_232
timestamp 1698175906
transform 1 0 13664 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_236
timestamp 1698175906
transform 1 0 13888 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_244
timestamp 1698175906
transform 1 0 14336 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_247
timestamp 1698175906
transform 1 0 14504 0 1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_311
timestamp 1698175906
transform 1 0 18088 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_317
timestamp 1698175906
transform 1 0 18424 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_321
timestamp 1698175906
transform 1 0 18648 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_2
timestamp 1698175906
transform 1 0 784 0 -1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_66
timestamp 1698175906
transform 1 0 4368 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_72
timestamp 1698175906
transform 1 0 4704 0 -1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_104
timestamp 1698175906
transform 1 0 6496 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_112
timestamp 1698175906
transform 1 0 6944 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_116
timestamp 1698175906
transform 1 0 7168 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_142
timestamp 1698175906
transform 1 0 8624 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_144
timestamp 1698175906
transform 1 0 8736 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_153
timestamp 1698175906
transform 1 0 9240 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_161
timestamp 1698175906
transform 1 0 9688 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_165
timestamp 1698175906
transform 1 0 9912 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_183
timestamp 1698175906
transform 1 0 10920 0 -1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_199
timestamp 1698175906
transform 1 0 11816 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_207
timestamp 1698175906
transform 1 0 12264 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_209
timestamp 1698175906
transform 1 0 12376 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_212
timestamp 1698175906
transform 1 0 12544 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_222
timestamp 1698175906
transform 1 0 13104 0 -1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_254
timestamp 1698175906
transform 1 0 14896 0 -1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_270
timestamp 1698175906
transform 1 0 15792 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_278
timestamp 1698175906
transform 1 0 16240 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_282
timestamp 1698175906
transform 1 0 16464 0 -1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_346
timestamp 1698175906
transform 1 0 20048 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_348
timestamp 1698175906
transform 1 0 20160 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_2
timestamp 1698175906
transform 1 0 784 0 1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698175906
transform 1 0 2576 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_37
timestamp 1698175906
transform 1 0 2744 0 1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_101
timestamp 1698175906
transform 1 0 6328 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_107
timestamp 1698175906
transform 1 0 6664 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_126
timestamp 1698175906
transform 1 0 7728 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_128
timestamp 1698175906
transform 1 0 7840 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_145
timestamp 1698175906
transform 1 0 8792 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_154
timestamp 1698175906
transform 1 0 9296 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_162
timestamp 1698175906
transform 1 0 9744 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_171
timestamp 1698175906
transform 1 0 10248 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_182
timestamp 1698175906
transform 1 0 10864 0 1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_214
timestamp 1698175906
transform 1 0 12656 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_218
timestamp 1698175906
transform 1 0 12880 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_230
timestamp 1698175906
transform 1 0 13552 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_232
timestamp 1698175906
transform 1 0 13664 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_239
timestamp 1698175906
transform 1 0 14056 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_243
timestamp 1698175906
transform 1 0 14280 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_247
timestamp 1698175906
transform 1 0 14504 0 1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_311
timestamp 1698175906
transform 1 0 18088 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_317
timestamp 1698175906
transform 1 0 18424 0 1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_2
timestamp 1698175906
transform 1 0 784 0 -1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_66
timestamp 1698175906
transform 1 0 4368 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_72
timestamp 1698175906
transform 1 0 4704 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_105
timestamp 1698175906
transform 1 0 6552 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_117
timestamp 1698175906
transform 1 0 7224 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_136
timestamp 1698175906
transform 1 0 8288 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_149
timestamp 1698175906
transform 1 0 9016 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_151
timestamp 1698175906
transform 1 0 9128 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_187
timestamp 1698175906
transform 1 0 11144 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_209
timestamp 1698175906
transform 1 0 12376 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_212
timestamp 1698175906
transform 1 0 12544 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_216
timestamp 1698175906
transform 1 0 12768 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_218
timestamp 1698175906
transform 1 0 12880 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_250
timestamp 1698175906
transform 1 0 14672 0 -1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_266
timestamp 1698175906
transform 1 0 15568 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_274
timestamp 1698175906
transform 1 0 16016 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_278
timestamp 1698175906
transform 1 0 16240 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_282
timestamp 1698175906
transform 1 0 16464 0 -1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_314
timestamp 1698175906
transform 1 0 18256 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_322
timestamp 1698175906
transform 1 0 18704 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_28
timestamp 1698175906
transform 1 0 2240 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_32
timestamp 1698175906
transform 1 0 2464 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698175906
transform 1 0 2576 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_37
timestamp 1698175906
transform 1 0 2744 0 1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_69
timestamp 1698175906
transform 1 0 4536 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_73
timestamp 1698175906
transform 1 0 4760 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_75
timestamp 1698175906
transform 1 0 4872 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_107
timestamp 1698175906
transform 1 0 6664 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_109
timestamp 1698175906
transform 1 0 6776 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_126
timestamp 1698175906
transform 1 0 7728 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_166
timestamp 1698175906
transform 1 0 9968 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_168
timestamp 1698175906
transform 1 0 10080 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_187
timestamp 1698175906
transform 1 0 11144 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_214
timestamp 1698175906
transform 1 0 12656 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_218
timestamp 1698175906
transform 1 0 12880 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_220
timestamp 1698175906
transform 1 0 12992 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_241
timestamp 1698175906
transform 1 0 14168 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_247
timestamp 1698175906
transform 1 0 14504 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_252
timestamp 1698175906
transform 1 0 14784 0 1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_284
timestamp 1698175906
transform 1 0 16576 0 1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_300
timestamp 1698175906
transform 1 0 17472 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_308
timestamp 1698175906
transform 1 0 17920 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_312
timestamp 1698175906
transform 1 0 18144 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_314
timestamp 1698175906
transform 1 0 18256 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_317
timestamp 1698175906
transform 1 0 18424 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_321
timestamp 1698175906
transform 1 0 18648 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_2
timestamp 1698175906
transform 1 0 784 0 -1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_66
timestamp 1698175906
transform 1 0 4368 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_72
timestamp 1698175906
transform 1 0 4704 0 -1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_104
timestamp 1698175906
transform 1 0 6496 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_107
timestamp 1698175906
transform 1 0 6664 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_109
timestamp 1698175906
transform 1 0 6776 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_122
timestamp 1698175906
transform 1 0 7504 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_142
timestamp 1698175906
transform 1 0 8624 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_144
timestamp 1698175906
transform 1 0 8736 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_225
timestamp 1698175906
transform 1 0 13272 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_258
timestamp 1698175906
transform 1 0 15120 0 -1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_274
timestamp 1698175906
transform 1 0 16016 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_278
timestamp 1698175906
transform 1 0 16240 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_282
timestamp 1698175906
transform 1 0 16464 0 -1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_346
timestamp 1698175906
transform 1 0 20048 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_348
timestamp 1698175906
transform 1 0 20160 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_2
timestamp 1698175906
transform 1 0 784 0 1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698175906
transform 1 0 2576 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_37
timestamp 1698175906
transform 1 0 2744 0 1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_101
timestamp 1698175906
transform 1 0 6328 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_107
timestamp 1698175906
transform 1 0 6664 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_115
timestamp 1698175906
transform 1 0 7112 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_117
timestamp 1698175906
transform 1 0 7224 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_120
timestamp 1698175906
transform 1 0 7392 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_185
timestamp 1698175906
transform 1 0 11032 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_236
timestamp 1698175906
transform 1 0 13888 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_244
timestamp 1698175906
transform 1 0 14336 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_247
timestamp 1698175906
transform 1 0 14504 0 1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_311
timestamp 1698175906
transform 1 0 18088 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_317
timestamp 1698175906
transform 1 0 18424 0 1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_2
timestamp 1698175906
transform 1 0 784 0 -1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_66
timestamp 1698175906
transform 1 0 4368 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_72
timestamp 1698175906
transform 1 0 4704 0 -1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_88
timestamp 1698175906
transform 1 0 5600 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_118
timestamp 1698175906
transform 1 0 7280 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_127
timestamp 1698175906
transform 1 0 7784 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_152
timestamp 1698175906
transform 1 0 9184 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_156
timestamp 1698175906
transform 1 0 9408 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_180
timestamp 1698175906
transform 1 0 10752 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_182
timestamp 1698175906
transform 1 0 10864 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_196
timestamp 1698175906
transform 1 0 11648 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_206
timestamp 1698175906
transform 1 0 12208 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_222
timestamp 1698175906
transform 1 0 13104 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_253
timestamp 1698175906
transform 1 0 14840 0 -1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_269
timestamp 1698175906
transform 1 0 15736 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_277
timestamp 1698175906
transform 1 0 16184 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_279
timestamp 1698175906
transform 1 0 16296 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_282
timestamp 1698175906
transform 1 0 16464 0 -1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_346
timestamp 1698175906
transform 1 0 20048 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_348
timestamp 1698175906
transform 1 0 20160 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_28
timestamp 1698175906
transform 1 0 2240 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_32
timestamp 1698175906
transform 1 0 2464 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698175906
transform 1 0 2576 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_37
timestamp 1698175906
transform 1 0 2744 0 1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_101
timestamp 1698175906
transform 1 0 6328 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_107
timestamp 1698175906
transform 1 0 6664 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_111
timestamp 1698175906
transform 1 0 6888 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_113
timestamp 1698175906
transform 1 0 7000 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_122
timestamp 1698175906
transform 1 0 7504 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_158
timestamp 1698175906
transform 1 0 9520 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_177
timestamp 1698175906
transform 1 0 10584 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_208
timestamp 1698175906
transform 1 0 12320 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_210
timestamp 1698175906
transform 1 0 12432 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_236
timestamp 1698175906
transform 1 0 13888 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_244
timestamp 1698175906
transform 1 0 14336 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_247
timestamp 1698175906
transform 1 0 14504 0 1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_311
timestamp 1698175906
transform 1 0 18088 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_317
timestamp 1698175906
transform 1 0 18424 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_321
timestamp 1698175906
transform 1 0 18648 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_2
timestamp 1698175906
transform 1 0 784 0 -1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_66
timestamp 1698175906
transform 1 0 4368 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_72
timestamp 1698175906
transform 1 0 4704 0 -1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_117
timestamp 1698175906
transform 1 0 7224 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_129
timestamp 1698175906
transform 1 0 7896 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_137
timestamp 1698175906
transform 1 0 8344 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_139
timestamp 1698175906
transform 1 0 8456 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_142
timestamp 1698175906
transform 1 0 8624 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_144
timestamp 1698175906
transform 1 0 8736 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_151
timestamp 1698175906
transform 1 0 9128 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_159
timestamp 1698175906
transform 1 0 9576 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_167
timestamp 1698175906
transform 1 0 10024 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_173
timestamp 1698175906
transform 1 0 10360 0 -1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_189
timestamp 1698175906
transform 1 0 11256 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_197
timestamp 1698175906
transform 1 0 11704 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_209
timestamp 1698175906
transform 1 0 12376 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_212
timestamp 1698175906
transform 1 0 12544 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_247
timestamp 1698175906
transform 1 0 14504 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_251
timestamp 1698175906
transform 1 0 14728 0 -1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_267
timestamp 1698175906
transform 1 0 15624 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_275
timestamp 1698175906
transform 1 0 16072 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_279
timestamp 1698175906
transform 1 0 16296 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_282
timestamp 1698175906
transform 1 0 16464 0 -1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_314
timestamp 1698175906
transform 1 0 18256 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_322
timestamp 1698175906
transform 1 0 18704 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_28
timestamp 1698175906
transform 1 0 2240 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_32
timestamp 1698175906
transform 1 0 2464 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698175906
transform 1 0 2576 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_37
timestamp 1698175906
transform 1 0 2744 0 1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_101
timestamp 1698175906
transform 1 0 6328 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_107
timestamp 1698175906
transform 1 0 6664 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_115
timestamp 1698175906
transform 1 0 7112 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_117
timestamp 1698175906
transform 1 0 7224 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_123
timestamp 1698175906
transform 1 0 7560 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_127
timestamp 1698175906
transform 1 0 7784 0 1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_143
timestamp 1698175906
transform 1 0 8680 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_151
timestamp 1698175906
transform 1 0 9128 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_155
timestamp 1698175906
transform 1 0 9352 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_157
timestamp 1698175906
transform 1 0 9464 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_163
timestamp 1698175906
transform 1 0 9800 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_171
timestamp 1698175906
transform 1 0 10248 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_177
timestamp 1698175906
transform 1 0 10584 0 1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_211
timestamp 1698175906
transform 1 0 12488 0 1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_243
timestamp 1698175906
transform 1 0 14280 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_247
timestamp 1698175906
transform 1 0 14504 0 1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_311
timestamp 1698175906
transform 1 0 18088 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_317
timestamp 1698175906
transform 1 0 18424 0 1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_2
timestamp 1698175906
transform 1 0 784 0 -1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_66
timestamp 1698175906
transform 1 0 4368 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_72
timestamp 1698175906
transform 1 0 4704 0 -1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_88
timestamp 1698175906
transform 1 0 5600 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_92
timestamp 1698175906
transform 1 0 5824 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_131
timestamp 1698175906
transform 1 0 8008 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_139
timestamp 1698175906
transform 1 0 8456 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_142
timestamp 1698175906
transform 1 0 8624 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_146
timestamp 1698175906
transform 1 0 8848 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_161
timestamp 1698175906
transform 1 0 9688 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_165
timestamp 1698175906
transform 1 0 9912 0 -1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_197
timestamp 1698175906
transform 1 0 11704 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_205
timestamp 1698175906
transform 1 0 12152 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_209
timestamp 1698175906
transform 1 0 12376 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_217
timestamp 1698175906
transform 1 0 12824 0 -1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_249
timestamp 1698175906
transform 1 0 14616 0 -1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_265
timestamp 1698175906
transform 1 0 15512 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_273
timestamp 1698175906
transform 1 0 15960 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_277
timestamp 1698175906
transform 1 0 16184 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_279
timestamp 1698175906
transform 1 0 16296 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_282
timestamp 1698175906
transform 1 0 16464 0 -1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_346
timestamp 1698175906
transform 1 0 20048 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_348
timestamp 1698175906
transform 1 0 20160 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_2
timestamp 1698175906
transform 1 0 784 0 1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698175906
transform 1 0 2576 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_37
timestamp 1698175906
transform 1 0 2744 0 1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_101
timestamp 1698175906
transform 1 0 6328 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_107
timestamp 1698175906
transform 1 0 6664 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_113
timestamp 1698175906
transform 1 0 7000 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_159
timestamp 1698175906
transform 1 0 9576 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_161
timestamp 1698175906
transform 1 0 9688 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_171
timestamp 1698175906
transform 1 0 10248 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_177
timestamp 1698175906
transform 1 0 10584 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_181
timestamp 1698175906
transform 1 0 10808 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_187
timestamp 1698175906
transform 1 0 11144 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_195
timestamp 1698175906
transform 1 0 11592 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_199
timestamp 1698175906
transform 1 0 11816 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_201
timestamp 1698175906
transform 1 0 11928 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_236
timestamp 1698175906
transform 1 0 13888 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_240
timestamp 1698175906
transform 1 0 14112 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_244
timestamp 1698175906
transform 1 0 14336 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_247
timestamp 1698175906
transform 1 0 14504 0 1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_311
timestamp 1698175906
transform 1 0 18088 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_317
timestamp 1698175906
transform 1 0 18424 0 1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_28
timestamp 1698175906
transform 1 0 2240 0 -1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_60
timestamp 1698175906
transform 1 0 4032 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_68
timestamp 1698175906
transform 1 0 4480 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_72
timestamp 1698175906
transform 1 0 4704 0 -1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_104
timestamp 1698175906
transform 1 0 6496 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_134
timestamp 1698175906
transform 1 0 8176 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_138
timestamp 1698175906
transform 1 0 8400 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_142
timestamp 1698175906
transform 1 0 8624 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_155
timestamp 1698175906
transform 1 0 9352 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_204
timestamp 1698175906
transform 1 0 12096 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_208
timestamp 1698175906
transform 1 0 12320 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_212
timestamp 1698175906
transform 1 0 12544 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_214
timestamp 1698175906
transform 1 0 12656 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_257
timestamp 1698175906
transform 1 0 15064 0 -1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_273
timestamp 1698175906
transform 1 0 15960 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_277
timestamp 1698175906
transform 1 0 16184 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_279
timestamp 1698175906
transform 1 0 16296 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_282
timestamp 1698175906
transform 1 0 16464 0 -1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_314
timestamp 1698175906
transform 1 0 18256 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_322
timestamp 1698175906
transform 1 0 18704 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_28
timestamp 1698175906
transform 1 0 2240 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_32
timestamp 1698175906
transform 1 0 2464 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698175906
transform 1 0 2576 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_37
timestamp 1698175906
transform 1 0 2744 0 1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_101
timestamp 1698175906
transform 1 0 6328 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_107
timestamp 1698175906
transform 1 0 6664 0 1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_139
timestamp 1698175906
transform 1 0 8456 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_143
timestamp 1698175906
transform 1 0 8680 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_183
timestamp 1698175906
transform 1 0 10920 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_223
timestamp 1698175906
transform 1 0 13160 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_230
timestamp 1698175906
transform 1 0 13552 0 1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_238
timestamp 1698175906
transform 1 0 14000 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_242
timestamp 1698175906
transform 1 0 14224 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_244
timestamp 1698175906
transform 1 0 14336 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_247
timestamp 1698175906
transform 1 0 14504 0 1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_311
timestamp 1698175906
transform 1 0 18088 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_317
timestamp 1698175906
transform 1 0 18424 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_321
timestamp 1698175906
transform 1 0 18648 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_2
timestamp 1698175906
transform 1 0 784 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_66
timestamp 1698175906
transform 1 0 4368 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_72
timestamp 1698175906
transform 1 0 4704 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_136
timestamp 1698175906
transform 1 0 8288 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_142
timestamp 1698175906
transform 1 0 8624 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_206
timestamp 1698175906
transform 1 0 12208 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_212
timestamp 1698175906
transform 1 0 12544 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_216
timestamp 1698175906
transform 1 0 12768 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_220
timestamp 1698175906
transform 1 0 12992 0 -1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_252
timestamp 1698175906
transform 1 0 14784 0 -1 14112
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_268
timestamp 1698175906
transform 1 0 15680 0 -1 14112
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_276
timestamp 1698175906
transform 1 0 16128 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_282
timestamp 1698175906
transform 1 0 16464 0 -1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_314
timestamp 1698175906
transform 1 0 18256 0 -1 14112
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_322
timestamp 1698175906
transform 1 0 18704 0 -1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_2
timestamp 1698175906
transform 1 0 784 0 1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698175906
transform 1 0 2576 0 1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_37
timestamp 1698175906
transform 1 0 2744 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_101
timestamp 1698175906
transform 1 0 6328 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_107
timestamp 1698175906
transform 1 0 6664 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_171
timestamp 1698175906
transform 1 0 10248 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_177
timestamp 1698175906
transform 1 0 10584 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_241
timestamp 1698175906
transform 1 0 14168 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_247
timestamp 1698175906
transform 1 0 14504 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_311
timestamp 1698175906
transform 1 0 18088 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_317
timestamp 1698175906
transform 1 0 18424 0 1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_2
timestamp 1698175906
transform 1 0 784 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_66
timestamp 1698175906
transform 1 0 4368 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_72
timestamp 1698175906
transform 1 0 4704 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_136
timestamp 1698175906
transform 1 0 8288 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_142
timestamp 1698175906
transform 1 0 8624 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_206
timestamp 1698175906
transform 1 0 12208 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_212
timestamp 1698175906
transform 1 0 12544 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_276
timestamp 1698175906
transform 1 0 16128 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_282
timestamp 1698175906
transform 1 0 16464 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_346
timestamp 1698175906
transform 1 0 20048 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_348
timestamp 1698175906
transform 1 0 20160 0 -1 14896
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698175906
transform 1 0 784 0 1 14896
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698175906
transform 1 0 2576 0 1 14896
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_37
timestamp 1698175906
transform 1 0 2744 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_101
timestamp 1698175906
transform 1 0 6328 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_107
timestamp 1698175906
transform 1 0 6664 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_171
timestamp 1698175906
transform 1 0 10248 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_177
timestamp 1698175906
transform 1 0 10584 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_241
timestamp 1698175906
transform 1 0 14168 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_247
timestamp 1698175906
transform 1 0 14504 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_311
timestamp 1698175906
transform 1 0 18088 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_317
timestamp 1698175906
transform 1 0 18424 0 1 14896
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2
timestamp 1698175906
transform 1 0 784 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_66
timestamp 1698175906
transform 1 0 4368 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_72
timestamp 1698175906
transform 1 0 4704 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_136
timestamp 1698175906
transform 1 0 8288 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_142
timestamp 1698175906
transform 1 0 8624 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_206
timestamp 1698175906
transform 1 0 12208 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_212
timestamp 1698175906
transform 1 0 12544 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_276
timestamp 1698175906
transform 1 0 16128 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_282
timestamp 1698175906
transform 1 0 16464 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_346
timestamp 1698175906
transform 1 0 20048 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_348
timestamp 1698175906
transform 1 0 20160 0 -1 15680
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_2
timestamp 1698175906
transform 1 0 784 0 1 15680
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698175906
transform 1 0 2576 0 1 15680
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_37
timestamp 1698175906
transform 1 0 2744 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_101
timestamp 1698175906
transform 1 0 6328 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_107
timestamp 1698175906
transform 1 0 6664 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_171
timestamp 1698175906
transform 1 0 10248 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_177
timestamp 1698175906
transform 1 0 10584 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_241
timestamp 1698175906
transform 1 0 14168 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_247
timestamp 1698175906
transform 1 0 14504 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_311
timestamp 1698175906
transform 1 0 18088 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_317
timestamp 1698175906
transform 1 0 18424 0 1 15680
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2
timestamp 1698175906
transform 1 0 784 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_66
timestamp 1698175906
transform 1 0 4368 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_72
timestamp 1698175906
transform 1 0 4704 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_136
timestamp 1698175906
transform 1 0 8288 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_142
timestamp 1698175906
transform 1 0 8624 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_206
timestamp 1698175906
transform 1 0 12208 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_212
timestamp 1698175906
transform 1 0 12544 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_276
timestamp 1698175906
transform 1 0 16128 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_282
timestamp 1698175906
transform 1 0 16464 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_346
timestamp 1698175906
transform 1 0 20048 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_348
timestamp 1698175906
transform 1 0 20160 0 -1 16464
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698175906
transform 1 0 784 0 1 16464
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698175906
transform 1 0 2576 0 1 16464
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_37
timestamp 1698175906
transform 1 0 2744 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_101
timestamp 1698175906
transform 1 0 6328 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_107
timestamp 1698175906
transform 1 0 6664 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_171
timestamp 1698175906
transform 1 0 10248 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_177
timestamp 1698175906
transform 1 0 10584 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_241
timestamp 1698175906
transform 1 0 14168 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_247
timestamp 1698175906
transform 1 0 14504 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_311
timestamp 1698175906
transform 1 0 18088 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_317
timestamp 1698175906
transform 1 0 18424 0 1 16464
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_2
timestamp 1698175906
transform 1 0 784 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_66
timestamp 1698175906
transform 1 0 4368 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_72
timestamp 1698175906
transform 1 0 4704 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_136
timestamp 1698175906
transform 1 0 8288 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_142
timestamp 1698175906
transform 1 0 8624 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_206
timestamp 1698175906
transform 1 0 12208 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_212
timestamp 1698175906
transform 1 0 12544 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_276
timestamp 1698175906
transform 1 0 16128 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_282
timestamp 1698175906
transform 1 0 16464 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_346
timestamp 1698175906
transform 1 0 20048 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_348
timestamp 1698175906
transform 1 0 20160 0 -1 17248
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698175906
transform 1 0 784 0 1 17248
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698175906
transform 1 0 2576 0 1 17248
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_37
timestamp 1698175906
transform 1 0 2744 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_101
timestamp 1698175906
transform 1 0 6328 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_107
timestamp 1698175906
transform 1 0 6664 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_171
timestamp 1698175906
transform 1 0 10248 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_177
timestamp 1698175906
transform 1 0 10584 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_241
timestamp 1698175906
transform 1 0 14168 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_247
timestamp 1698175906
transform 1 0 14504 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_311
timestamp 1698175906
transform 1 0 18088 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_317
timestamp 1698175906
transform 1 0 18424 0 1 17248
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_333
timestamp 1698175906
transform 1 0 19320 0 1 17248
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_341
timestamp 1698175906
transform 1 0 19768 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2
timestamp 1698175906
transform 1 0 784 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1698175906
transform 1 0 4368 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_72
timestamp 1698175906
transform 1 0 4704 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_136
timestamp 1698175906
transform 1 0 8288 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_142
timestamp 1698175906
transform 1 0 8624 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_206
timestamp 1698175906
transform 1 0 12208 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_212
timestamp 1698175906
transform 1 0 12544 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_276
timestamp 1698175906
transform 1 0 16128 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_282
timestamp 1698175906
transform 1 0 16464 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_346
timestamp 1698175906
transform 1 0 20048 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_348
timestamp 1698175906
transform 1 0 20160 0 -1 18032
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_2
timestamp 1698175906
transform 1 0 784 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698175906
transform 1 0 2576 0 1 18032
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_37
timestamp 1698175906
transform 1 0 2744 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_101
timestamp 1698175906
transform 1 0 6328 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_107
timestamp 1698175906
transform 1 0 6664 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_171
timestamp 1698175906
transform 1 0 10248 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_177
timestamp 1698175906
transform 1 0 10584 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_241
timestamp 1698175906
transform 1 0 14168 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_247
timestamp 1698175906
transform 1 0 14504 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_311
timestamp 1698175906
transform 1 0 18088 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_317
timestamp 1698175906
transform 1 0 18424 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_2
timestamp 1698175906
transform 1 0 784 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_66
timestamp 1698175906
transform 1 0 4368 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_72
timestamp 1698175906
transform 1 0 4704 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_136
timestamp 1698175906
transform 1 0 8288 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_142
timestamp 1698175906
transform 1 0 8624 0 -1 18816
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_158
timestamp 1698175906
transform 1 0 9520 0 -1 18816
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_166
timestamp 1698175906
transform 1 0 9968 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_168
timestamp 1698175906
transform 1 0 10080 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_195
timestamp 1698175906
transform 1 0 11592 0 -1 18816
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_203
timestamp 1698175906
transform 1 0 12040 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_207
timestamp 1698175906
transform 1 0 12264 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_209
timestamp 1698175906
transform 1 0 12376 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_212
timestamp 1698175906
transform 1 0 12544 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_216
timestamp 1698175906
transform 1 0 12768 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_243
timestamp 1698175906
transform 1 0 14280 0 -1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_275
timestamp 1698175906
transform 1 0 16072 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_279
timestamp 1698175906
transform 1 0 16296 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_282
timestamp 1698175906
transform 1 0 16464 0 -1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_314
timestamp 1698175906
transform 1 0 18256 0 -1 18816
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_330
timestamp 1698175906
transform 1 0 19152 0 -1 18816
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_338
timestamp 1698175906
transform 1 0 19600 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_342
timestamp 1698175906
transform 1 0 19824 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_344
timestamp 1698175906
transform 1 0 19936 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_2
timestamp 1698175906
transform 1 0 784 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_36
timestamp 1698175906
transform 1 0 2688 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_70
timestamp 1698175906
transform 1 0 4592 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_104
timestamp 1698175906
transform 1 0 6496 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_138
timestamp 1698175906
transform 1 0 8400 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_142
timestamp 1698175906
transform 1 0 8624 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_172
timestamp 1698175906
transform 1 0 10304 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_174
timestamp 1698175906
transform 1 0 10416 0 1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_201
timestamp 1698175906
transform 1 0 11928 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_203
timestamp 1698175906
transform 1 0 12040 0 1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_232
timestamp 1698175906
transform 1 0 13664 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_236
timestamp 1698175906
transform 1 0 13888 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_240
timestamp 1698175906
transform 1 0 14112 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_274
timestamp 1698175906
transform 1 0 16016 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_308
timestamp 1698175906
transform 1 0 17920 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_342
timestamp 1698175906
transform 1 0 19824 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_346
timestamp 1698175906
transform 1 0 20048 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_348
timestamp 1698175906
transform 1 0 20160 0 1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita30_24 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19992 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita30_25
timestamp 1698175906
transform -1 0 17752 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita30_26
timestamp 1698175906
transform 1 0 19992 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8736 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output2
timestamp 1698175906
transform 1 0 18760 0 1 7840
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output3
timestamp 1698175906
transform 1 0 18760 0 -1 7840
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output4
timestamp 1698175906
transform 1 0 18760 0 -1 11760
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output5
timestamp 1698175906
transform 1 0 10472 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output6
timestamp 1698175906
transform 1 0 18760 0 -1 13328
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output7
timestamp 1698175906
transform 1 0 10136 0 -1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output8
timestamp 1698175906
transform 1 0 8736 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output9
timestamp 1698175906
transform 1 0 18760 0 -1 9408
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output10
timestamp 1698175906
transform 1 0 12208 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output11
timestamp 1698175906
transform 1 0 18760 0 1 10976
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output12
timestamp 1698175906
transform -1 0 2240 0 -1 13328
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output13
timestamp 1698175906
transform 1 0 10472 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output14
timestamp 1698175906
transform -1 0 2240 0 1 9408
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output15
timestamp 1698175906
transform -1 0 2240 0 1 10976
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output16
timestamp 1698175906
transform -1 0 2240 0 1 13328
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output17
timestamp 1698175906
transform 1 0 12208 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output18
timestamp 1698175906
transform 1 0 12824 0 -1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output19
timestamp 1698175906
transform -1 0 2240 0 1 11760
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output20
timestamp 1698175906
transform 1 0 18760 0 1 13328
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output21
timestamp 1698175906
transform 1 0 18760 0 -1 14112
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output22
timestamp 1698175906
transform 1 0 12544 0 -1 2352
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output23
timestamp 1698175906
transform 1 0 18760 0 1 9408
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_45 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 672 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698175906
transform -1 0 20328 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_46
timestamp 1698175906
transform 1 0 672 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698175906
transform -1 0 20328 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_47
timestamp 1698175906
transform 1 0 672 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698175906
transform -1 0 20328 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_48
timestamp 1698175906
transform 1 0 672 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698175906
transform -1 0 20328 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_49
timestamp 1698175906
transform 1 0 672 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698175906
transform -1 0 20328 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_50
timestamp 1698175906
transform 1 0 672 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698175906
transform -1 0 20328 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_51
timestamp 1698175906
transform 1 0 672 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698175906
transform -1 0 20328 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_52
timestamp 1698175906
transform 1 0 672 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698175906
transform -1 0 20328 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_53
timestamp 1698175906
transform 1 0 672 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698175906
transform -1 0 20328 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_54
timestamp 1698175906
transform 1 0 672 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698175906
transform -1 0 20328 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_55
timestamp 1698175906
transform 1 0 672 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698175906
transform -1 0 20328 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_56
timestamp 1698175906
transform 1 0 672 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698175906
transform -1 0 20328 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_57
timestamp 1698175906
transform 1 0 672 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698175906
transform -1 0 20328 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_58
timestamp 1698175906
transform 1 0 672 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698175906
transform -1 0 20328 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_59
timestamp 1698175906
transform 1 0 672 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698175906
transform -1 0 20328 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_60
timestamp 1698175906
transform 1 0 672 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698175906
transform -1 0 20328 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_61
timestamp 1698175906
transform 1 0 672 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698175906
transform -1 0 20328 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_62
timestamp 1698175906
transform 1 0 672 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698175906
transform -1 0 20328 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_63
timestamp 1698175906
transform 1 0 672 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698175906
transform -1 0 20328 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_64
timestamp 1698175906
transform 1 0 672 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698175906
transform -1 0 20328 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_65
timestamp 1698175906
transform 1 0 672 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698175906
transform -1 0 20328 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_66
timestamp 1698175906
transform 1 0 672 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698175906
transform -1 0 20328 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_67
timestamp 1698175906
transform 1 0 672 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698175906
transform -1 0 20328 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_68
timestamp 1698175906
transform 1 0 672 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698175906
transform -1 0 20328 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_69
timestamp 1698175906
transform 1 0 672 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698175906
transform -1 0 20328 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_70
timestamp 1698175906
transform 1 0 672 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698175906
transform -1 0 20328 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_71
timestamp 1698175906
transform 1 0 672 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698175906
transform -1 0 20328 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_72
timestamp 1698175906
transform 1 0 672 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698175906
transform -1 0 20328 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_73
timestamp 1698175906
transform 1 0 672 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698175906
transform -1 0 20328 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_74
timestamp 1698175906
transform 1 0 672 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698175906
transform -1 0 20328 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_75
timestamp 1698175906
transform 1 0 672 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698175906
transform -1 0 20328 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_76
timestamp 1698175906
transform 1 0 672 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698175906
transform -1 0 20328 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_77
timestamp 1698175906
transform 1 0 672 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698175906
transform -1 0 20328 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_78
timestamp 1698175906
transform 1 0 672 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698175906
transform -1 0 20328 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_79
timestamp 1698175906
transform 1 0 672 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698175906
transform -1 0 20328 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_80
timestamp 1698175906
transform 1 0 672 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698175906
transform -1 0 20328 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_81
timestamp 1698175906
transform 1 0 672 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698175906
transform -1 0 20328 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_82
timestamp 1698175906
transform 1 0 672 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698175906
transform -1 0 20328 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_83
timestamp 1698175906
transform 1 0 672 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698175906
transform -1 0 20328 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_84
timestamp 1698175906
transform 1 0 672 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698175906
transform -1 0 20328 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_85
timestamp 1698175906
transform 1 0 672 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698175906
transform -1 0 20328 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_86
timestamp 1698175906
transform 1 0 672 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698175906
transform -1 0 20328 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_87
timestamp 1698175906
transform 1 0 672 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698175906
transform -1 0 20328 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_88
timestamp 1698175906
transform 1 0 672 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698175906
transform -1 0 20328 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_89
timestamp 1698175906
transform 1 0 672 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698175906
transform -1 0 20328 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_90 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 2576 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_91
timestamp 1698175906
transform 1 0 4480 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_92
timestamp 1698175906
transform 1 0 6384 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_93
timestamp 1698175906
transform 1 0 8288 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_94
timestamp 1698175906
transform 1 0 10192 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_95
timestamp 1698175906
transform 1 0 12096 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_96
timestamp 1698175906
transform 1 0 14000 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_97
timestamp 1698175906
transform 1 0 15904 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_98
timestamp 1698175906
transform 1 0 17808 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_99
timestamp 1698175906
transform 1 0 19712 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_100
timestamp 1698175906
transform 1 0 4592 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_101
timestamp 1698175906
transform 1 0 8512 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_102
timestamp 1698175906
transform 1 0 12432 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_103
timestamp 1698175906
transform 1 0 16352 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_104
timestamp 1698175906
transform 1 0 2632 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_105
timestamp 1698175906
transform 1 0 6552 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_106
timestamp 1698175906
transform 1 0 10472 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_107
timestamp 1698175906
transform 1 0 14392 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_108
timestamp 1698175906
transform 1 0 18312 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_109
timestamp 1698175906
transform 1 0 4592 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_110
timestamp 1698175906
transform 1 0 8512 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_111
timestamp 1698175906
transform 1 0 12432 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_112
timestamp 1698175906
transform 1 0 16352 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_113
timestamp 1698175906
transform 1 0 2632 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_114
timestamp 1698175906
transform 1 0 6552 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_115
timestamp 1698175906
transform 1 0 10472 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_116
timestamp 1698175906
transform 1 0 14392 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_117
timestamp 1698175906
transform 1 0 18312 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_118
timestamp 1698175906
transform 1 0 4592 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_119
timestamp 1698175906
transform 1 0 8512 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_120
timestamp 1698175906
transform 1 0 12432 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_121
timestamp 1698175906
transform 1 0 16352 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_122
timestamp 1698175906
transform 1 0 2632 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_123
timestamp 1698175906
transform 1 0 6552 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_124
timestamp 1698175906
transform 1 0 10472 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_125
timestamp 1698175906
transform 1 0 14392 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_126
timestamp 1698175906
transform 1 0 18312 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_127
timestamp 1698175906
transform 1 0 4592 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_128
timestamp 1698175906
transform 1 0 8512 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_129
timestamp 1698175906
transform 1 0 12432 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_130
timestamp 1698175906
transform 1 0 16352 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_131
timestamp 1698175906
transform 1 0 2632 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_132
timestamp 1698175906
transform 1 0 6552 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_133
timestamp 1698175906
transform 1 0 10472 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_134
timestamp 1698175906
transform 1 0 14392 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_135
timestamp 1698175906
transform 1 0 18312 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_136
timestamp 1698175906
transform 1 0 4592 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_137
timestamp 1698175906
transform 1 0 8512 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_138
timestamp 1698175906
transform 1 0 12432 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_139
timestamp 1698175906
transform 1 0 16352 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_140
timestamp 1698175906
transform 1 0 2632 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_141
timestamp 1698175906
transform 1 0 6552 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_142
timestamp 1698175906
transform 1 0 10472 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_143
timestamp 1698175906
transform 1 0 14392 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_144
timestamp 1698175906
transform 1 0 18312 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_145
timestamp 1698175906
transform 1 0 4592 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_146
timestamp 1698175906
transform 1 0 8512 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_147
timestamp 1698175906
transform 1 0 12432 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_148
timestamp 1698175906
transform 1 0 16352 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_149
timestamp 1698175906
transform 1 0 2632 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_150
timestamp 1698175906
transform 1 0 6552 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_151
timestamp 1698175906
transform 1 0 10472 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_152
timestamp 1698175906
transform 1 0 14392 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_153
timestamp 1698175906
transform 1 0 18312 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_154
timestamp 1698175906
transform 1 0 4592 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_155
timestamp 1698175906
transform 1 0 8512 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_156
timestamp 1698175906
transform 1 0 12432 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_157
timestamp 1698175906
transform 1 0 16352 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_158
timestamp 1698175906
transform 1 0 2632 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_159
timestamp 1698175906
transform 1 0 6552 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_160
timestamp 1698175906
transform 1 0 10472 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_161
timestamp 1698175906
transform 1 0 14392 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_162
timestamp 1698175906
transform 1 0 18312 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_163
timestamp 1698175906
transform 1 0 4592 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_164
timestamp 1698175906
transform 1 0 8512 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_165
timestamp 1698175906
transform 1 0 12432 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_166
timestamp 1698175906
transform 1 0 16352 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_167
timestamp 1698175906
transform 1 0 2632 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_168
timestamp 1698175906
transform 1 0 6552 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_169
timestamp 1698175906
transform 1 0 10472 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_170
timestamp 1698175906
transform 1 0 14392 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_171
timestamp 1698175906
transform 1 0 18312 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_172
timestamp 1698175906
transform 1 0 4592 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_173
timestamp 1698175906
transform 1 0 8512 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_174
timestamp 1698175906
transform 1 0 12432 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_175
timestamp 1698175906
transform 1 0 16352 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_176
timestamp 1698175906
transform 1 0 2632 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_177
timestamp 1698175906
transform 1 0 6552 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_178
timestamp 1698175906
transform 1 0 10472 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_179
timestamp 1698175906
transform 1 0 14392 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_180
timestamp 1698175906
transform 1 0 18312 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_181
timestamp 1698175906
transform 1 0 4592 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_182
timestamp 1698175906
transform 1 0 8512 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_183
timestamp 1698175906
transform 1 0 12432 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_184
timestamp 1698175906
transform 1 0 16352 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_185
timestamp 1698175906
transform 1 0 2632 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_186
timestamp 1698175906
transform 1 0 6552 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_187
timestamp 1698175906
transform 1 0 10472 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_188
timestamp 1698175906
transform 1 0 14392 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_189
timestamp 1698175906
transform 1 0 18312 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_190
timestamp 1698175906
transform 1 0 4592 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_191
timestamp 1698175906
transform 1 0 8512 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_192
timestamp 1698175906
transform 1 0 12432 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_193
timestamp 1698175906
transform 1 0 16352 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_194
timestamp 1698175906
transform 1 0 2632 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_195
timestamp 1698175906
transform 1 0 6552 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_196
timestamp 1698175906
transform 1 0 10472 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_197
timestamp 1698175906
transform 1 0 14392 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_198
timestamp 1698175906
transform 1 0 18312 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_199
timestamp 1698175906
transform 1 0 4592 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_200
timestamp 1698175906
transform 1 0 8512 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_201
timestamp 1698175906
transform 1 0 12432 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_202
timestamp 1698175906
transform 1 0 16352 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_203
timestamp 1698175906
transform 1 0 2632 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_204
timestamp 1698175906
transform 1 0 6552 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_205
timestamp 1698175906
transform 1 0 10472 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_206
timestamp 1698175906
transform 1 0 14392 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_207
timestamp 1698175906
transform 1 0 18312 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_208
timestamp 1698175906
transform 1 0 4592 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_209
timestamp 1698175906
transform 1 0 8512 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_210
timestamp 1698175906
transform 1 0 12432 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_211
timestamp 1698175906
transform 1 0 16352 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_212
timestamp 1698175906
transform 1 0 2632 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_213
timestamp 1698175906
transform 1 0 6552 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_214
timestamp 1698175906
transform 1 0 10472 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_215
timestamp 1698175906
transform 1 0 14392 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_216
timestamp 1698175906
transform 1 0 18312 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_217
timestamp 1698175906
transform 1 0 4592 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_218
timestamp 1698175906
transform 1 0 8512 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_219
timestamp 1698175906
transform 1 0 12432 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_220
timestamp 1698175906
transform 1 0 16352 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_221
timestamp 1698175906
transform 1 0 2632 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_222
timestamp 1698175906
transform 1 0 6552 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_223
timestamp 1698175906
transform 1 0 10472 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_224
timestamp 1698175906
transform 1 0 14392 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_225
timestamp 1698175906
transform 1 0 18312 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_226
timestamp 1698175906
transform 1 0 4592 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_227
timestamp 1698175906
transform 1 0 8512 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_228
timestamp 1698175906
transform 1 0 12432 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_229
timestamp 1698175906
transform 1 0 16352 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_230
timestamp 1698175906
transform 1 0 2632 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_231
timestamp 1698175906
transform 1 0 6552 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_232
timestamp 1698175906
transform 1 0 10472 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_233
timestamp 1698175906
transform 1 0 14392 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_234
timestamp 1698175906
transform 1 0 18312 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_235
timestamp 1698175906
transform 1 0 4592 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_236
timestamp 1698175906
transform 1 0 8512 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_237
timestamp 1698175906
transform 1 0 12432 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_238
timestamp 1698175906
transform 1 0 16352 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_239
timestamp 1698175906
transform 1 0 2632 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_240
timestamp 1698175906
transform 1 0 6552 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_241
timestamp 1698175906
transform 1 0 10472 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_242
timestamp 1698175906
transform 1 0 14392 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_243
timestamp 1698175906
transform 1 0 18312 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_244
timestamp 1698175906
transform 1 0 4592 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_245
timestamp 1698175906
transform 1 0 8512 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_246
timestamp 1698175906
transform 1 0 12432 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_247
timestamp 1698175906
transform 1 0 16352 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_248
timestamp 1698175906
transform 1 0 2632 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_249
timestamp 1698175906
transform 1 0 6552 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_250
timestamp 1698175906
transform 1 0 10472 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_251
timestamp 1698175906
transform 1 0 14392 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_252
timestamp 1698175906
transform 1 0 18312 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_253
timestamp 1698175906
transform 1 0 4592 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_254
timestamp 1698175906
transform 1 0 8512 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_255
timestamp 1698175906
transform 1 0 12432 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_256
timestamp 1698175906
transform 1 0 16352 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_257
timestamp 1698175906
transform 1 0 2632 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_258
timestamp 1698175906
transform 1 0 6552 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_259
timestamp 1698175906
transform 1 0 10472 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_260
timestamp 1698175906
transform 1 0 14392 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_261
timestamp 1698175906
transform 1 0 18312 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_262
timestamp 1698175906
transform 1 0 4592 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_263
timestamp 1698175906
transform 1 0 8512 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_264
timestamp 1698175906
transform 1 0 12432 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_265
timestamp 1698175906
transform 1 0 16352 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_266
timestamp 1698175906
transform 1 0 2632 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_267
timestamp 1698175906
transform 1 0 6552 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_268
timestamp 1698175906
transform 1 0 10472 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_269
timestamp 1698175906
transform 1 0 14392 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_270
timestamp 1698175906
transform 1 0 18312 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_271
timestamp 1698175906
transform 1 0 4592 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_272
timestamp 1698175906
transform 1 0 8512 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_273
timestamp 1698175906
transform 1 0 12432 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_274
timestamp 1698175906
transform 1 0 16352 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_275
timestamp 1698175906
transform 1 0 2632 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_276
timestamp 1698175906
transform 1 0 6552 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_277
timestamp 1698175906
transform 1 0 10472 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_278
timestamp 1698175906
transform 1 0 14392 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_279
timestamp 1698175906
transform 1 0 18312 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_280
timestamp 1698175906
transform 1 0 4592 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_281
timestamp 1698175906
transform 1 0 8512 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_282
timestamp 1698175906
transform 1 0 12432 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_283
timestamp 1698175906
transform 1 0 16352 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_284
timestamp 1698175906
transform 1 0 2632 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_285
timestamp 1698175906
transform 1 0 6552 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_286
timestamp 1698175906
transform 1 0 10472 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_287
timestamp 1698175906
transform 1 0 14392 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_288
timestamp 1698175906
transform 1 0 18312 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_289
timestamp 1698175906
transform 1 0 4592 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_290
timestamp 1698175906
transform 1 0 8512 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_291
timestamp 1698175906
transform 1 0 12432 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_292
timestamp 1698175906
transform 1 0 16352 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_293
timestamp 1698175906
transform 1 0 2576 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_294
timestamp 1698175906
transform 1 0 4480 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_295
timestamp 1698175906
transform 1 0 6384 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_296
timestamp 1698175906
transform 1 0 8288 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_297
timestamp 1698175906
transform 1 0 10192 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_298
timestamp 1698175906
transform 1 0 12096 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_299
timestamp 1698175906
transform 1 0 14000 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_300
timestamp 1698175906
transform 1 0 15904 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_301
timestamp 1698175906
transform 1 0 17808 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_302
timestamp 1698175906
transform 1 0 19712 0 1 18816
box -43 -43 155 435
<< labels >>
flabel metal3 s 0 13440 400 13496 0 FreeSans 224 0 0 0 clk
port 0 nsew signal input
flabel metal3 s 20600 18480 21000 18536 0 FreeSans 224 0 0 0 segm[0]
port 1 nsew signal tristate
flabel metal2 s 9072 0 9128 400 0 FreeSans 224 90 0 0 segm[10]
port 2 nsew signal tristate
flabel metal3 s 20600 7728 21000 7784 0 FreeSans 224 0 0 0 segm[11]
port 3 nsew signal tristate
flabel metal3 s 20600 7392 21000 7448 0 FreeSans 224 0 0 0 segm[12]
port 4 nsew signal tristate
flabel metal3 s 20600 11424 21000 11480 0 FreeSans 224 0 0 0 segm[13]
port 5 nsew signal tristate
flabel metal2 s 10416 20600 10472 21000 0 FreeSans 224 90 0 0 segm[1]
port 6 nsew signal tristate
flabel metal3 s 20600 12768 21000 12824 0 FreeSans 224 0 0 0 segm[2]
port 7 nsew signal tristate
flabel metal2 s 17472 0 17528 400 0 FreeSans 224 90 0 0 segm[3]
port 8 nsew signal tristate
flabel metal2 s 10080 20600 10136 21000 0 FreeSans 224 90 0 0 segm[4]
port 9 nsew signal tristate
flabel metal3 s 20600 17136 21000 17192 0 FreeSans 224 0 0 0 segm[5]
port 10 nsew signal tristate
flabel metal2 s 9408 20600 9464 21000 0 FreeSans 224 90 0 0 segm[6]
port 11 nsew signal tristate
flabel metal3 s 20600 9072 21000 9128 0 FreeSans 224 0 0 0 segm[7]
port 12 nsew signal tristate
flabel metal2 s 11424 0 11480 400 0 FreeSans 224 90 0 0 segm[8]
port 13 nsew signal tristate
flabel metal3 s 20600 11088 21000 11144 0 FreeSans 224 0 0 0 segm[9]
port 14 nsew signal tristate
flabel metal3 s 0 12768 400 12824 0 FreeSans 224 0 0 0 sel[0]
port 15 nsew signal tristate
flabel metal2 s 10416 0 10472 400 0 FreeSans 224 90 0 0 sel[10]
port 16 nsew signal tristate
flabel metal3 s 0 9408 400 9464 0 FreeSans 224 0 0 0 sel[11]
port 17 nsew signal tristate
flabel metal3 s 0 11088 400 11144 0 FreeSans 224 0 0 0 sel[1]
port 18 nsew signal tristate
flabel metal3 s 0 13104 400 13160 0 FreeSans 224 0 0 0 sel[2]
port 19 nsew signal tristate
flabel metal2 s 11424 20600 11480 21000 0 FreeSans 224 90 0 0 sel[3]
port 20 nsew signal tristate
flabel metal2 s 12768 20600 12824 21000 0 FreeSans 224 90 0 0 sel[4]
port 21 nsew signal tristate
flabel metal3 s 0 11760 400 11816 0 FreeSans 224 0 0 0 sel[5]
port 22 nsew signal tristate
flabel metal3 s 20600 13104 21000 13160 0 FreeSans 224 0 0 0 sel[6]
port 23 nsew signal tristate
flabel metal3 s 20600 13440 21000 13496 0 FreeSans 224 0 0 0 sel[7]
port 24 nsew signal tristate
flabel metal2 s 12432 0 12488 400 0 FreeSans 224 90 0 0 sel[8]
port 25 nsew signal tristate
flabel metal3 s 20600 9408 21000 9464 0 FreeSans 224 0 0 0 sel[9]
port 26 nsew signal tristate
flabel metal4 s 2224 1538 2384 19238 0 FreeSans 640 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 17584 1538 17744 19238 0 FreeSans 640 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 9904 1538 10064 19238 0 FreeSans 640 90 0 0 vss
port 28 nsew ground bidirectional
rlabel metal1 10500 19208 10500 19208 0 vdd
rlabel metal1 10500 18816 10500 18816 0 vss
rlabel metal3 7350 8764 7350 8764 0 _000_
rlabel metal2 6972 8596 6972 8596 0 _001_
rlabel metal3 7364 9156 7364 9156 0 _002_
rlabel metal2 11172 11004 11172 11004 0 _003_
rlabel metal2 12572 12572 12572 12572 0 _004_
rlabel metal3 7056 11060 7056 11060 0 _005_
rlabel metal2 11732 13454 11732 13454 0 _006_
rlabel metal2 10892 12908 10892 12908 0 _007_
rlabel metal3 7462 12684 7462 12684 0 _008_
rlabel metal2 6804 11172 6804 11172 0 _009_
rlabel metal2 7028 12516 7028 12516 0 _010_
rlabel metal2 13468 8932 13468 8932 0 _011_
rlabel metal2 11032 7308 11032 7308 0 _012_
rlabel metal2 13692 10948 13692 10948 0 _013_
rlabel metal2 13636 12908 13636 12908 0 _014_
rlabel metal2 11620 6748 11620 6748 0 _015_
rlabel metal2 9604 6944 9604 6944 0 _016_
rlabel metal2 6076 9520 6076 9520 0 _017_
rlabel metal2 10136 12852 10136 12852 0 _018_
rlabel metal2 9044 12572 9044 12572 0 _019_
rlabel metal2 8092 6720 8092 6720 0 _020_
rlabel metal2 13188 7728 13188 7728 0 _021_
rlabel metal3 12600 7308 12600 7308 0 _022_
rlabel metal2 12740 11004 12740 11004 0 _023_
rlabel metal2 13356 9800 13356 9800 0 _024_
rlabel metal3 11060 12740 11060 12740 0 _025_
rlabel metal3 12460 13524 12460 13524 0 _026_
rlabel metal2 9212 9576 9212 9576 0 _027_
rlabel metal2 10052 10864 10052 10864 0 _028_
rlabel metal2 11004 13076 11004 13076 0 _029_
rlabel metal2 8652 11144 8652 11144 0 _030_
rlabel metal2 10388 10836 10388 10836 0 _031_
rlabel metal2 7980 11928 7980 11928 0 _032_
rlabel metal2 7448 12796 7448 12796 0 _033_
rlabel metal2 7644 11368 7644 11368 0 _034_
rlabel metal2 7532 11144 7532 11144 0 _035_
rlabel metal2 12628 10444 12628 10444 0 _036_
rlabel metal2 11284 10724 11284 10724 0 _037_
rlabel metal2 10164 11368 10164 11368 0 _038_
rlabel metal2 11508 10976 11508 10976 0 _039_
rlabel metal2 11340 10668 11340 10668 0 _040_
rlabel metal2 6860 12600 6860 12600 0 _041_
rlabel metal2 13076 8932 13076 8932 0 _042_
rlabel metal3 13580 8820 13580 8820 0 _043_
rlabel metal3 13048 8036 13048 8036 0 _044_
rlabel metal2 10864 7700 10864 7700 0 _045_
rlabel metal2 11732 7154 11732 7154 0 _046_
rlabel metal2 11284 7532 11284 7532 0 _047_
rlabel metal2 13636 11060 13636 11060 0 _048_
rlabel metal3 13622 11172 13622 11172 0 _049_
rlabel metal2 13748 12208 13748 12208 0 _050_
rlabel metal2 13804 13076 13804 13076 0 _051_
rlabel metal3 11872 6860 11872 6860 0 _052_
rlabel metal2 9772 7336 9772 7336 0 _053_
rlabel metal2 9268 7392 9268 7392 0 _054_
rlabel metal3 9940 7168 9940 7168 0 _055_
rlabel metal2 7084 9800 7084 9800 0 _056_
rlabel metal2 9772 12292 9772 12292 0 _057_
rlabel metal2 9828 12936 9828 12936 0 _058_
rlabel metal3 13692 7980 13692 7980 0 _059_
rlabel metal2 8932 12012 8932 12012 0 _060_
rlabel metal2 9324 12740 9324 12740 0 _061_
rlabel metal2 9072 9324 9072 9324 0 _062_
rlabel metal2 9268 6580 9268 6580 0 _063_
rlabel metal3 9128 6860 9128 6860 0 _064_
rlabel metal3 8596 6860 8596 6860 0 _065_
rlabel metal2 10052 8400 10052 8400 0 _066_
rlabel metal2 10612 9156 10612 9156 0 _067_
rlabel metal2 12908 8960 12908 8960 0 _068_
rlabel metal2 13076 7980 13076 7980 0 _069_
rlabel metal2 12124 7840 12124 7840 0 _070_
rlabel metal2 7476 9044 7476 9044 0 _071_
rlabel metal3 10892 7700 10892 7700 0 _072_
rlabel metal3 12936 11060 12936 11060 0 _073_
rlabel metal3 12488 11172 12488 11172 0 _074_
rlabel metal2 12712 11172 12712 11172 0 _075_
rlabel metal2 7868 8288 7868 8288 0 _076_
rlabel metal2 7980 10948 7980 10948 0 _077_
rlabel metal3 9856 9996 9856 9996 0 _078_
rlabel metal2 6888 9996 6888 9996 0 _079_
rlabel metal2 8764 9576 8764 9576 0 _080_
rlabel metal2 8008 9884 8008 9884 0 _081_
rlabel metal3 10388 7224 10388 7224 0 _082_
rlabel metal2 13524 10612 13524 10612 0 _083_
rlabel metal2 7252 8568 7252 8568 0 _084_
rlabel metal2 8876 10276 8876 10276 0 _085_
rlabel metal2 10500 9380 10500 9380 0 _086_
rlabel metal3 14364 9604 14364 9604 0 _087_
rlabel metal2 9716 10472 9716 10472 0 _088_
rlabel metal2 7140 9184 7140 9184 0 _089_
rlabel metal2 12516 9800 12516 9800 0 _090_
rlabel metal3 11956 9324 11956 9324 0 _091_
rlabel metal2 13916 9352 13916 9352 0 _092_
rlabel metal2 13860 9660 13860 9660 0 _093_
rlabel metal2 13496 9660 13496 9660 0 _094_
rlabel metal2 7476 8036 7476 8036 0 _095_
rlabel metal2 7196 8736 7196 8736 0 _096_
rlabel metal2 7168 8932 7168 8932 0 _097_
rlabel metal3 10360 9604 10360 9604 0 _098_
rlabel metal2 9436 9184 9436 9184 0 _099_
rlabel metal3 7252 10052 7252 10052 0 _100_
rlabel metal2 7308 9688 7308 9688 0 _101_
rlabel metal2 9156 9324 9156 9324 0 _102_
rlabel metal2 8960 9324 8960 9324 0 _103_
rlabel metal3 10612 9212 10612 9212 0 _104_
rlabel metal2 9268 8960 9268 8960 0 _105_
rlabel metal3 12488 10892 12488 10892 0 _106_
rlabel metal2 12292 9184 12292 9184 0 _107_
rlabel metal2 12292 9912 12292 9912 0 _108_
rlabel metal2 7700 9408 7700 9408 0 _109_
rlabel metal2 9548 11620 9548 11620 0 _110_
rlabel metal3 10640 13468 10640 13468 0 _111_
rlabel metal2 12768 12404 12768 12404 0 _112_
rlabel metal2 7420 10864 7420 10864 0 _113_
rlabel metal2 7476 12236 7476 12236 0 _114_
rlabel metal2 7084 11508 7084 11508 0 _115_
rlabel metal3 9072 11676 9072 11676 0 _116_
rlabel metal2 9996 9296 9996 9296 0 _117_
rlabel metal3 1239 13468 1239 13468 0 clk
rlabel metal2 11172 10220 11172 10220 0 clknet_0_clk
rlabel metal2 8876 13468 8876 13468 0 clknet_1_0__leaf_clk
rlabel metal2 11396 13496 11396 13496 0 clknet_1_1__leaf_clk
rlabel metal2 7308 8260 7308 8260 0 dut30.count\[0\]
rlabel metal2 8204 7434 8204 7434 0 dut30.count\[1\]
rlabel metal2 6860 9212 6860 9212 0 dut30.count\[2\]
rlabel metal2 10892 10416 10892 10416 0 dut30.count\[3\]
rlabel metal3 8988 6524 8988 6524 0 net1
rlabel metal2 12292 2982 12292 2982 0 net10
rlabel metal2 14756 10752 14756 10752 0 net11
rlabel metal2 5964 12712 5964 12712 0 net12
rlabel metal2 10556 2982 10556 2982 0 net13
rlabel metal3 3178 9604 3178 9604 0 net14
rlabel metal2 2156 11004 2156 11004 0 net15
rlabel metal2 6636 13300 6636 13300 0 net16
rlabel metal2 11704 14140 11704 14140 0 net17
rlabel metal2 12796 13776 12796 13776 0 net18
rlabel metal2 5684 11732 5684 11732 0 net19
rlabel metal2 18956 7812 18956 7812 0 net2
rlabel metal3 15470 13188 15470 13188 0 net20
rlabel metal2 13524 12824 13524 12824 0 net21
rlabel metal2 12656 6524 12656 6524 0 net22
rlabel metal2 14700 9800 14700 9800 0 net23
rlabel metal2 20132 18592 20132 18592 0 net24
rlabel metal2 17500 1015 17500 1015 0 net25
rlabel metal2 20132 17248 20132 17248 0 net26
rlabel metal2 14084 7588 14084 7588 0 net3
rlabel metal3 15190 11508 15190 11508 0 net4
rlabel metal2 10668 16240 10668 16240 0 net5
rlabel metal2 14644 13272 14644 13272 0 net6
rlabel metal2 10388 16100 10388 16100 0 net7
rlabel metal2 9044 17486 9044 17486 0 net8
rlabel metal2 13972 8988 13972 8988 0 net9
rlabel metal2 9100 1099 9100 1099 0 segm[10]
rlabel metal2 20020 7924 20020 7924 0 segm[11]
rlabel metal2 20020 7504 20020 7504 0 segm[12]
rlabel metal3 20321 11452 20321 11452 0 segm[13]
rlabel metal2 10444 19873 10444 19873 0 segm[1]
rlabel metal2 20020 12908 20020 12908 0 segm[2]
rlabel metal2 10108 19677 10108 19677 0 segm[4]
rlabel metal2 9436 19845 9436 19845 0 segm[6]
rlabel metal3 20321 9100 20321 9100 0 segm[7]
rlabel metal2 11452 1099 11452 1099 0 segm[8]
rlabel metal2 20020 11172 20020 11172 0 segm[9]
rlabel metal3 679 12796 679 12796 0 sel[0]
rlabel metal2 10444 1099 10444 1099 0 sel[10]
rlabel metal3 679 9436 679 9436 0 sel[11]
rlabel metal3 679 11116 679 11116 0 sel[1]
rlabel metal3 679 13132 679 13132 0 sel[2]
rlabel metal2 11452 19873 11452 19873 0 sel[3]
rlabel metal2 12796 19957 12796 19957 0 sel[4]
rlabel metal3 679 11788 679 11788 0 sel[5]
rlabel metal2 20020 13356 20020 13356 0 sel[6]
rlabel metal2 19964 13664 19964 13664 0 sel[7]
rlabel metal2 12460 1211 12460 1211 0 sel[8]
rlabel metal2 20020 9548 20020 9548 0 sel[9]
<< properties >>
string FIXED_BBOX 0 0 21000 21000
<< end >>
