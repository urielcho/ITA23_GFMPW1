magic
tech gf180mcuD
magscale 1 5
timestamp 1699645460
<< obsm1 >>
rect 672 1538 20328 19305
<< metal2 >>
rect 8736 20600 8792 21000
rect 9072 20600 9128 21000
rect 9408 20600 9464 21000
rect 11088 20600 11144 21000
rect 11424 20600 11480 21000
rect 12432 20600 12488 21000
rect 13440 20600 13496 21000
rect 8064 0 8120 400
rect 8400 0 8456 400
rect 12432 0 12488 400
<< obsm2 >>
rect 854 20570 8706 20600
rect 8822 20570 9042 20600
rect 9158 20570 9378 20600
rect 9494 20570 11058 20600
rect 11174 20570 11394 20600
rect 11510 20570 12402 20600
rect 12518 20570 13410 20600
rect 13526 20570 20034 20600
rect 854 430 20034 20570
rect 854 400 8034 430
rect 8150 400 8370 430
rect 8486 400 12402 430
rect 12518 400 20034 430
<< metal3 >>
rect 0 18144 400 18200
rect 0 14112 400 14168
rect 0 12768 400 12824
rect 0 12096 400 12152
rect 20600 12096 21000 12152
rect 0 11760 400 11816
rect 20600 11760 21000 11816
rect 0 11424 400 11480
rect 20600 11424 21000 11480
rect 0 11088 400 11144
rect 0 10752 400 10808
rect 20600 10080 21000 10136
rect 0 9072 400 9128
rect 20600 9072 21000 9128
rect 20600 8064 21000 8120
rect 20600 7728 21000 7784
rect 20600 7392 21000 7448
<< obsm3 >>
rect 400 18230 20600 19222
rect 430 18114 20600 18230
rect 400 14198 20600 18114
rect 430 14082 20600 14198
rect 400 12854 20600 14082
rect 430 12738 20600 12854
rect 400 12182 20600 12738
rect 430 12066 20570 12182
rect 400 11846 20600 12066
rect 430 11730 20570 11846
rect 400 11510 20600 11730
rect 430 11394 20570 11510
rect 400 11174 20600 11394
rect 430 11058 20600 11174
rect 400 10838 20600 11058
rect 430 10722 20600 10838
rect 400 10166 20600 10722
rect 400 10050 20570 10166
rect 400 9158 20600 10050
rect 430 9042 20570 9158
rect 400 8150 20600 9042
rect 400 8034 20570 8150
rect 400 7814 20600 8034
rect 400 7698 20570 7814
rect 400 7478 20600 7698
rect 400 7362 20570 7478
rect 400 1554 20600 7362
<< metal4 >>
rect 2224 1538 2384 19238
rect 9904 1538 10064 19238
rect 17584 1538 17744 19238
<< obsm4 >>
rect 11214 11265 11410 11751
<< labels >>
rlabel metal3 s 0 14112 400 14168 6 clk
port 1 nsew signal input
rlabel metal3 s 0 11760 400 11816 6 segm[0]
port 2 nsew signal output
rlabel metal2 s 12432 0 12488 400 6 segm[10]
port 3 nsew signal output
rlabel metal2 s 8736 20600 8792 21000 6 segm[11]
port 4 nsew signal output
rlabel metal2 s 12432 20600 12488 21000 6 segm[12]
port 5 nsew signal output
rlabel metal3 s 20600 11760 21000 11816 6 segm[13]
port 6 nsew signal output
rlabel metal2 s 13440 20600 13496 21000 6 segm[1]
port 7 nsew signal output
rlabel metal3 s 20600 7728 21000 7784 6 segm[2]
port 8 nsew signal output
rlabel metal3 s 0 11088 400 11144 6 segm[3]
port 9 nsew signal output
rlabel metal3 s 0 18144 400 18200 6 segm[4]
port 10 nsew signal output
rlabel metal2 s 9072 20600 9128 21000 6 segm[5]
port 11 nsew signal output
rlabel metal3 s 0 12096 400 12152 6 segm[6]
port 12 nsew signal output
rlabel metal2 s 9408 20600 9464 21000 6 segm[7]
port 13 nsew signal output
rlabel metal3 s 0 10752 400 10808 6 segm[8]
port 14 nsew signal output
rlabel metal2 s 11424 20600 11480 21000 6 segm[9]
port 15 nsew signal output
rlabel metal3 s 20600 12096 21000 12152 6 sel[0]
port 16 nsew signal output
rlabel metal3 s 0 12768 400 12824 6 sel[10]
port 17 nsew signal output
rlabel metal2 s 8400 0 8456 400 6 sel[11]
port 18 nsew signal output
rlabel metal3 s 20600 11424 21000 11480 6 sel[1]
port 19 nsew signal output
rlabel metal3 s 20600 10080 21000 10136 6 sel[2]
port 20 nsew signal output
rlabel metal3 s 20600 9072 21000 9128 6 sel[3]
port 21 nsew signal output
rlabel metal3 s 20600 8064 21000 8120 6 sel[4]
port 22 nsew signal output
rlabel metal2 s 11088 20600 11144 21000 6 sel[5]
port 23 nsew signal output
rlabel metal3 s 20600 7392 21000 7448 6 sel[6]
port 24 nsew signal output
rlabel metal2 s 8064 0 8120 400 6 sel[7]
port 25 nsew signal output
rlabel metal3 s 0 9072 400 9128 6 sel[8]
port 26 nsew signal output
rlabel metal3 s 0 11424 400 11480 6 sel[9]
port 27 nsew signal output
rlabel metal4 s 2224 1538 2384 19238 6 vdd
port 28 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 19238 6 vdd
port 28 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 19238 6 vss
port 29 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 21000 21000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 496442
string GDS_FILE /home/urielcho/Proyectos_caravel/ITA23_GFMPW1b/openlane/ita28/runs/23_11_10_13_42/results/signoff/ita28.magic.gds
string GDS_START 165790
<< end >>

