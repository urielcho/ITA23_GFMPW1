magic
tech gf180mcuD
magscale 1 5
timestamp 1699641638
<< metal1 >>
rect 672 19221 20328 19238
rect 672 19195 2239 19221
rect 2265 19195 2291 19221
rect 2317 19195 2343 19221
rect 2369 19195 17599 19221
rect 17625 19195 17651 19221
rect 17677 19195 17703 19221
rect 17729 19195 20328 19221
rect 672 19178 20328 19195
rect 8975 19137 9001 19143
rect 8975 19105 9001 19111
rect 11047 19137 11073 19143
rect 11047 19105 11073 19111
rect 12783 19137 12809 19143
rect 12783 19105 12809 19111
rect 8465 18999 8471 19025
rect 8497 18999 8503 19025
rect 10537 18999 10543 19025
rect 10569 18999 10575 19025
rect 12273 18999 12279 19025
rect 12305 18999 12311 19025
rect 672 18829 20328 18846
rect 672 18803 9919 18829
rect 9945 18803 9971 18829
rect 9997 18803 10023 18829
rect 10049 18803 20328 18829
rect 672 18786 20328 18803
rect 10039 18745 10065 18751
rect 10039 18713 10065 18719
rect 13735 18745 13761 18751
rect 13735 18713 13761 18719
rect 9585 18607 9591 18633
rect 9617 18607 9623 18633
rect 13225 18607 13231 18633
rect 13257 18607 13263 18633
rect 672 18437 20328 18454
rect 672 18411 2239 18437
rect 2265 18411 2291 18437
rect 2317 18411 2343 18437
rect 2369 18411 17599 18437
rect 17625 18411 17651 18437
rect 17677 18411 17703 18437
rect 17729 18411 20328 18437
rect 672 18394 20328 18411
rect 8359 18353 8385 18359
rect 8359 18321 8385 18327
rect 8073 18215 8079 18241
rect 8105 18215 8111 18241
rect 672 18045 20328 18062
rect 672 18019 9919 18045
rect 9945 18019 9971 18045
rect 9997 18019 10023 18045
rect 10049 18019 20328 18045
rect 672 18002 20328 18019
rect 672 17653 20328 17670
rect 672 17627 2239 17653
rect 2265 17627 2291 17653
rect 2317 17627 2343 17653
rect 2369 17627 17599 17653
rect 17625 17627 17651 17653
rect 17677 17627 17703 17653
rect 17729 17627 20328 17653
rect 672 17610 20328 17627
rect 672 17261 20328 17278
rect 672 17235 9919 17261
rect 9945 17235 9971 17261
rect 9997 17235 10023 17261
rect 10049 17235 20328 17261
rect 672 17218 20328 17235
rect 672 16869 20328 16886
rect 672 16843 2239 16869
rect 2265 16843 2291 16869
rect 2317 16843 2343 16869
rect 2369 16843 17599 16869
rect 17625 16843 17651 16869
rect 17677 16843 17703 16869
rect 17729 16843 20328 16869
rect 672 16826 20328 16843
rect 672 16477 20328 16494
rect 672 16451 9919 16477
rect 9945 16451 9971 16477
rect 9997 16451 10023 16477
rect 10049 16451 20328 16477
rect 672 16434 20328 16451
rect 672 16085 20328 16102
rect 672 16059 2239 16085
rect 2265 16059 2291 16085
rect 2317 16059 2343 16085
rect 2369 16059 17599 16085
rect 17625 16059 17651 16085
rect 17677 16059 17703 16085
rect 17729 16059 20328 16085
rect 672 16042 20328 16059
rect 672 15693 20328 15710
rect 672 15667 9919 15693
rect 9945 15667 9971 15693
rect 9997 15667 10023 15693
rect 10049 15667 20328 15693
rect 672 15650 20328 15667
rect 672 15301 20328 15318
rect 672 15275 2239 15301
rect 2265 15275 2291 15301
rect 2317 15275 2343 15301
rect 2369 15275 17599 15301
rect 17625 15275 17651 15301
rect 17677 15275 17703 15301
rect 17729 15275 20328 15301
rect 672 15258 20328 15275
rect 672 14909 20328 14926
rect 672 14883 9919 14909
rect 9945 14883 9971 14909
rect 9997 14883 10023 14909
rect 10049 14883 20328 14909
rect 672 14866 20328 14883
rect 672 14517 20328 14534
rect 672 14491 2239 14517
rect 2265 14491 2291 14517
rect 2317 14491 2343 14517
rect 2369 14491 17599 14517
rect 17625 14491 17651 14517
rect 17677 14491 17703 14517
rect 17729 14491 20328 14517
rect 672 14474 20328 14491
rect 8247 14209 8273 14215
rect 8247 14177 8273 14183
rect 672 14125 20328 14142
rect 672 14099 9919 14125
rect 9945 14099 9971 14125
rect 9997 14099 10023 14125
rect 10049 14099 20328 14125
rect 672 14082 20328 14099
rect 8247 14041 8273 14047
rect 8409 14015 8415 14041
rect 8441 14015 8447 14041
rect 8247 14009 8273 14015
rect 12671 13985 12697 13991
rect 12671 13953 12697 13959
rect 12615 13929 12641 13935
rect 6673 13903 6679 13929
rect 6705 13903 6711 13929
rect 8969 13903 8975 13929
rect 9001 13903 9007 13929
rect 18825 13903 18831 13929
rect 18857 13903 18863 13929
rect 12615 13897 12641 13903
rect 10655 13873 10681 13879
rect 7009 13847 7015 13873
rect 7041 13847 7047 13873
rect 8073 13847 8079 13873
rect 8105 13847 8111 13873
rect 9361 13847 9367 13873
rect 9393 13847 9399 13873
rect 10425 13847 10431 13873
rect 10457 13847 10463 13873
rect 10655 13841 10681 13847
rect 13735 13873 13761 13879
rect 13735 13841 13761 13847
rect 12671 13817 12697 13823
rect 12671 13785 12697 13791
rect 13679 13817 13705 13823
rect 13679 13785 13705 13791
rect 20007 13817 20033 13823
rect 20007 13785 20033 13791
rect 672 13733 20328 13750
rect 672 13707 2239 13733
rect 2265 13707 2291 13733
rect 2317 13707 2343 13733
rect 2369 13707 17599 13733
rect 17625 13707 17651 13733
rect 17677 13707 17703 13733
rect 17729 13707 20328 13733
rect 672 13690 20328 13707
rect 7407 13649 7433 13655
rect 7407 13617 7433 13623
rect 7575 13593 7601 13599
rect 10263 13593 10289 13599
rect 7793 13567 7799 13593
rect 7825 13567 7831 13593
rect 9585 13567 9591 13593
rect 9617 13567 9623 13593
rect 12049 13567 12055 13593
rect 12081 13567 12087 13593
rect 13113 13567 13119 13593
rect 13145 13567 13151 13593
rect 7575 13561 7601 13567
rect 10263 13561 10289 13567
rect 9871 13537 9897 13543
rect 8129 13511 8135 13537
rect 8161 13511 8167 13537
rect 9871 13505 9897 13511
rect 11215 13537 11241 13543
rect 11713 13511 11719 13537
rect 11745 13511 11751 13537
rect 11215 13505 11241 13511
rect 7463 13481 7489 13487
rect 7463 13449 7489 13455
rect 7855 13481 7881 13487
rect 7855 13449 7881 13455
rect 7967 13481 7993 13487
rect 9759 13481 9785 13487
rect 8521 13455 8527 13481
rect 8553 13455 8559 13481
rect 7967 13449 7993 13455
rect 9759 13449 9785 13455
rect 11495 13481 11521 13487
rect 11495 13449 11521 13455
rect 9815 13425 9841 13431
rect 9815 13393 9841 13399
rect 9983 13425 10009 13431
rect 9983 13393 10009 13399
rect 11383 13425 11409 13431
rect 11383 13393 11409 13399
rect 11551 13425 11577 13431
rect 11551 13393 11577 13399
rect 13343 13425 13369 13431
rect 13343 13393 13369 13399
rect 672 13341 20328 13358
rect 672 13315 9919 13341
rect 9945 13315 9971 13341
rect 9997 13315 10023 13341
rect 10049 13315 20328 13341
rect 672 13298 20328 13315
rect 8975 13257 9001 13263
rect 8975 13225 9001 13231
rect 9479 13257 9505 13263
rect 9479 13225 9505 13231
rect 9703 13201 9729 13207
rect 9703 13169 9729 13175
rect 10375 13201 10401 13207
rect 10375 13169 10401 13175
rect 8863 13145 8889 13151
rect 7569 13119 7575 13145
rect 7601 13119 7607 13145
rect 8863 13113 8889 13119
rect 9031 13145 9057 13151
rect 9031 13113 9057 13119
rect 9143 13145 9169 13151
rect 9143 13113 9169 13119
rect 9367 13145 9393 13151
rect 9367 13113 9393 13119
rect 9535 13145 9561 13151
rect 9535 13113 9561 13119
rect 9815 13145 9841 13151
rect 9815 13113 9841 13119
rect 9983 13145 10009 13151
rect 9983 13113 10009 13119
rect 10263 13145 10289 13151
rect 10263 13113 10289 13119
rect 10431 13145 10457 13151
rect 10817 13119 10823 13145
rect 10849 13119 10855 13145
rect 12777 13119 12783 13145
rect 12809 13119 12815 13145
rect 10431 13113 10457 13119
rect 14463 13089 14489 13095
rect 11153 13063 11159 13089
rect 11185 13063 11191 13089
rect 12217 13063 12223 13089
rect 12249 13063 12255 13089
rect 13169 13063 13175 13089
rect 13201 13063 13207 13089
rect 14233 13063 14239 13089
rect 14265 13063 14271 13089
rect 14463 13057 14489 13063
rect 7575 13033 7601 13039
rect 7575 13001 7601 13007
rect 7743 13033 7769 13039
rect 7743 13001 7769 13007
rect 9759 13033 9785 13039
rect 9759 13001 9785 13007
rect 10095 13033 10121 13039
rect 10095 13001 10121 13007
rect 672 12949 20328 12966
rect 672 12923 2239 12949
rect 2265 12923 2291 12949
rect 2317 12923 2343 12949
rect 2369 12923 17599 12949
rect 17625 12923 17651 12949
rect 17677 12923 17703 12949
rect 17729 12923 20328 12949
rect 672 12906 20328 12923
rect 967 12809 993 12815
rect 12223 12809 12249 12815
rect 20007 12809 20033 12815
rect 6729 12783 6735 12809
rect 6761 12783 6767 12809
rect 12553 12783 12559 12809
rect 12585 12783 12591 12809
rect 13113 12783 13119 12809
rect 13145 12783 13151 12809
rect 967 12777 993 12783
rect 12223 12777 12249 12783
rect 20007 12777 20033 12783
rect 8359 12753 8385 12759
rect 2137 12727 2143 12753
rect 2169 12727 2175 12753
rect 8129 12727 8135 12753
rect 8161 12727 8167 12753
rect 8359 12721 8385 12727
rect 11327 12753 11353 12759
rect 11327 12721 11353 12727
rect 11495 12753 11521 12759
rect 13063 12753 13089 12759
rect 12497 12727 12503 12753
rect 12529 12727 12535 12753
rect 18825 12727 18831 12753
rect 18857 12727 18863 12753
rect 11495 12721 11521 12727
rect 13063 12721 13089 12727
rect 12391 12697 12417 12703
rect 7793 12671 7799 12697
rect 7825 12671 7831 12697
rect 8521 12671 8527 12697
rect 8553 12671 8559 12697
rect 12391 12665 12417 12671
rect 12615 12697 12641 12703
rect 12615 12665 12641 12671
rect 12839 12697 12865 12703
rect 12839 12665 12865 12671
rect 13119 12697 13145 12703
rect 13119 12665 13145 12671
rect 13791 12697 13817 12703
rect 13791 12665 13817 12671
rect 13847 12697 13873 12703
rect 13847 12665 13873 12671
rect 8751 12641 8777 12647
rect 8751 12609 8777 12615
rect 11439 12641 11465 12647
rect 11439 12609 11465 12615
rect 12951 12641 12977 12647
rect 12951 12609 12977 12615
rect 13959 12641 13985 12647
rect 13959 12609 13985 12615
rect 672 12557 20328 12574
rect 672 12531 9919 12557
rect 9945 12531 9971 12557
rect 9997 12531 10023 12557
rect 10049 12531 20328 12557
rect 672 12514 20328 12531
rect 7295 12473 7321 12479
rect 12105 12447 12111 12473
rect 12137 12447 12143 12473
rect 7295 12441 7321 12447
rect 7239 12361 7265 12367
rect 2137 12335 2143 12361
rect 2169 12335 2175 12361
rect 7239 12329 7265 12335
rect 7351 12361 7377 12367
rect 7351 12329 7377 12335
rect 7575 12361 7601 12367
rect 9529 12335 9535 12361
rect 9561 12335 9567 12361
rect 12217 12335 12223 12361
rect 12249 12335 12255 12361
rect 13617 12335 13623 12361
rect 13649 12335 13655 12361
rect 7575 12329 7601 12335
rect 7463 12305 7489 12311
rect 11159 12305 11185 12311
rect 15247 12305 15273 12311
rect 9865 12279 9871 12305
rect 9897 12279 9903 12305
rect 10929 12279 10935 12305
rect 10961 12279 10967 12305
rect 13953 12279 13959 12305
rect 13985 12279 13991 12305
rect 15017 12279 15023 12305
rect 15049 12279 15055 12305
rect 7463 12273 7489 12279
rect 11159 12273 11185 12279
rect 15247 12273 15273 12279
rect 967 12249 993 12255
rect 967 12217 993 12223
rect 672 12165 20328 12182
rect 672 12139 2239 12165
rect 2265 12139 2291 12165
rect 2317 12139 2343 12165
rect 2369 12139 17599 12165
rect 17625 12139 17651 12165
rect 17677 12139 17703 12165
rect 17729 12139 20328 12165
rect 672 12122 20328 12139
rect 967 12025 993 12031
rect 967 11993 993 11999
rect 9647 12025 9673 12031
rect 9647 11993 9673 11999
rect 20007 12025 20033 12031
rect 20007 11993 20033 11999
rect 8863 11969 8889 11975
rect 2025 11943 2031 11969
rect 2057 11943 2063 11969
rect 7009 11943 7015 11969
rect 7041 11943 7047 11969
rect 8863 11937 8889 11943
rect 9591 11969 9617 11975
rect 9591 11937 9617 11943
rect 9815 11969 9841 11975
rect 14071 11969 14097 11975
rect 9865 11943 9871 11969
rect 9897 11943 9903 11969
rect 18825 11943 18831 11969
rect 18857 11943 18863 11969
rect 9815 11937 9841 11943
rect 14071 11937 14097 11943
rect 8695 11913 8721 11919
rect 6897 11887 6903 11913
rect 6929 11887 6935 11913
rect 8695 11881 8721 11887
rect 8975 11913 9001 11919
rect 11215 11913 11241 11919
rect 13791 11913 13817 11919
rect 9697 11887 9703 11913
rect 9729 11887 9735 11913
rect 10649 11887 10655 11913
rect 10681 11887 10687 11913
rect 12497 11887 12503 11913
rect 12529 11887 12535 11913
rect 8975 11881 9001 11887
rect 11215 11881 11241 11887
rect 13791 11881 13817 11887
rect 13903 11913 13929 11919
rect 13903 11881 13929 11887
rect 7295 11857 7321 11863
rect 7295 11825 7321 11831
rect 8751 11857 8777 11863
rect 8751 11825 8777 11831
rect 10823 11857 10849 11863
rect 10823 11825 10849 11831
rect 11383 11857 11409 11863
rect 11383 11825 11409 11831
rect 11551 11857 11577 11863
rect 12671 11857 12697 11863
rect 11713 11831 11719 11857
rect 11745 11831 11751 11857
rect 11551 11825 11577 11831
rect 12671 11825 12697 11831
rect 13959 11857 13985 11863
rect 13959 11825 13985 11831
rect 672 11773 20328 11790
rect 672 11747 9919 11773
rect 9945 11747 9971 11773
rect 9997 11747 10023 11773
rect 10049 11747 20328 11773
rect 672 11730 20328 11747
rect 9031 11689 9057 11695
rect 9031 11657 9057 11663
rect 9255 11689 9281 11695
rect 9255 11657 9281 11663
rect 10095 11689 10121 11695
rect 10095 11657 10121 11663
rect 10655 11689 10681 11695
rect 10655 11657 10681 11663
rect 7127 11633 7153 11639
rect 7127 11601 7153 11607
rect 7239 11633 7265 11639
rect 7239 11601 7265 11607
rect 7351 11633 7377 11639
rect 7351 11601 7377 11607
rect 7687 11633 7713 11639
rect 7687 11601 7713 11607
rect 9871 11633 9897 11639
rect 10481 11607 10487 11633
rect 10513 11607 10519 11633
rect 11657 11607 11663 11633
rect 11689 11607 11695 11633
rect 9871 11601 9897 11607
rect 7463 11577 7489 11583
rect 2137 11551 2143 11577
rect 2169 11551 2175 11577
rect 6897 11551 6903 11577
rect 6929 11551 6935 11577
rect 7463 11545 7489 11551
rect 9143 11577 9169 11583
rect 9143 11545 9169 11551
rect 10263 11577 10289 11583
rect 10263 11545 10289 11551
rect 11495 11577 11521 11583
rect 13393 11551 13399 11577
rect 13425 11551 13431 11577
rect 11495 11545 11521 11551
rect 7631 11521 7657 11527
rect 5497 11495 5503 11521
rect 5529 11495 5535 11521
rect 6561 11495 6567 11521
rect 6593 11495 6599 11521
rect 7631 11489 7657 11495
rect 9087 11521 9113 11527
rect 9087 11489 9113 11495
rect 9535 11521 9561 11527
rect 9535 11489 9561 11495
rect 10823 11521 10849 11527
rect 15023 11521 15049 11527
rect 13729 11495 13735 11521
rect 13761 11495 13767 11521
rect 14793 11495 14799 11521
rect 14825 11495 14831 11521
rect 10823 11489 10849 11495
rect 15023 11489 15049 11495
rect 967 11465 993 11471
rect 967 11433 993 11439
rect 7575 11465 7601 11471
rect 7575 11433 7601 11439
rect 9759 11465 9785 11471
rect 9759 11433 9785 11439
rect 9927 11465 9953 11471
rect 9927 11433 9953 11439
rect 10879 11465 10905 11471
rect 10879 11433 10905 11439
rect 672 11381 20328 11398
rect 672 11355 2239 11381
rect 2265 11355 2291 11381
rect 2317 11355 2343 11381
rect 2369 11355 17599 11381
rect 17625 11355 17651 11381
rect 17677 11355 17703 11381
rect 17729 11355 20328 11381
rect 672 11338 20328 11355
rect 9311 11297 9337 11303
rect 7121 11271 7127 11297
rect 7153 11271 7159 11297
rect 9311 11265 9337 11271
rect 13903 11241 13929 11247
rect 7681 11215 7687 11241
rect 7713 11215 7719 11241
rect 8745 11215 8751 11241
rect 8777 11215 8783 11241
rect 10817 11215 10823 11241
rect 10849 11215 10855 11241
rect 12665 11215 12671 11241
rect 12697 11215 12703 11241
rect 13903 11209 13929 11215
rect 20007 11241 20033 11247
rect 20007 11209 20033 11215
rect 6791 11185 6817 11191
rect 9479 11185 9505 11191
rect 9137 11159 9143 11185
rect 9169 11159 9175 11185
rect 6791 11153 6817 11159
rect 9479 11153 9505 11159
rect 10375 11185 10401 11191
rect 13175 11185 13201 11191
rect 13511 11185 13537 11191
rect 10761 11159 10767 11185
rect 10793 11159 10799 11185
rect 11265 11159 11271 11185
rect 11297 11159 11303 11185
rect 13393 11159 13399 11185
rect 13425 11159 13431 11185
rect 10375 11153 10401 11159
rect 13175 11153 13201 11159
rect 13511 11153 13537 11159
rect 13623 11185 13649 11191
rect 18825 11159 18831 11185
rect 18857 11159 18863 11185
rect 13623 11153 13649 11159
rect 6847 11129 6873 11135
rect 6847 11097 6873 11103
rect 6903 11129 6929 11135
rect 6903 11097 6929 11103
rect 9591 11129 9617 11135
rect 11047 11129 11073 11135
rect 12839 11129 12865 11135
rect 9977 11103 9983 11129
rect 10009 11103 10015 11129
rect 10201 11103 10207 11129
rect 10233 11103 10239 11129
rect 11601 11103 11607 11129
rect 11633 11103 11639 11129
rect 9591 11097 9617 11103
rect 11047 11097 11073 11103
rect 12839 11097 12865 11103
rect 12895 11129 12921 11135
rect 12895 11097 12921 11103
rect 13007 11129 13033 11135
rect 13007 11097 13033 11103
rect 13847 11129 13873 11135
rect 13847 11097 13873 11103
rect 13959 11129 13985 11135
rect 13959 11097 13985 11103
rect 13455 11073 13481 11079
rect 10145 11047 10151 11073
rect 10177 11047 10183 11073
rect 13455 11041 13481 11047
rect 672 10989 20328 11006
rect 672 10963 9919 10989
rect 9945 10963 9971 10989
rect 9997 10963 10023 10989
rect 10049 10963 20328 10989
rect 672 10946 20328 10963
rect 11551 10905 11577 10911
rect 11551 10873 11577 10879
rect 11495 10849 11521 10855
rect 11495 10817 11521 10823
rect 12615 10849 12641 10855
rect 13119 10849 13145 10855
rect 12945 10823 12951 10849
rect 12977 10823 12983 10849
rect 12615 10817 12641 10823
rect 13119 10817 13145 10823
rect 13343 10849 13369 10855
rect 13343 10817 13369 10823
rect 13791 10793 13817 10799
rect 2137 10767 2143 10793
rect 2169 10767 2175 10793
rect 11321 10767 11327 10793
rect 11353 10767 11359 10793
rect 11657 10767 11663 10793
rect 11689 10767 11695 10793
rect 12721 10767 12727 10793
rect 12753 10767 12759 10793
rect 14009 10767 14015 10793
rect 14041 10767 14047 10793
rect 13791 10761 13817 10767
rect 13287 10737 13313 10743
rect 9473 10711 9479 10737
rect 9505 10711 9511 10737
rect 13287 10705 13313 10711
rect 13847 10737 13873 10743
rect 15695 10737 15721 10743
rect 14401 10711 14407 10737
rect 14433 10711 14439 10737
rect 15465 10711 15471 10737
rect 15497 10711 15503 10737
rect 13847 10705 13873 10711
rect 15695 10705 15721 10711
rect 967 10681 993 10687
rect 967 10649 993 10655
rect 13623 10681 13649 10687
rect 13623 10649 13649 10655
rect 13679 10681 13705 10687
rect 13679 10649 13705 10655
rect 672 10597 20328 10614
rect 672 10571 2239 10597
rect 2265 10571 2291 10597
rect 2317 10571 2343 10597
rect 2369 10571 17599 10597
rect 17625 10571 17651 10597
rect 17677 10571 17703 10597
rect 17729 10571 20328 10597
rect 672 10554 20328 10571
rect 8471 10513 8497 10519
rect 8863 10513 8889 10519
rect 8689 10487 8695 10513
rect 8721 10487 8727 10513
rect 9865 10487 9871 10513
rect 9897 10487 9903 10513
rect 8471 10481 8497 10487
rect 8863 10481 8889 10487
rect 8975 10457 9001 10463
rect 14127 10457 14153 10463
rect 4993 10431 4999 10457
rect 5025 10431 5031 10457
rect 9249 10431 9255 10457
rect 9281 10431 9287 10457
rect 8975 10425 9001 10431
rect 14127 10425 14153 10431
rect 20007 10457 20033 10463
rect 20007 10425 20033 10431
rect 6735 10401 6761 10407
rect 10431 10401 10457 10407
rect 14071 10401 14097 10407
rect 6393 10375 6399 10401
rect 6425 10375 6431 10401
rect 9305 10375 9311 10401
rect 9337 10375 9343 10401
rect 9585 10375 9591 10401
rect 9617 10375 9623 10401
rect 9697 10375 9703 10401
rect 9729 10375 9735 10401
rect 9809 10375 9815 10401
rect 9841 10375 9847 10401
rect 10649 10375 10655 10401
rect 10681 10375 10687 10401
rect 13561 10375 13567 10401
rect 13593 10375 13599 10401
rect 14233 10375 14239 10401
rect 14265 10375 14271 10401
rect 18825 10375 18831 10401
rect 18857 10375 18863 10401
rect 6735 10369 6761 10375
rect 10431 10369 10457 10375
rect 14071 10369 14097 10375
rect 6847 10345 6873 10351
rect 6057 10319 6063 10345
rect 6089 10319 6095 10345
rect 6847 10313 6873 10319
rect 6903 10345 6929 10351
rect 8415 10345 8441 10351
rect 6953 10319 6959 10345
rect 6985 10319 6991 10345
rect 6903 10313 6929 10319
rect 8415 10313 8441 10319
rect 8471 10345 8497 10351
rect 12553 10319 12559 10345
rect 12585 10319 12591 10345
rect 8471 10313 8497 10319
rect 6791 10289 6817 10295
rect 13449 10263 13455 10289
rect 13481 10263 13487 10289
rect 6791 10257 6817 10263
rect 672 10205 20328 10222
rect 672 10179 9919 10205
rect 9945 10179 9971 10205
rect 9997 10179 10023 10205
rect 10049 10179 20328 10205
rect 672 10162 20328 10179
rect 10879 10121 10905 10127
rect 9249 10095 9255 10121
rect 9281 10095 9287 10121
rect 10879 10089 10905 10095
rect 6119 10065 6145 10071
rect 6119 10033 6145 10039
rect 6231 10065 6257 10071
rect 6231 10033 6257 10039
rect 8863 10065 8889 10071
rect 8863 10033 8889 10039
rect 10207 10065 10233 10071
rect 12279 10065 12305 10071
rect 11041 10039 11047 10065
rect 11073 10039 11079 10065
rect 10207 10033 10233 10039
rect 12279 10033 12305 10039
rect 8919 10009 8945 10015
rect 2137 9983 2143 10009
rect 2169 9983 2175 10009
rect 6785 9983 6791 10009
rect 6817 9983 6823 10009
rect 8919 9977 8945 9983
rect 9087 10009 9113 10015
rect 9087 9977 9113 9983
rect 9703 10009 9729 10015
rect 11215 10009 11241 10015
rect 10649 9983 10655 10009
rect 10681 9983 10687 10009
rect 10761 9983 10767 10009
rect 10793 9983 10799 10009
rect 9703 9977 9729 9983
rect 11215 9977 11241 9983
rect 12223 10009 12249 10015
rect 12609 9983 12615 10009
rect 12641 9983 12647 10009
rect 12223 9977 12249 9983
rect 6567 9953 6593 9959
rect 9423 9953 9449 9959
rect 6057 9927 6063 9953
rect 6089 9927 6095 9953
rect 7177 9927 7183 9953
rect 7209 9927 7215 9953
rect 8241 9927 8247 9953
rect 8273 9927 8279 9953
rect 6567 9921 6593 9927
rect 9423 9921 9449 9927
rect 9927 9953 9953 9959
rect 10817 9927 10823 9953
rect 10849 9927 10855 9953
rect 14457 9927 14463 9953
rect 14489 9927 14495 9953
rect 9927 9921 9953 9927
rect 967 9897 993 9903
rect 967 9865 993 9871
rect 12279 9897 12305 9903
rect 12279 9865 12305 9871
rect 672 9813 20328 9830
rect 672 9787 2239 9813
rect 2265 9787 2291 9813
rect 2317 9787 2343 9813
rect 2369 9787 17599 9813
rect 17625 9787 17651 9813
rect 17677 9787 17703 9813
rect 17729 9787 20328 9813
rect 672 9770 20328 9787
rect 10655 9729 10681 9735
rect 10655 9697 10681 9703
rect 10823 9729 10849 9735
rect 10823 9697 10849 9703
rect 13175 9729 13201 9735
rect 13175 9697 13201 9703
rect 14127 9729 14153 9735
rect 14127 9697 14153 9703
rect 12615 9673 12641 9679
rect 4937 9647 4943 9673
rect 4969 9647 4975 9673
rect 9753 9647 9759 9673
rect 9785 9647 9791 9673
rect 12615 9641 12641 9647
rect 13063 9673 13089 9679
rect 13063 9641 13089 9647
rect 8919 9617 8945 9623
rect 12727 9617 12753 9623
rect 6393 9591 6399 9617
rect 6425 9591 6431 9617
rect 6729 9591 6735 9617
rect 6761 9591 6767 9617
rect 9361 9591 9367 9617
rect 9393 9591 9399 9617
rect 9641 9591 9647 9617
rect 9673 9591 9679 9617
rect 10201 9591 10207 9617
rect 10233 9591 10239 9617
rect 10649 9591 10655 9617
rect 10681 9591 10687 9617
rect 12105 9591 12111 9617
rect 12137 9591 12143 9617
rect 8919 9585 8945 9591
rect 12727 9585 12753 9591
rect 13511 9617 13537 9623
rect 13511 9585 13537 9591
rect 13847 9617 13873 9623
rect 14239 9617 14265 9623
rect 14009 9591 14015 9617
rect 14041 9591 14047 9617
rect 13847 9585 13873 9591
rect 14239 9585 14265 9591
rect 6903 9561 6929 9567
rect 10991 9561 11017 9567
rect 14295 9561 14321 9567
rect 6001 9535 6007 9561
rect 6033 9535 6039 9561
rect 9137 9535 9143 9561
rect 9169 9535 9175 9561
rect 9697 9535 9703 9561
rect 9729 9535 9735 9561
rect 11153 9535 11159 9561
rect 11185 9535 11191 9561
rect 11769 9535 11775 9561
rect 11801 9535 11807 9561
rect 12049 9535 12055 9561
rect 12081 9535 12087 9561
rect 6903 9529 6929 9535
rect 10991 9529 11017 9535
rect 14295 9529 14321 9535
rect 14575 9561 14601 9567
rect 14575 9529 14601 9535
rect 6847 9505 6873 9511
rect 6847 9473 6873 9479
rect 8359 9505 8385 9511
rect 8359 9473 8385 9479
rect 8751 9505 8777 9511
rect 8751 9473 8777 9479
rect 8863 9505 8889 9511
rect 13735 9505 13761 9511
rect 9361 9479 9367 9505
rect 9393 9479 9399 9505
rect 11713 9479 11719 9505
rect 11745 9479 11751 9505
rect 12889 9479 12895 9505
rect 12921 9479 12927 9505
rect 13337 9479 13343 9505
rect 13369 9479 13375 9505
rect 8863 9473 8889 9479
rect 13735 9473 13761 9479
rect 13791 9505 13817 9511
rect 13791 9473 13817 9479
rect 14631 9505 14657 9511
rect 14631 9473 14657 9479
rect 14687 9505 14713 9511
rect 14687 9473 14713 9479
rect 672 9421 20328 9438
rect 672 9395 9919 9421
rect 9945 9395 9971 9421
rect 9997 9395 10023 9421
rect 10049 9395 20328 9421
rect 672 9378 20328 9395
rect 9703 9337 9729 9343
rect 9703 9305 9729 9311
rect 6175 9281 6201 9287
rect 8303 9281 8329 9287
rect 11439 9281 11465 9287
rect 7793 9255 7799 9281
rect 7825 9255 7831 9281
rect 9865 9255 9871 9281
rect 9897 9255 9903 9281
rect 10313 9255 10319 9281
rect 10345 9255 10351 9281
rect 6175 9249 6201 9255
rect 8303 9249 8329 9255
rect 11439 9249 11465 9255
rect 11551 9281 11577 9287
rect 13567 9281 13593 9287
rect 11769 9255 11775 9281
rect 11801 9255 11807 9281
rect 12049 9255 12055 9281
rect 12081 9255 12087 9281
rect 13001 9255 13007 9281
rect 13033 9255 13039 9281
rect 14401 9255 14407 9281
rect 14433 9255 14439 9281
rect 11551 9249 11577 9255
rect 13567 9249 13593 9255
rect 6231 9225 6257 9231
rect 6231 9193 6257 9199
rect 6343 9225 6369 9231
rect 7407 9225 7433 9231
rect 8639 9225 8665 9231
rect 6449 9199 6455 9225
rect 6481 9199 6487 9225
rect 7737 9199 7743 9225
rect 7769 9199 7775 9225
rect 6343 9193 6369 9199
rect 7407 9193 7433 9199
rect 8639 9193 8665 9199
rect 8807 9225 8833 9231
rect 9535 9225 9561 9231
rect 9025 9199 9031 9225
rect 9057 9199 9063 9225
rect 8807 9193 8833 9199
rect 9535 9193 9561 9199
rect 10151 9225 10177 9231
rect 11383 9225 11409 9231
rect 11153 9199 11159 9225
rect 11185 9199 11191 9225
rect 12105 9199 12111 9225
rect 12137 9199 12143 9225
rect 12945 9199 12951 9225
rect 12977 9199 12983 9225
rect 13505 9199 13511 9225
rect 13537 9199 13543 9225
rect 14009 9199 14015 9225
rect 14041 9199 14047 9225
rect 10151 9193 10177 9199
rect 11383 9193 11409 9199
rect 6679 9169 6705 9175
rect 9479 9169 9505 9175
rect 15695 9169 15721 9175
rect 8913 9143 8919 9169
rect 8945 9143 8951 9169
rect 13057 9143 13063 9169
rect 13089 9143 13095 9169
rect 15465 9143 15471 9169
rect 15497 9143 15503 9169
rect 6679 9137 6705 9143
rect 9479 9137 9505 9143
rect 15695 9137 15721 9143
rect 7239 9113 7265 9119
rect 7239 9081 7265 9087
rect 8247 9113 8273 9119
rect 8247 9081 8273 9087
rect 8415 9113 8441 9119
rect 8415 9081 8441 9087
rect 11271 9113 11297 9119
rect 11271 9081 11297 9087
rect 672 9029 20328 9046
rect 672 9003 2239 9029
rect 2265 9003 2291 9029
rect 2317 9003 2343 9029
rect 2369 9003 17599 9029
rect 17625 9003 17651 9029
rect 17677 9003 17703 9029
rect 17729 9003 20328 9029
rect 672 8986 20328 9003
rect 6287 8945 6313 8951
rect 6287 8913 6313 8919
rect 7855 8945 7881 8951
rect 7855 8913 7881 8919
rect 8023 8945 8049 8951
rect 8023 8913 8049 8919
rect 13623 8945 13649 8951
rect 13623 8913 13649 8919
rect 967 8889 993 8895
rect 14183 8889 14209 8895
rect 6449 8863 6455 8889
rect 6481 8863 6487 8889
rect 6953 8863 6959 8889
rect 6985 8863 6991 8889
rect 8409 8863 8415 8889
rect 8441 8863 8447 8889
rect 967 8857 993 8863
rect 14183 8857 14209 8863
rect 14799 8889 14825 8895
rect 14799 8857 14825 8863
rect 20007 8889 20033 8895
rect 20007 8857 20033 8863
rect 7127 8833 7153 8839
rect 2137 8807 2143 8833
rect 2169 8807 2175 8833
rect 7127 8801 7153 8807
rect 7463 8833 7489 8839
rect 9423 8833 9449 8839
rect 8241 8807 8247 8833
rect 8273 8807 8279 8833
rect 8745 8807 8751 8833
rect 8777 8807 8783 8833
rect 8913 8807 8919 8833
rect 8945 8807 8951 8833
rect 7463 8801 7489 8807
rect 9423 8801 9449 8807
rect 10375 8833 10401 8839
rect 11607 8833 11633 8839
rect 13119 8833 13145 8839
rect 10705 8807 10711 8833
rect 10737 8807 10743 8833
rect 12161 8807 12167 8833
rect 12193 8807 12199 8833
rect 13001 8807 13007 8833
rect 13033 8807 13039 8833
rect 10375 8801 10401 8807
rect 11607 8801 11633 8807
rect 13119 8801 13145 8807
rect 13175 8833 13201 8839
rect 13567 8833 13593 8839
rect 14015 8833 14041 8839
rect 14239 8833 14265 8839
rect 13393 8807 13399 8833
rect 13425 8807 13431 8833
rect 13841 8807 13847 8833
rect 13873 8807 13879 8833
rect 14121 8807 14127 8833
rect 14153 8807 14159 8833
rect 13175 8801 13201 8807
rect 13567 8801 13593 8807
rect 14015 8801 14041 8807
rect 14239 8801 14265 8807
rect 14575 8833 14601 8839
rect 14575 8801 14601 8807
rect 14967 8833 14993 8839
rect 14967 8801 14993 8807
rect 15135 8833 15161 8839
rect 15135 8801 15161 8807
rect 15303 8833 15329 8839
rect 18825 8807 18831 8833
rect 18857 8807 18863 8833
rect 15303 8801 15329 8807
rect 6399 8777 6425 8783
rect 6399 8745 6425 8751
rect 7015 8777 7041 8783
rect 7015 8745 7041 8751
rect 7239 8777 7265 8783
rect 11271 8777 11297 8783
rect 9193 8751 9199 8777
rect 9225 8751 9231 8777
rect 10761 8751 10767 8777
rect 10793 8751 10799 8777
rect 10929 8751 10935 8777
rect 10961 8751 10967 8777
rect 7239 8745 7265 8751
rect 11271 8745 11297 8751
rect 11943 8777 11969 8783
rect 11943 8745 11969 8751
rect 13623 8777 13649 8783
rect 13623 8745 13649 8751
rect 14687 8777 14713 8783
rect 14687 8745 14713 8751
rect 14855 8777 14881 8783
rect 14855 8745 14881 8751
rect 6959 8721 6985 8727
rect 6959 8689 6985 8695
rect 7407 8721 7433 8727
rect 7407 8689 7433 8695
rect 7911 8721 7937 8727
rect 11775 8721 11801 8727
rect 8689 8695 8695 8721
rect 8721 8695 8727 8721
rect 9585 8695 9591 8721
rect 9617 8695 9623 8721
rect 10201 8695 10207 8721
rect 10233 8695 10239 8721
rect 11433 8695 11439 8721
rect 11465 8695 11471 8721
rect 7911 8689 7937 8695
rect 11775 8689 11801 8695
rect 11831 8721 11857 8727
rect 11831 8689 11857 8695
rect 11887 8721 11913 8727
rect 11887 8689 11913 8695
rect 15079 8721 15105 8727
rect 15079 8689 15105 8695
rect 672 8637 20328 8654
rect 672 8611 9919 8637
rect 9945 8611 9971 8637
rect 9997 8611 10023 8637
rect 10049 8611 20328 8637
rect 672 8594 20328 8611
rect 11215 8553 11241 8559
rect 11215 8521 11241 8527
rect 15527 8553 15553 8559
rect 15527 8521 15553 8527
rect 7463 8497 7489 8503
rect 6617 8471 6623 8497
rect 6649 8471 6655 8497
rect 7463 8465 7489 8471
rect 11159 8497 11185 8503
rect 14233 8471 14239 8497
rect 14265 8471 14271 8497
rect 11159 8465 11185 8471
rect 7239 8441 7265 8447
rect 7009 8415 7015 8441
rect 7041 8415 7047 8441
rect 7239 8409 7265 8415
rect 7631 8441 7657 8447
rect 7631 8409 7657 8415
rect 7799 8441 7825 8447
rect 8135 8441 8161 8447
rect 7905 8415 7911 8441
rect 7937 8415 7943 8441
rect 7799 8409 7825 8415
rect 8135 8409 8161 8415
rect 8303 8441 8329 8447
rect 8303 8409 8329 8415
rect 8919 8441 8945 8447
rect 8919 8409 8945 8415
rect 9199 8441 9225 8447
rect 9199 8409 9225 8415
rect 11327 8441 11353 8447
rect 13897 8415 13903 8441
rect 13929 8415 13935 8441
rect 18825 8415 18831 8441
rect 18857 8415 18863 8441
rect 11327 8409 11353 8415
rect 7687 8385 7713 8391
rect 5553 8359 5559 8385
rect 5585 8359 5591 8385
rect 7687 8353 7713 8359
rect 8247 8385 8273 8391
rect 20007 8385 20033 8391
rect 15297 8359 15303 8385
rect 15329 8359 15335 8385
rect 8247 8353 8273 8359
rect 20007 8353 20033 8359
rect 8023 8329 8049 8335
rect 8023 8297 8049 8303
rect 672 8245 20328 8262
rect 672 8219 2239 8245
rect 2265 8219 2291 8245
rect 2317 8219 2343 8245
rect 2369 8219 17599 8245
rect 17625 8219 17651 8245
rect 17677 8219 17703 8245
rect 17729 8219 20328 8245
rect 672 8202 20328 8219
rect 10935 8161 10961 8167
rect 10935 8129 10961 8135
rect 7519 8049 7545 8055
rect 8639 8049 8665 8055
rect 8353 8023 8359 8049
rect 8385 8023 8391 8049
rect 7519 8017 7545 8023
rect 8639 8017 8665 8023
rect 10095 8049 10121 8055
rect 10711 8049 10737 8055
rect 10257 8023 10263 8049
rect 10289 8023 10295 8049
rect 10095 8017 10121 8023
rect 10711 8017 10737 8023
rect 11047 8049 11073 8055
rect 11047 8017 11073 8023
rect 11663 8049 11689 8055
rect 11663 8017 11689 8023
rect 8695 7993 8721 7999
rect 8695 7961 8721 7967
rect 10431 7993 10457 7999
rect 10431 7961 10457 7967
rect 10655 7993 10681 7999
rect 10655 7961 10681 7967
rect 10823 7993 10849 7999
rect 10823 7961 10849 7967
rect 7351 7937 7377 7943
rect 7351 7905 7377 7911
rect 10375 7937 10401 7943
rect 11825 7911 11831 7937
rect 11857 7911 11863 7937
rect 10375 7905 10401 7911
rect 672 7853 20328 7870
rect 672 7827 9919 7853
rect 9945 7827 9971 7853
rect 9997 7827 10023 7853
rect 10049 7827 20328 7853
rect 672 7810 20328 7827
rect 10935 7769 10961 7775
rect 10935 7737 10961 7743
rect 11999 7769 12025 7775
rect 11999 7737 12025 7743
rect 12111 7769 12137 7775
rect 12111 7737 12137 7743
rect 13343 7769 13369 7775
rect 13343 7737 13369 7743
rect 15695 7769 15721 7775
rect 15695 7737 15721 7743
rect 8695 7713 8721 7719
rect 7121 7687 7127 7713
rect 7153 7687 7159 7713
rect 8695 7681 8721 7687
rect 8863 7713 8889 7719
rect 11271 7713 11297 7719
rect 9697 7687 9703 7713
rect 9729 7687 9735 7713
rect 8863 7681 8889 7687
rect 11271 7681 11297 7687
rect 11551 7713 11577 7719
rect 11551 7681 11577 7687
rect 13119 7713 13145 7719
rect 14401 7687 14407 7713
rect 14433 7687 14439 7713
rect 13119 7681 13145 7687
rect 10991 7657 11017 7663
rect 12335 7657 12361 7663
rect 13231 7657 13257 7663
rect 6785 7631 6791 7657
rect 6817 7631 6823 7657
rect 9361 7631 9367 7657
rect 9393 7631 9399 7657
rect 11657 7631 11663 7657
rect 11689 7631 11695 7657
rect 11769 7631 11775 7657
rect 11801 7631 11807 7657
rect 12945 7631 12951 7657
rect 12977 7631 12983 7657
rect 10991 7625 11017 7631
rect 12335 7625 12361 7631
rect 13231 7625 13257 7631
rect 13399 7657 13425 7663
rect 13399 7625 13425 7631
rect 13511 7657 13537 7663
rect 14009 7631 14015 7657
rect 14041 7631 14047 7657
rect 18825 7631 18831 7657
rect 18857 7631 18863 7657
rect 13511 7625 13537 7631
rect 8415 7601 8441 7607
rect 11103 7601 11129 7607
rect 8185 7575 8191 7601
rect 8217 7575 8223 7601
rect 10761 7575 10767 7601
rect 10793 7575 10799 7601
rect 8415 7569 8441 7575
rect 11103 7569 11129 7575
rect 12055 7601 12081 7607
rect 12055 7569 12081 7575
rect 13063 7601 13089 7607
rect 20007 7601 20033 7607
rect 15465 7575 15471 7601
rect 15497 7575 15503 7601
rect 13063 7569 13089 7575
rect 20007 7569 20033 7575
rect 11383 7545 11409 7551
rect 11383 7513 11409 7519
rect 11495 7545 11521 7551
rect 11495 7513 11521 7519
rect 672 7461 20328 7478
rect 672 7435 2239 7461
rect 2265 7435 2291 7461
rect 2317 7435 2343 7461
rect 2369 7435 17599 7461
rect 17625 7435 17651 7461
rect 17677 7435 17703 7461
rect 17729 7435 20328 7461
rect 672 7418 20328 7435
rect 9031 7321 9057 7327
rect 9031 7289 9057 7295
rect 10207 7321 10233 7327
rect 10207 7289 10233 7295
rect 10879 7321 10905 7327
rect 12273 7295 12279 7321
rect 12305 7295 12311 7321
rect 13337 7295 13343 7321
rect 13369 7295 13375 7321
rect 10879 7289 10905 7295
rect 9143 7265 9169 7271
rect 9143 7233 9169 7239
rect 9927 7265 9953 7271
rect 9927 7233 9953 7239
rect 11439 7265 11465 7271
rect 11439 7233 11465 7239
rect 11775 7265 11801 7271
rect 11937 7239 11943 7265
rect 11969 7239 11975 7265
rect 11775 7233 11801 7239
rect 11495 7153 11521 7159
rect 9305 7127 9311 7153
rect 9337 7127 9343 7153
rect 11495 7121 11521 7127
rect 11551 7153 11577 7159
rect 11551 7121 11577 7127
rect 13567 7153 13593 7159
rect 13567 7121 13593 7127
rect 672 7069 20328 7086
rect 672 7043 9919 7069
rect 9945 7043 9971 7069
rect 9997 7043 10023 7069
rect 10049 7043 20328 7069
rect 672 7026 20328 7043
rect 12727 6985 12753 6991
rect 12727 6953 12753 6959
rect 14743 6985 14769 6991
rect 14743 6953 14769 6959
rect 12167 6929 12193 6935
rect 10705 6903 10711 6929
rect 10737 6903 10743 6929
rect 12167 6897 12193 6903
rect 12279 6929 12305 6935
rect 12279 6897 12305 6903
rect 12839 6929 12865 6935
rect 13449 6903 13455 6929
rect 13481 6903 13487 6929
rect 12839 6897 12865 6903
rect 11999 6873 12025 6879
rect 10369 6847 10375 6873
rect 10401 6847 10407 6873
rect 11999 6841 12025 6847
rect 12559 6873 12585 6879
rect 13113 6847 13119 6873
rect 13145 6847 13151 6873
rect 12559 6841 12585 6847
rect 12111 6817 12137 6823
rect 11769 6791 11775 6817
rect 11801 6791 11807 6817
rect 12111 6785 12137 6791
rect 12671 6817 12697 6823
rect 14513 6791 14519 6817
rect 14545 6791 14551 6817
rect 12671 6785 12697 6791
rect 672 6677 20328 6694
rect 672 6651 2239 6677
rect 2265 6651 2291 6677
rect 2317 6651 2343 6677
rect 2369 6651 17599 6677
rect 17625 6651 17651 6677
rect 17677 6651 17703 6677
rect 17729 6651 20328 6677
rect 672 6634 20328 6651
rect 9815 6537 9841 6543
rect 12783 6537 12809 6543
rect 8465 6511 8471 6537
rect 8497 6511 8503 6537
rect 9529 6511 9535 6537
rect 9561 6511 9567 6537
rect 11489 6511 11495 6537
rect 11521 6511 11527 6537
rect 12553 6511 12559 6537
rect 12585 6511 12591 6537
rect 9815 6505 9841 6511
rect 12783 6505 12809 6511
rect 8129 6455 8135 6481
rect 8161 6455 8167 6481
rect 11097 6455 11103 6481
rect 11129 6455 11135 6481
rect 672 6285 20328 6302
rect 672 6259 9919 6285
rect 9945 6259 9971 6285
rect 9997 6259 10023 6285
rect 10049 6259 20328 6285
rect 672 6242 20328 6259
rect 11943 6201 11969 6207
rect 11943 6169 11969 6175
rect 672 5893 20328 5910
rect 672 5867 2239 5893
rect 2265 5867 2291 5893
rect 2317 5867 2343 5893
rect 2369 5867 17599 5893
rect 17625 5867 17651 5893
rect 17677 5867 17703 5893
rect 17729 5867 20328 5893
rect 672 5850 20328 5867
rect 672 5501 20328 5518
rect 672 5475 9919 5501
rect 9945 5475 9971 5501
rect 9997 5475 10023 5501
rect 10049 5475 20328 5501
rect 672 5458 20328 5475
rect 672 5109 20328 5126
rect 672 5083 2239 5109
rect 2265 5083 2291 5109
rect 2317 5083 2343 5109
rect 2369 5083 17599 5109
rect 17625 5083 17651 5109
rect 17677 5083 17703 5109
rect 17729 5083 20328 5109
rect 672 5066 20328 5083
rect 672 4717 20328 4734
rect 672 4691 9919 4717
rect 9945 4691 9971 4717
rect 9997 4691 10023 4717
rect 10049 4691 20328 4717
rect 672 4674 20328 4691
rect 672 4325 20328 4342
rect 672 4299 2239 4325
rect 2265 4299 2291 4325
rect 2317 4299 2343 4325
rect 2369 4299 17599 4325
rect 17625 4299 17651 4325
rect 17677 4299 17703 4325
rect 17729 4299 20328 4325
rect 672 4282 20328 4299
rect 672 3933 20328 3950
rect 672 3907 9919 3933
rect 9945 3907 9971 3933
rect 9997 3907 10023 3933
rect 10049 3907 20328 3933
rect 672 3890 20328 3907
rect 672 3541 20328 3558
rect 672 3515 2239 3541
rect 2265 3515 2291 3541
rect 2317 3515 2343 3541
rect 2369 3515 17599 3541
rect 17625 3515 17651 3541
rect 17677 3515 17703 3541
rect 17729 3515 20328 3541
rect 672 3498 20328 3515
rect 672 3149 20328 3166
rect 672 3123 9919 3149
rect 9945 3123 9971 3149
rect 9997 3123 10023 3149
rect 10049 3123 20328 3149
rect 672 3106 20328 3123
rect 672 2757 20328 2774
rect 672 2731 2239 2757
rect 2265 2731 2291 2757
rect 2317 2731 2343 2757
rect 2369 2731 17599 2757
rect 17625 2731 17651 2757
rect 17677 2731 17703 2757
rect 17729 2731 20328 2757
rect 672 2714 20328 2731
rect 13399 2617 13425 2623
rect 13399 2585 13425 2591
rect 12889 2535 12895 2561
rect 12921 2535 12927 2561
rect 672 2365 20328 2382
rect 672 2339 9919 2365
rect 9945 2339 9971 2365
rect 9997 2339 10023 2365
rect 10049 2339 20328 2365
rect 672 2322 20328 2339
rect 12609 2143 12615 2169
rect 12641 2143 12647 2169
rect 13119 2057 13145 2063
rect 13119 2025 13145 2031
rect 672 1973 20328 1990
rect 672 1947 2239 1973
rect 2265 1947 2291 1973
rect 2317 1947 2343 1973
rect 2369 1947 17599 1973
rect 17625 1947 17651 1973
rect 17677 1947 17703 1973
rect 17729 1947 20328 1973
rect 672 1930 20328 1947
rect 11215 1833 11241 1839
rect 11215 1801 11241 1807
rect 12783 1833 12809 1839
rect 12783 1801 12809 1807
rect 8521 1751 8527 1777
rect 8553 1751 8559 1777
rect 10817 1751 10823 1777
rect 10849 1751 10855 1777
rect 12273 1751 12279 1777
rect 12305 1751 12311 1777
rect 9031 1665 9057 1671
rect 9031 1633 9057 1639
rect 672 1581 20328 1598
rect 672 1555 9919 1581
rect 9945 1555 9971 1581
rect 9997 1555 10023 1581
rect 10049 1555 20328 1581
rect 672 1538 20328 1555
<< via1 >>
rect 2239 19195 2265 19221
rect 2291 19195 2317 19221
rect 2343 19195 2369 19221
rect 17599 19195 17625 19221
rect 17651 19195 17677 19221
rect 17703 19195 17729 19221
rect 8975 19111 9001 19137
rect 11047 19111 11073 19137
rect 12783 19111 12809 19137
rect 8471 18999 8497 19025
rect 10543 18999 10569 19025
rect 12279 18999 12305 19025
rect 9919 18803 9945 18829
rect 9971 18803 9997 18829
rect 10023 18803 10049 18829
rect 10039 18719 10065 18745
rect 13735 18719 13761 18745
rect 9591 18607 9617 18633
rect 13231 18607 13257 18633
rect 2239 18411 2265 18437
rect 2291 18411 2317 18437
rect 2343 18411 2369 18437
rect 17599 18411 17625 18437
rect 17651 18411 17677 18437
rect 17703 18411 17729 18437
rect 8359 18327 8385 18353
rect 8079 18215 8105 18241
rect 9919 18019 9945 18045
rect 9971 18019 9997 18045
rect 10023 18019 10049 18045
rect 2239 17627 2265 17653
rect 2291 17627 2317 17653
rect 2343 17627 2369 17653
rect 17599 17627 17625 17653
rect 17651 17627 17677 17653
rect 17703 17627 17729 17653
rect 9919 17235 9945 17261
rect 9971 17235 9997 17261
rect 10023 17235 10049 17261
rect 2239 16843 2265 16869
rect 2291 16843 2317 16869
rect 2343 16843 2369 16869
rect 17599 16843 17625 16869
rect 17651 16843 17677 16869
rect 17703 16843 17729 16869
rect 9919 16451 9945 16477
rect 9971 16451 9997 16477
rect 10023 16451 10049 16477
rect 2239 16059 2265 16085
rect 2291 16059 2317 16085
rect 2343 16059 2369 16085
rect 17599 16059 17625 16085
rect 17651 16059 17677 16085
rect 17703 16059 17729 16085
rect 9919 15667 9945 15693
rect 9971 15667 9997 15693
rect 10023 15667 10049 15693
rect 2239 15275 2265 15301
rect 2291 15275 2317 15301
rect 2343 15275 2369 15301
rect 17599 15275 17625 15301
rect 17651 15275 17677 15301
rect 17703 15275 17729 15301
rect 9919 14883 9945 14909
rect 9971 14883 9997 14909
rect 10023 14883 10049 14909
rect 2239 14491 2265 14517
rect 2291 14491 2317 14517
rect 2343 14491 2369 14517
rect 17599 14491 17625 14517
rect 17651 14491 17677 14517
rect 17703 14491 17729 14517
rect 8247 14183 8273 14209
rect 9919 14099 9945 14125
rect 9971 14099 9997 14125
rect 10023 14099 10049 14125
rect 8247 14015 8273 14041
rect 8415 14015 8441 14041
rect 12671 13959 12697 13985
rect 6679 13903 6705 13929
rect 8975 13903 9001 13929
rect 12615 13903 12641 13929
rect 18831 13903 18857 13929
rect 7015 13847 7041 13873
rect 8079 13847 8105 13873
rect 9367 13847 9393 13873
rect 10431 13847 10457 13873
rect 10655 13847 10681 13873
rect 13735 13847 13761 13873
rect 12671 13791 12697 13817
rect 13679 13791 13705 13817
rect 20007 13791 20033 13817
rect 2239 13707 2265 13733
rect 2291 13707 2317 13733
rect 2343 13707 2369 13733
rect 17599 13707 17625 13733
rect 17651 13707 17677 13733
rect 17703 13707 17729 13733
rect 7407 13623 7433 13649
rect 7575 13567 7601 13593
rect 7799 13567 7825 13593
rect 9591 13567 9617 13593
rect 10263 13567 10289 13593
rect 12055 13567 12081 13593
rect 13119 13567 13145 13593
rect 8135 13511 8161 13537
rect 9871 13511 9897 13537
rect 11215 13511 11241 13537
rect 11719 13511 11745 13537
rect 7463 13455 7489 13481
rect 7855 13455 7881 13481
rect 7967 13455 7993 13481
rect 8527 13455 8553 13481
rect 9759 13455 9785 13481
rect 11495 13455 11521 13481
rect 9815 13399 9841 13425
rect 9983 13399 10009 13425
rect 11383 13399 11409 13425
rect 11551 13399 11577 13425
rect 13343 13399 13369 13425
rect 9919 13315 9945 13341
rect 9971 13315 9997 13341
rect 10023 13315 10049 13341
rect 8975 13231 9001 13257
rect 9479 13231 9505 13257
rect 9703 13175 9729 13201
rect 10375 13175 10401 13201
rect 7575 13119 7601 13145
rect 8863 13119 8889 13145
rect 9031 13119 9057 13145
rect 9143 13119 9169 13145
rect 9367 13119 9393 13145
rect 9535 13119 9561 13145
rect 9815 13119 9841 13145
rect 9983 13119 10009 13145
rect 10263 13119 10289 13145
rect 10431 13119 10457 13145
rect 10823 13119 10849 13145
rect 12783 13119 12809 13145
rect 11159 13063 11185 13089
rect 12223 13063 12249 13089
rect 13175 13063 13201 13089
rect 14239 13063 14265 13089
rect 14463 13063 14489 13089
rect 7575 13007 7601 13033
rect 7743 13007 7769 13033
rect 9759 13007 9785 13033
rect 10095 13007 10121 13033
rect 2239 12923 2265 12949
rect 2291 12923 2317 12949
rect 2343 12923 2369 12949
rect 17599 12923 17625 12949
rect 17651 12923 17677 12949
rect 17703 12923 17729 12949
rect 967 12783 993 12809
rect 6735 12783 6761 12809
rect 12223 12783 12249 12809
rect 12559 12783 12585 12809
rect 13119 12783 13145 12809
rect 20007 12783 20033 12809
rect 2143 12727 2169 12753
rect 8135 12727 8161 12753
rect 8359 12727 8385 12753
rect 11327 12727 11353 12753
rect 11495 12727 11521 12753
rect 12503 12727 12529 12753
rect 13063 12727 13089 12753
rect 18831 12727 18857 12753
rect 7799 12671 7825 12697
rect 8527 12671 8553 12697
rect 12391 12671 12417 12697
rect 12615 12671 12641 12697
rect 12839 12671 12865 12697
rect 13119 12671 13145 12697
rect 13791 12671 13817 12697
rect 13847 12671 13873 12697
rect 8751 12615 8777 12641
rect 11439 12615 11465 12641
rect 12951 12615 12977 12641
rect 13959 12615 13985 12641
rect 9919 12531 9945 12557
rect 9971 12531 9997 12557
rect 10023 12531 10049 12557
rect 7295 12447 7321 12473
rect 12111 12447 12137 12473
rect 2143 12335 2169 12361
rect 7239 12335 7265 12361
rect 7351 12335 7377 12361
rect 7575 12335 7601 12361
rect 9535 12335 9561 12361
rect 12223 12335 12249 12361
rect 13623 12335 13649 12361
rect 7463 12279 7489 12305
rect 9871 12279 9897 12305
rect 10935 12279 10961 12305
rect 11159 12279 11185 12305
rect 13959 12279 13985 12305
rect 15023 12279 15049 12305
rect 15247 12279 15273 12305
rect 967 12223 993 12249
rect 2239 12139 2265 12165
rect 2291 12139 2317 12165
rect 2343 12139 2369 12165
rect 17599 12139 17625 12165
rect 17651 12139 17677 12165
rect 17703 12139 17729 12165
rect 967 11999 993 12025
rect 9647 11999 9673 12025
rect 20007 11999 20033 12025
rect 2031 11943 2057 11969
rect 7015 11943 7041 11969
rect 8863 11943 8889 11969
rect 9591 11943 9617 11969
rect 9815 11943 9841 11969
rect 9871 11943 9897 11969
rect 14071 11943 14097 11969
rect 18831 11943 18857 11969
rect 6903 11887 6929 11913
rect 8695 11887 8721 11913
rect 8975 11887 9001 11913
rect 9703 11887 9729 11913
rect 10655 11887 10681 11913
rect 11215 11887 11241 11913
rect 12503 11887 12529 11913
rect 13791 11887 13817 11913
rect 13903 11887 13929 11913
rect 7295 11831 7321 11857
rect 8751 11831 8777 11857
rect 10823 11831 10849 11857
rect 11383 11831 11409 11857
rect 11551 11831 11577 11857
rect 11719 11831 11745 11857
rect 12671 11831 12697 11857
rect 13959 11831 13985 11857
rect 9919 11747 9945 11773
rect 9971 11747 9997 11773
rect 10023 11747 10049 11773
rect 9031 11663 9057 11689
rect 9255 11663 9281 11689
rect 10095 11663 10121 11689
rect 10655 11663 10681 11689
rect 7127 11607 7153 11633
rect 7239 11607 7265 11633
rect 7351 11607 7377 11633
rect 7687 11607 7713 11633
rect 9871 11607 9897 11633
rect 10487 11607 10513 11633
rect 11663 11607 11689 11633
rect 2143 11551 2169 11577
rect 6903 11551 6929 11577
rect 7463 11551 7489 11577
rect 9143 11551 9169 11577
rect 10263 11551 10289 11577
rect 11495 11551 11521 11577
rect 13399 11551 13425 11577
rect 5503 11495 5529 11521
rect 6567 11495 6593 11521
rect 7631 11495 7657 11521
rect 9087 11495 9113 11521
rect 9535 11495 9561 11521
rect 10823 11495 10849 11521
rect 13735 11495 13761 11521
rect 14799 11495 14825 11521
rect 15023 11495 15049 11521
rect 967 11439 993 11465
rect 7575 11439 7601 11465
rect 9759 11439 9785 11465
rect 9927 11439 9953 11465
rect 10879 11439 10905 11465
rect 2239 11355 2265 11381
rect 2291 11355 2317 11381
rect 2343 11355 2369 11381
rect 17599 11355 17625 11381
rect 17651 11355 17677 11381
rect 17703 11355 17729 11381
rect 7127 11271 7153 11297
rect 9311 11271 9337 11297
rect 7687 11215 7713 11241
rect 8751 11215 8777 11241
rect 10823 11215 10849 11241
rect 12671 11215 12697 11241
rect 13903 11215 13929 11241
rect 20007 11215 20033 11241
rect 6791 11159 6817 11185
rect 9143 11159 9169 11185
rect 9479 11159 9505 11185
rect 10375 11159 10401 11185
rect 10767 11159 10793 11185
rect 11271 11159 11297 11185
rect 13175 11159 13201 11185
rect 13399 11159 13425 11185
rect 13511 11159 13537 11185
rect 13623 11159 13649 11185
rect 18831 11159 18857 11185
rect 6847 11103 6873 11129
rect 6903 11103 6929 11129
rect 9591 11103 9617 11129
rect 9983 11103 10009 11129
rect 10207 11103 10233 11129
rect 11047 11103 11073 11129
rect 11607 11103 11633 11129
rect 12839 11103 12865 11129
rect 12895 11103 12921 11129
rect 13007 11103 13033 11129
rect 13847 11103 13873 11129
rect 13959 11103 13985 11129
rect 10151 11047 10177 11073
rect 13455 11047 13481 11073
rect 9919 10963 9945 10989
rect 9971 10963 9997 10989
rect 10023 10963 10049 10989
rect 11551 10879 11577 10905
rect 11495 10823 11521 10849
rect 12615 10823 12641 10849
rect 12951 10823 12977 10849
rect 13119 10823 13145 10849
rect 13343 10823 13369 10849
rect 2143 10767 2169 10793
rect 11327 10767 11353 10793
rect 11663 10767 11689 10793
rect 12727 10767 12753 10793
rect 13791 10767 13817 10793
rect 14015 10767 14041 10793
rect 9479 10711 9505 10737
rect 13287 10711 13313 10737
rect 13847 10711 13873 10737
rect 14407 10711 14433 10737
rect 15471 10711 15497 10737
rect 15695 10711 15721 10737
rect 967 10655 993 10681
rect 13623 10655 13649 10681
rect 13679 10655 13705 10681
rect 2239 10571 2265 10597
rect 2291 10571 2317 10597
rect 2343 10571 2369 10597
rect 17599 10571 17625 10597
rect 17651 10571 17677 10597
rect 17703 10571 17729 10597
rect 8471 10487 8497 10513
rect 8695 10487 8721 10513
rect 8863 10487 8889 10513
rect 9871 10487 9897 10513
rect 4999 10431 5025 10457
rect 8975 10431 9001 10457
rect 9255 10431 9281 10457
rect 14127 10431 14153 10457
rect 20007 10431 20033 10457
rect 6399 10375 6425 10401
rect 6735 10375 6761 10401
rect 9311 10375 9337 10401
rect 9591 10375 9617 10401
rect 9703 10375 9729 10401
rect 9815 10375 9841 10401
rect 10431 10375 10457 10401
rect 10655 10375 10681 10401
rect 13567 10375 13593 10401
rect 14071 10375 14097 10401
rect 14239 10375 14265 10401
rect 18831 10375 18857 10401
rect 6063 10319 6089 10345
rect 6847 10319 6873 10345
rect 6903 10319 6929 10345
rect 6959 10319 6985 10345
rect 8415 10319 8441 10345
rect 8471 10319 8497 10345
rect 12559 10319 12585 10345
rect 6791 10263 6817 10289
rect 13455 10263 13481 10289
rect 9919 10179 9945 10205
rect 9971 10179 9997 10205
rect 10023 10179 10049 10205
rect 9255 10095 9281 10121
rect 10879 10095 10905 10121
rect 6119 10039 6145 10065
rect 6231 10039 6257 10065
rect 8863 10039 8889 10065
rect 10207 10039 10233 10065
rect 11047 10039 11073 10065
rect 12279 10039 12305 10065
rect 2143 9983 2169 10009
rect 6791 9983 6817 10009
rect 8919 9983 8945 10009
rect 9087 9983 9113 10009
rect 9703 9983 9729 10009
rect 10655 9983 10681 10009
rect 10767 9983 10793 10009
rect 11215 9983 11241 10009
rect 12223 9983 12249 10009
rect 12615 9983 12641 10009
rect 6063 9927 6089 9953
rect 6567 9927 6593 9953
rect 7183 9927 7209 9953
rect 8247 9927 8273 9953
rect 9423 9927 9449 9953
rect 9927 9927 9953 9953
rect 10823 9927 10849 9953
rect 14463 9927 14489 9953
rect 967 9871 993 9897
rect 12279 9871 12305 9897
rect 2239 9787 2265 9813
rect 2291 9787 2317 9813
rect 2343 9787 2369 9813
rect 17599 9787 17625 9813
rect 17651 9787 17677 9813
rect 17703 9787 17729 9813
rect 10655 9703 10681 9729
rect 10823 9703 10849 9729
rect 13175 9703 13201 9729
rect 14127 9703 14153 9729
rect 4943 9647 4969 9673
rect 9759 9647 9785 9673
rect 12615 9647 12641 9673
rect 13063 9647 13089 9673
rect 6399 9591 6425 9617
rect 6735 9591 6761 9617
rect 8919 9591 8945 9617
rect 9367 9591 9393 9617
rect 9647 9591 9673 9617
rect 10207 9591 10233 9617
rect 10655 9591 10681 9617
rect 12111 9591 12137 9617
rect 12727 9591 12753 9617
rect 13511 9591 13537 9617
rect 13847 9591 13873 9617
rect 14015 9591 14041 9617
rect 14239 9591 14265 9617
rect 6007 9535 6033 9561
rect 6903 9535 6929 9561
rect 9143 9535 9169 9561
rect 9703 9535 9729 9561
rect 10991 9535 11017 9561
rect 11159 9535 11185 9561
rect 11775 9535 11801 9561
rect 12055 9535 12081 9561
rect 14295 9535 14321 9561
rect 14575 9535 14601 9561
rect 6847 9479 6873 9505
rect 8359 9479 8385 9505
rect 8751 9479 8777 9505
rect 8863 9479 8889 9505
rect 9367 9479 9393 9505
rect 11719 9479 11745 9505
rect 12895 9479 12921 9505
rect 13343 9479 13369 9505
rect 13735 9479 13761 9505
rect 13791 9479 13817 9505
rect 14631 9479 14657 9505
rect 14687 9479 14713 9505
rect 9919 9395 9945 9421
rect 9971 9395 9997 9421
rect 10023 9395 10049 9421
rect 9703 9311 9729 9337
rect 6175 9255 6201 9281
rect 7799 9255 7825 9281
rect 8303 9255 8329 9281
rect 9871 9255 9897 9281
rect 10319 9255 10345 9281
rect 11439 9255 11465 9281
rect 11551 9255 11577 9281
rect 11775 9255 11801 9281
rect 12055 9255 12081 9281
rect 13007 9255 13033 9281
rect 13567 9255 13593 9281
rect 14407 9255 14433 9281
rect 6231 9199 6257 9225
rect 6343 9199 6369 9225
rect 6455 9199 6481 9225
rect 7407 9199 7433 9225
rect 7743 9199 7769 9225
rect 8639 9199 8665 9225
rect 8807 9199 8833 9225
rect 9031 9199 9057 9225
rect 9535 9199 9561 9225
rect 10151 9199 10177 9225
rect 11159 9199 11185 9225
rect 11383 9199 11409 9225
rect 12111 9199 12137 9225
rect 12951 9199 12977 9225
rect 13511 9199 13537 9225
rect 14015 9199 14041 9225
rect 6679 9143 6705 9169
rect 8919 9143 8945 9169
rect 9479 9143 9505 9169
rect 13063 9143 13089 9169
rect 15471 9143 15497 9169
rect 15695 9143 15721 9169
rect 7239 9087 7265 9113
rect 8247 9087 8273 9113
rect 8415 9087 8441 9113
rect 11271 9087 11297 9113
rect 2239 9003 2265 9029
rect 2291 9003 2317 9029
rect 2343 9003 2369 9029
rect 17599 9003 17625 9029
rect 17651 9003 17677 9029
rect 17703 9003 17729 9029
rect 6287 8919 6313 8945
rect 7855 8919 7881 8945
rect 8023 8919 8049 8945
rect 13623 8919 13649 8945
rect 967 8863 993 8889
rect 6455 8863 6481 8889
rect 6959 8863 6985 8889
rect 8415 8863 8441 8889
rect 14183 8863 14209 8889
rect 14799 8863 14825 8889
rect 20007 8863 20033 8889
rect 2143 8807 2169 8833
rect 7127 8807 7153 8833
rect 7463 8807 7489 8833
rect 8247 8807 8273 8833
rect 8751 8807 8777 8833
rect 8919 8807 8945 8833
rect 9423 8807 9449 8833
rect 10375 8807 10401 8833
rect 10711 8807 10737 8833
rect 11607 8807 11633 8833
rect 12167 8807 12193 8833
rect 13007 8807 13033 8833
rect 13119 8807 13145 8833
rect 13175 8807 13201 8833
rect 13399 8807 13425 8833
rect 13567 8807 13593 8833
rect 13847 8807 13873 8833
rect 14015 8807 14041 8833
rect 14127 8807 14153 8833
rect 14239 8807 14265 8833
rect 14575 8807 14601 8833
rect 14967 8807 14993 8833
rect 15135 8807 15161 8833
rect 15303 8807 15329 8833
rect 18831 8807 18857 8833
rect 6399 8751 6425 8777
rect 7015 8751 7041 8777
rect 7239 8751 7265 8777
rect 9199 8751 9225 8777
rect 10767 8751 10793 8777
rect 10935 8751 10961 8777
rect 11271 8751 11297 8777
rect 11943 8751 11969 8777
rect 13623 8751 13649 8777
rect 14687 8751 14713 8777
rect 14855 8751 14881 8777
rect 6959 8695 6985 8721
rect 7407 8695 7433 8721
rect 7911 8695 7937 8721
rect 8695 8695 8721 8721
rect 9591 8695 9617 8721
rect 10207 8695 10233 8721
rect 11439 8695 11465 8721
rect 11775 8695 11801 8721
rect 11831 8695 11857 8721
rect 11887 8695 11913 8721
rect 15079 8695 15105 8721
rect 9919 8611 9945 8637
rect 9971 8611 9997 8637
rect 10023 8611 10049 8637
rect 11215 8527 11241 8553
rect 15527 8527 15553 8553
rect 6623 8471 6649 8497
rect 7463 8471 7489 8497
rect 11159 8471 11185 8497
rect 14239 8471 14265 8497
rect 7015 8415 7041 8441
rect 7239 8415 7265 8441
rect 7631 8415 7657 8441
rect 7799 8415 7825 8441
rect 7911 8415 7937 8441
rect 8135 8415 8161 8441
rect 8303 8415 8329 8441
rect 8919 8415 8945 8441
rect 9199 8415 9225 8441
rect 11327 8415 11353 8441
rect 13903 8415 13929 8441
rect 18831 8415 18857 8441
rect 5559 8359 5585 8385
rect 7687 8359 7713 8385
rect 8247 8359 8273 8385
rect 15303 8359 15329 8385
rect 20007 8359 20033 8385
rect 8023 8303 8049 8329
rect 2239 8219 2265 8245
rect 2291 8219 2317 8245
rect 2343 8219 2369 8245
rect 17599 8219 17625 8245
rect 17651 8219 17677 8245
rect 17703 8219 17729 8245
rect 10935 8135 10961 8161
rect 7519 8023 7545 8049
rect 8359 8023 8385 8049
rect 8639 8023 8665 8049
rect 10095 8023 10121 8049
rect 10263 8023 10289 8049
rect 10711 8023 10737 8049
rect 11047 8023 11073 8049
rect 11663 8023 11689 8049
rect 8695 7967 8721 7993
rect 10431 7967 10457 7993
rect 10655 7967 10681 7993
rect 10823 7967 10849 7993
rect 7351 7911 7377 7937
rect 10375 7911 10401 7937
rect 11831 7911 11857 7937
rect 9919 7827 9945 7853
rect 9971 7827 9997 7853
rect 10023 7827 10049 7853
rect 10935 7743 10961 7769
rect 11999 7743 12025 7769
rect 12111 7743 12137 7769
rect 13343 7743 13369 7769
rect 15695 7743 15721 7769
rect 7127 7687 7153 7713
rect 8695 7687 8721 7713
rect 8863 7687 8889 7713
rect 9703 7687 9729 7713
rect 11271 7687 11297 7713
rect 11551 7687 11577 7713
rect 13119 7687 13145 7713
rect 14407 7687 14433 7713
rect 6791 7631 6817 7657
rect 9367 7631 9393 7657
rect 10991 7631 11017 7657
rect 11663 7631 11689 7657
rect 11775 7631 11801 7657
rect 12335 7631 12361 7657
rect 12951 7631 12977 7657
rect 13231 7631 13257 7657
rect 13399 7631 13425 7657
rect 13511 7631 13537 7657
rect 14015 7631 14041 7657
rect 18831 7631 18857 7657
rect 8191 7575 8217 7601
rect 8415 7575 8441 7601
rect 10767 7575 10793 7601
rect 11103 7575 11129 7601
rect 12055 7575 12081 7601
rect 13063 7575 13089 7601
rect 15471 7575 15497 7601
rect 20007 7575 20033 7601
rect 11383 7519 11409 7545
rect 11495 7519 11521 7545
rect 2239 7435 2265 7461
rect 2291 7435 2317 7461
rect 2343 7435 2369 7461
rect 17599 7435 17625 7461
rect 17651 7435 17677 7461
rect 17703 7435 17729 7461
rect 9031 7295 9057 7321
rect 10207 7295 10233 7321
rect 10879 7295 10905 7321
rect 12279 7295 12305 7321
rect 13343 7295 13369 7321
rect 9143 7239 9169 7265
rect 9927 7239 9953 7265
rect 11439 7239 11465 7265
rect 11775 7239 11801 7265
rect 11943 7239 11969 7265
rect 9311 7127 9337 7153
rect 11495 7127 11521 7153
rect 11551 7127 11577 7153
rect 13567 7127 13593 7153
rect 9919 7043 9945 7069
rect 9971 7043 9997 7069
rect 10023 7043 10049 7069
rect 12727 6959 12753 6985
rect 14743 6959 14769 6985
rect 10711 6903 10737 6929
rect 12167 6903 12193 6929
rect 12279 6903 12305 6929
rect 12839 6903 12865 6929
rect 13455 6903 13481 6929
rect 10375 6847 10401 6873
rect 11999 6847 12025 6873
rect 12559 6847 12585 6873
rect 13119 6847 13145 6873
rect 11775 6791 11801 6817
rect 12111 6791 12137 6817
rect 12671 6791 12697 6817
rect 14519 6791 14545 6817
rect 2239 6651 2265 6677
rect 2291 6651 2317 6677
rect 2343 6651 2369 6677
rect 17599 6651 17625 6677
rect 17651 6651 17677 6677
rect 17703 6651 17729 6677
rect 8471 6511 8497 6537
rect 9535 6511 9561 6537
rect 9815 6511 9841 6537
rect 11495 6511 11521 6537
rect 12559 6511 12585 6537
rect 12783 6511 12809 6537
rect 8135 6455 8161 6481
rect 11103 6455 11129 6481
rect 9919 6259 9945 6285
rect 9971 6259 9997 6285
rect 10023 6259 10049 6285
rect 11943 6175 11969 6201
rect 2239 5867 2265 5893
rect 2291 5867 2317 5893
rect 2343 5867 2369 5893
rect 17599 5867 17625 5893
rect 17651 5867 17677 5893
rect 17703 5867 17729 5893
rect 9919 5475 9945 5501
rect 9971 5475 9997 5501
rect 10023 5475 10049 5501
rect 2239 5083 2265 5109
rect 2291 5083 2317 5109
rect 2343 5083 2369 5109
rect 17599 5083 17625 5109
rect 17651 5083 17677 5109
rect 17703 5083 17729 5109
rect 9919 4691 9945 4717
rect 9971 4691 9997 4717
rect 10023 4691 10049 4717
rect 2239 4299 2265 4325
rect 2291 4299 2317 4325
rect 2343 4299 2369 4325
rect 17599 4299 17625 4325
rect 17651 4299 17677 4325
rect 17703 4299 17729 4325
rect 9919 3907 9945 3933
rect 9971 3907 9997 3933
rect 10023 3907 10049 3933
rect 2239 3515 2265 3541
rect 2291 3515 2317 3541
rect 2343 3515 2369 3541
rect 17599 3515 17625 3541
rect 17651 3515 17677 3541
rect 17703 3515 17729 3541
rect 9919 3123 9945 3149
rect 9971 3123 9997 3149
rect 10023 3123 10049 3149
rect 2239 2731 2265 2757
rect 2291 2731 2317 2757
rect 2343 2731 2369 2757
rect 17599 2731 17625 2757
rect 17651 2731 17677 2757
rect 17703 2731 17729 2757
rect 13399 2591 13425 2617
rect 12895 2535 12921 2561
rect 9919 2339 9945 2365
rect 9971 2339 9997 2365
rect 10023 2339 10049 2365
rect 12615 2143 12641 2169
rect 13119 2031 13145 2057
rect 2239 1947 2265 1973
rect 2291 1947 2317 1973
rect 2343 1947 2369 1973
rect 17599 1947 17625 1973
rect 17651 1947 17677 1973
rect 17703 1947 17729 1973
rect 11215 1807 11241 1833
rect 12783 1807 12809 1833
rect 8527 1751 8553 1777
rect 10823 1751 10849 1777
rect 12279 1751 12305 1777
rect 9031 1639 9057 1665
rect 9919 1555 9945 1581
rect 9971 1555 9997 1581
rect 10023 1555 10049 1581
<< metal2 >>
rect 7728 20600 7784 21000
rect 8064 20600 8120 21000
rect 9408 20600 9464 21000
rect 10416 20600 10472 21000
rect 12096 20600 12152 21000
rect 13104 20600 13160 21000
rect 2238 19222 2370 19227
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2238 19189 2370 19194
rect 2238 18438 2370 18443
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2238 18405 2370 18410
rect 7742 18354 7770 20600
rect 8078 19138 8106 20600
rect 8078 19105 8106 19110
rect 8974 19138 9002 19143
rect 8974 19091 9002 19110
rect 8470 19025 8498 19031
rect 8470 18999 8471 19025
rect 8497 18999 8498 19025
rect 7742 18321 7770 18326
rect 8358 18354 8386 18359
rect 8358 18307 8386 18326
rect 8078 18241 8106 18247
rect 8078 18215 8079 18241
rect 8105 18215 8106 18241
rect 2238 17654 2370 17659
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2238 17621 2370 17626
rect 2238 16870 2370 16875
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2238 16837 2370 16842
rect 2238 16086 2370 16091
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2238 16053 2370 16058
rect 2238 15302 2370 15307
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2238 15269 2370 15274
rect 2238 14518 2370 14523
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2238 14485 2370 14490
rect 8078 14098 8106 18215
rect 8470 15974 8498 18999
rect 9422 18746 9450 20600
rect 10430 19138 10458 20600
rect 10430 19105 10458 19110
rect 11046 19138 11074 19143
rect 11046 19091 11074 19110
rect 12110 19138 12138 20600
rect 12110 19105 12138 19110
rect 12782 19138 12810 19143
rect 12782 19091 12810 19110
rect 10542 19025 10570 19031
rect 10542 18999 10543 19025
rect 10569 18999 10570 19025
rect 9918 18830 10050 18835
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 9918 18797 10050 18802
rect 9422 18713 9450 18718
rect 10038 18746 10066 18751
rect 10038 18699 10066 18718
rect 8414 15946 8498 15974
rect 9590 18633 9618 18639
rect 9590 18607 9591 18633
rect 9617 18607 9618 18633
rect 8246 14210 8274 14215
rect 8246 14209 8330 14210
rect 8246 14183 8247 14209
rect 8273 14183 8330 14209
rect 8246 14182 8330 14183
rect 8246 14177 8274 14182
rect 8078 14070 8274 14098
rect 6678 13930 6706 13935
rect 6678 13883 6706 13902
rect 7014 13874 7042 13879
rect 8078 13874 8106 14070
rect 8246 14041 8274 14070
rect 8246 14015 8247 14041
rect 8273 14015 8274 14041
rect 8246 14009 8274 14015
rect 7014 13873 7434 13874
rect 7014 13847 7015 13873
rect 7041 13847 7434 13873
rect 7014 13846 7434 13847
rect 7014 13841 7042 13846
rect 2238 13734 2370 13739
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2238 13701 2370 13706
rect 7406 13649 7434 13846
rect 7406 13623 7407 13649
rect 7433 13623 7434 13649
rect 7406 13617 7434 13623
rect 7854 13873 8106 13874
rect 7854 13847 8079 13873
rect 8105 13847 8106 13873
rect 7854 13846 8106 13847
rect 7574 13594 7602 13599
rect 7798 13594 7826 13599
rect 7574 13593 7826 13594
rect 7574 13567 7575 13593
rect 7601 13567 7799 13593
rect 7825 13567 7826 13593
rect 7574 13566 7826 13567
rect 7574 13561 7602 13566
rect 7798 13561 7826 13566
rect 2086 13482 2114 13487
rect 966 12809 994 12815
rect 966 12783 967 12809
rect 993 12783 994 12809
rect 966 12474 994 12783
rect 966 12441 994 12446
rect 966 12250 994 12255
rect 966 12203 994 12222
rect 966 12025 994 12031
rect 966 11999 967 12025
rect 993 11999 994 12025
rect 966 11802 994 11999
rect 966 11769 994 11774
rect 2030 11969 2058 11975
rect 2030 11943 2031 11969
rect 2057 11943 2058 11969
rect 2030 11522 2058 11943
rect 2030 11489 2058 11494
rect 966 11466 994 11471
rect 966 11419 994 11438
rect 966 10681 994 10687
rect 966 10655 967 10681
rect 993 10655 994 10681
rect 966 10458 994 10655
rect 966 10425 994 10430
rect 2086 10402 2114 13454
rect 7462 13481 7490 13487
rect 7462 13455 7463 13481
rect 7489 13455 7490 13481
rect 2238 12950 2370 12955
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2238 12917 2370 12922
rect 6734 12809 6762 12815
rect 6734 12783 6735 12809
rect 6761 12783 6762 12809
rect 2142 12754 2170 12759
rect 2142 12707 2170 12726
rect 6734 12754 6762 12783
rect 6734 12721 6762 12726
rect 7294 12698 7322 12703
rect 7294 12473 7322 12670
rect 7294 12447 7295 12473
rect 7321 12447 7322 12473
rect 7294 12441 7322 12447
rect 2142 12362 2170 12367
rect 2142 12315 2170 12334
rect 6902 12362 6930 12367
rect 7238 12362 7266 12367
rect 2238 12166 2370 12171
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2238 12133 2370 12138
rect 6902 11913 6930 12334
rect 7182 12361 7266 12362
rect 7182 12335 7239 12361
rect 7265 12335 7266 12361
rect 7182 12334 7266 12335
rect 7126 12250 7154 12255
rect 6902 11887 6903 11913
rect 6929 11887 6930 11913
rect 6902 11881 6930 11887
rect 7014 11969 7042 11975
rect 7014 11943 7015 11969
rect 7041 11943 7042 11969
rect 2142 11746 2170 11751
rect 2142 11577 2170 11718
rect 7014 11634 7042 11943
rect 7014 11601 7042 11606
rect 7126 11633 7154 12222
rect 7126 11607 7127 11633
rect 7153 11607 7154 11633
rect 7126 11601 7154 11607
rect 6902 11578 6930 11583
rect 2142 11551 2143 11577
rect 2169 11551 2170 11577
rect 2142 11545 2170 11551
rect 6734 11550 6902 11578
rect 5502 11522 5530 11527
rect 5502 11475 5530 11494
rect 6566 11522 6594 11527
rect 6566 11475 6594 11494
rect 2238 11382 2370 11387
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2238 11349 2370 11354
rect 6734 10962 6762 11550
rect 6902 11531 6930 11550
rect 7126 11466 7154 11471
rect 7126 11297 7154 11438
rect 7126 11271 7127 11297
rect 7153 11271 7154 11297
rect 7126 11265 7154 11271
rect 6790 11214 6986 11242
rect 6790 11185 6818 11214
rect 6790 11159 6791 11185
rect 6817 11159 6818 11185
rect 6790 11153 6818 11159
rect 6678 10934 6762 10962
rect 6846 11129 6874 11135
rect 6846 11103 6847 11129
rect 6873 11103 6874 11129
rect 2142 10794 2170 10799
rect 2142 10747 2170 10766
rect 4998 10794 5026 10799
rect 2238 10598 2370 10603
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2238 10565 2370 10570
rect 2086 10369 2114 10374
rect 4998 10457 5026 10766
rect 4998 10431 4999 10457
rect 5025 10431 5026 10457
rect 4998 10346 5026 10431
rect 6398 10401 6426 10407
rect 6398 10375 6399 10401
rect 6425 10375 6426 10401
rect 4998 10313 5026 10318
rect 6062 10345 6090 10351
rect 6062 10319 6063 10345
rect 6089 10319 6090 10345
rect 2142 10010 2170 10015
rect 2142 9963 2170 9982
rect 4942 10010 4970 10015
rect 966 9898 994 9903
rect 966 9851 994 9870
rect 2238 9814 2370 9819
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2238 9781 2370 9786
rect 4942 9673 4970 9982
rect 6062 9953 6090 10319
rect 6230 10290 6258 10295
rect 6062 9927 6063 9953
rect 6089 9927 6090 9953
rect 6062 9921 6090 9927
rect 6118 10065 6146 10071
rect 6118 10039 6119 10065
rect 6145 10039 6146 10065
rect 4942 9647 4943 9673
rect 4969 9647 4970 9673
rect 4942 9618 4970 9647
rect 6118 9618 6146 10039
rect 6230 10065 6258 10262
rect 6230 10039 6231 10065
rect 6257 10039 6258 10065
rect 6230 10033 6258 10039
rect 6398 9954 6426 10375
rect 6678 10094 6706 10934
rect 6846 10626 6874 11103
rect 6846 10593 6874 10598
rect 6902 11129 6930 11135
rect 6902 11103 6903 11129
rect 6929 11103 6930 11129
rect 6902 10514 6930 11103
rect 6566 10066 6706 10094
rect 6734 10486 6930 10514
rect 6958 10514 6986 11214
rect 7182 11186 7210 12334
rect 7238 12329 7266 12334
rect 7350 12361 7378 12367
rect 7350 12335 7351 12361
rect 7377 12335 7378 12361
rect 7350 12306 7378 12335
rect 7350 12273 7378 12278
rect 7462 12305 7490 13455
rect 7854 13481 7882 13846
rect 8078 13841 8106 13846
rect 8134 13930 8162 13935
rect 8302 13930 8330 14182
rect 8414 14041 8442 15946
rect 8414 14015 8415 14041
rect 8441 14015 8442 14041
rect 8414 14009 8442 14015
rect 8162 13902 8330 13930
rect 8750 13930 8778 13935
rect 8134 13537 8162 13902
rect 8134 13511 8135 13537
rect 8161 13511 8162 13537
rect 7854 13455 7855 13481
rect 7881 13455 7882 13481
rect 7854 13449 7882 13455
rect 7966 13482 7994 13487
rect 7966 13435 7994 13454
rect 7574 13146 7602 13151
rect 7574 13145 7658 13146
rect 7574 13119 7575 13145
rect 7601 13119 7658 13145
rect 7574 13118 7658 13119
rect 7574 13113 7602 13118
rect 7574 13033 7602 13039
rect 7574 13007 7575 13033
rect 7601 13007 7602 13033
rect 7574 12361 7602 13007
rect 7630 12754 7658 13118
rect 7742 13034 7770 13039
rect 7742 12987 7770 13006
rect 7630 12721 7658 12726
rect 8134 12753 8162 13511
rect 8470 13482 8498 13487
rect 8134 12727 8135 12753
rect 8161 12727 8162 12753
rect 8134 12721 8162 12727
rect 8358 13034 8386 13039
rect 8358 12754 8386 13006
rect 8358 12707 8386 12726
rect 7798 12698 7826 12703
rect 8470 12698 8498 13454
rect 8526 13481 8554 13487
rect 8526 13455 8527 13481
rect 8553 13455 8554 13481
rect 8526 13258 8554 13455
rect 8526 13225 8554 13230
rect 8526 12698 8554 12703
rect 8470 12697 8554 12698
rect 8470 12671 8527 12697
rect 8553 12671 8554 12697
rect 8470 12670 8554 12671
rect 7798 12651 7826 12670
rect 8526 12665 8554 12670
rect 8750 12642 8778 13902
rect 8974 13930 9002 13935
rect 8974 13883 9002 13902
rect 9366 13873 9394 13879
rect 9366 13847 9367 13873
rect 9393 13847 9394 13873
rect 9086 13482 9114 13487
rect 9366 13454 9394 13847
rect 9590 13594 9618 18607
rect 9918 18046 10050 18051
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 9918 18013 10050 18018
rect 9918 17262 10050 17267
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 9918 17229 10050 17234
rect 9918 16478 10050 16483
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 9918 16445 10050 16450
rect 10542 15974 10570 18999
rect 12278 19025 12306 19031
rect 12278 18999 12279 19025
rect 12305 18999 12306 19025
rect 12278 15974 12306 18999
rect 13118 18746 13146 20600
rect 17598 19222 17730 19227
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17598 19189 17730 19194
rect 13118 18713 13146 18718
rect 13734 18746 13762 18751
rect 13734 18699 13762 18718
rect 13230 18633 13258 18639
rect 13230 18607 13231 18633
rect 13257 18607 13258 18633
rect 13230 15974 13258 18607
rect 17598 18438 17730 18443
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17598 18405 17730 18410
rect 17598 17654 17730 17659
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17598 17621 17730 17626
rect 17598 16870 17730 16875
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17598 16837 17730 16842
rect 17598 16086 17730 16091
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17598 16053 17730 16058
rect 10430 15946 10570 15974
rect 12222 15946 12306 15974
rect 13118 15946 13258 15974
rect 9918 15694 10050 15699
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 9918 15661 10050 15666
rect 9918 14910 10050 14915
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 9918 14877 10050 14882
rect 9918 14126 10050 14131
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 9918 14093 10050 14098
rect 10262 13874 10290 13879
rect 9478 13593 9618 13594
rect 9478 13567 9591 13593
rect 9617 13567 9618 13593
rect 9478 13566 9618 13567
rect 9086 13426 9170 13454
rect 9366 13426 9450 13454
rect 8974 13258 9002 13263
rect 8974 13211 9002 13230
rect 8750 12595 8778 12614
rect 8862 13145 8890 13151
rect 8862 13119 8863 13145
rect 8889 13119 8890 13145
rect 7574 12335 7575 12361
rect 7601 12335 7602 12361
rect 7574 12329 7602 12335
rect 7462 12279 7463 12305
rect 7489 12279 7490 12305
rect 7462 12250 7490 12279
rect 7462 12217 7490 12222
rect 8862 11969 8890 13119
rect 9030 13146 9058 13151
rect 9030 13099 9058 13118
rect 9142 13145 9170 13426
rect 9142 13119 9143 13145
rect 9169 13119 9170 13145
rect 8862 11943 8863 11969
rect 8889 11943 8890 11969
rect 8694 11913 8722 11919
rect 8694 11887 8695 11913
rect 8721 11887 8722 11913
rect 7294 11857 7322 11863
rect 7294 11831 7295 11857
rect 7321 11831 7322 11857
rect 7238 11634 7266 11639
rect 7238 11587 7266 11606
rect 7294 11578 7322 11831
rect 7350 11634 7378 11639
rect 7350 11587 7378 11606
rect 7686 11634 7714 11639
rect 7686 11587 7714 11606
rect 7294 11545 7322 11550
rect 7462 11577 7490 11583
rect 7462 11551 7463 11577
rect 7489 11551 7490 11577
rect 7070 11158 7210 11186
rect 6734 10401 6762 10486
rect 6734 10375 6735 10401
rect 6761 10375 6762 10401
rect 6734 10094 6762 10375
rect 6846 10346 6874 10351
rect 6846 10299 6874 10318
rect 6902 10345 6930 10351
rect 6902 10319 6903 10345
rect 6929 10319 6930 10345
rect 6790 10290 6818 10295
rect 6790 10243 6818 10262
rect 6902 10234 6930 10319
rect 6958 10345 6986 10486
rect 6958 10319 6959 10345
rect 6985 10319 6986 10345
rect 6958 10313 6986 10319
rect 7014 10570 7042 10575
rect 7014 10234 7042 10542
rect 6902 10206 7042 10234
rect 7070 10094 7098 11158
rect 7462 11130 7490 11551
rect 7630 11522 7658 11527
rect 7630 11475 7658 11494
rect 7574 11466 7602 11471
rect 7574 11419 7602 11438
rect 7686 11466 7714 11471
rect 7686 11241 7714 11438
rect 7686 11215 7687 11241
rect 7713 11215 7714 11241
rect 7686 11209 7714 11215
rect 7462 11097 7490 11102
rect 8526 10570 8554 10575
rect 8470 10514 8498 10519
rect 8470 10467 8498 10486
rect 8414 10345 8442 10351
rect 8414 10319 8415 10345
rect 8441 10319 8442 10345
rect 7182 10290 7210 10295
rect 6734 10066 6930 10094
rect 7070 10066 7154 10094
rect 6566 9954 6594 10066
rect 6678 10010 6706 10066
rect 6790 10010 6818 10015
rect 6678 10009 6818 10010
rect 6678 9983 6791 10009
rect 6817 9983 6818 10009
rect 6678 9982 6818 9983
rect 6790 9977 6818 9982
rect 6398 9953 6594 9954
rect 6398 9927 6567 9953
rect 6593 9927 6594 9953
rect 6398 9926 6594 9927
rect 6118 9590 6258 9618
rect 4942 9585 4970 9590
rect 6006 9562 6034 9567
rect 6006 9561 6202 9562
rect 6006 9535 6007 9561
rect 6033 9535 6202 9561
rect 6006 9534 6202 9535
rect 6006 9529 6034 9534
rect 6174 9281 6202 9534
rect 6174 9255 6175 9281
rect 6201 9255 6202 9281
rect 6174 9249 6202 9255
rect 6230 9338 6258 9590
rect 6398 9617 6426 9926
rect 6566 9921 6594 9926
rect 6398 9591 6399 9617
rect 6425 9591 6426 9617
rect 6398 9506 6426 9591
rect 6734 9618 6762 9623
rect 6734 9571 6762 9590
rect 6902 9561 6930 10066
rect 6902 9535 6903 9561
rect 6929 9535 6930 9561
rect 6398 9473 6426 9478
rect 6678 9506 6706 9511
rect 6230 9226 6258 9310
rect 6342 9282 6370 9287
rect 6230 9225 6314 9226
rect 6230 9199 6231 9225
rect 6257 9199 6314 9225
rect 6230 9198 6314 9199
rect 6230 9193 6258 9198
rect 2238 9030 2370 9035
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2238 8997 2370 9002
rect 6286 8945 6314 9198
rect 6342 9225 6370 9254
rect 6342 9199 6343 9225
rect 6369 9199 6370 9225
rect 6342 9193 6370 9199
rect 6454 9226 6482 9231
rect 6454 9179 6482 9198
rect 6286 8919 6287 8945
rect 6313 8919 6314 8945
rect 6286 8913 6314 8919
rect 6678 9169 6706 9478
rect 6846 9505 6874 9511
rect 6846 9479 6847 9505
rect 6873 9479 6874 9505
rect 6846 9282 6874 9479
rect 6846 9249 6874 9254
rect 6678 9143 6679 9169
rect 6705 9143 6706 9169
rect 966 8889 994 8895
rect 966 8863 967 8889
rect 993 8863 994 8889
rect 966 8442 994 8863
rect 6398 8890 6426 8895
rect 2142 8834 2170 8839
rect 2142 8787 2170 8806
rect 5558 8834 5586 8839
rect 966 8409 994 8414
rect 5558 8385 5586 8806
rect 6398 8777 6426 8862
rect 6454 8890 6482 8895
rect 6454 8889 6650 8890
rect 6454 8863 6455 8889
rect 6481 8863 6650 8889
rect 6454 8862 6650 8863
rect 6454 8857 6482 8862
rect 6398 8751 6399 8777
rect 6425 8751 6426 8777
rect 6398 8745 6426 8751
rect 6622 8497 6650 8862
rect 6622 8471 6623 8497
rect 6649 8471 6650 8497
rect 6622 8465 6650 8471
rect 6678 8442 6706 9143
rect 6902 8834 6930 9535
rect 7126 9226 7154 10066
rect 7182 9953 7210 10262
rect 8414 10010 8442 10319
rect 8470 10346 8498 10351
rect 8526 10346 8554 10542
rect 8694 10513 8722 11887
rect 8750 11857 8778 11863
rect 8750 11831 8751 11857
rect 8777 11831 8778 11857
rect 8750 11241 8778 11831
rect 8862 11410 8890 11943
rect 9030 12754 9058 12759
rect 8974 11913 9002 11919
rect 8974 11887 8975 11913
rect 9001 11887 9002 11913
rect 8974 11522 9002 11887
rect 9030 11690 9058 12726
rect 9142 11914 9170 13119
rect 9366 13146 9394 13151
rect 9366 13099 9394 13118
rect 9422 13034 9450 13426
rect 9478 13257 9506 13566
rect 9590 13561 9618 13566
rect 9870 13818 9898 13823
rect 9870 13537 9898 13790
rect 10262 13593 10290 13846
rect 10430 13873 10458 15946
rect 10430 13847 10431 13873
rect 10457 13847 10458 13873
rect 10430 13818 10458 13847
rect 10654 13874 10682 13879
rect 10654 13827 10682 13846
rect 10430 13785 10458 13790
rect 12054 13818 12082 13823
rect 10262 13567 10263 13593
rect 10289 13567 10290 13593
rect 10262 13561 10290 13567
rect 12054 13593 12082 13790
rect 12054 13567 12055 13593
rect 12081 13567 12082 13593
rect 12054 13561 12082 13567
rect 11214 13538 11242 13543
rect 9870 13511 9871 13537
rect 9897 13511 9898 13537
rect 9870 13505 9898 13511
rect 11102 13537 11242 13538
rect 11102 13511 11215 13537
rect 11241 13511 11242 13537
rect 11102 13510 11242 13511
rect 9758 13482 9786 13487
rect 9758 13435 9786 13454
rect 9478 13231 9479 13257
rect 9505 13231 9506 13257
rect 9478 13225 9506 13231
rect 9534 13426 9562 13431
rect 9422 13001 9450 13006
rect 9534 13145 9562 13398
rect 9814 13425 9842 13431
rect 9814 13399 9815 13425
rect 9841 13399 9842 13425
rect 9814 13258 9842 13399
rect 9870 13426 9898 13431
rect 9982 13426 10010 13431
rect 9898 13425 10010 13426
rect 9898 13399 9983 13425
rect 10009 13399 10010 13425
rect 9898 13398 10010 13399
rect 9870 13393 9898 13398
rect 9982 13393 10010 13398
rect 9918 13342 10050 13347
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 9918 13309 10050 13314
rect 9758 13230 9842 13258
rect 9702 13202 9730 13207
rect 9758 13202 9786 13230
rect 9702 13201 9786 13202
rect 9702 13175 9703 13201
rect 9729 13175 9786 13201
rect 9702 13174 9786 13175
rect 10374 13201 10402 13207
rect 10374 13175 10375 13201
rect 10401 13175 10402 13201
rect 9702 13169 9730 13174
rect 9534 13119 9535 13145
rect 9561 13119 9562 13145
rect 9534 12698 9562 13119
rect 9814 13145 9842 13151
rect 9814 13119 9815 13145
rect 9841 13119 9842 13145
rect 9758 13034 9786 13039
rect 9758 12987 9786 13006
rect 9142 11881 9170 11886
rect 9478 12670 9562 12698
rect 9254 11690 9282 11695
rect 9030 11689 9226 11690
rect 9030 11663 9031 11689
rect 9057 11663 9226 11689
rect 9030 11662 9226 11663
rect 9030 11657 9058 11662
rect 9142 11577 9170 11583
rect 9142 11551 9143 11577
rect 9169 11551 9170 11577
rect 8974 11489 9002 11494
rect 9086 11521 9114 11527
rect 9086 11495 9087 11521
rect 9113 11495 9114 11521
rect 8862 11377 8890 11382
rect 9086 11298 9114 11495
rect 9142 11466 9170 11551
rect 9142 11433 9170 11438
rect 8750 11215 8751 11241
rect 8777 11215 8778 11241
rect 8750 11209 8778 11215
rect 8862 11270 9114 11298
rect 8694 10487 8695 10513
rect 8721 10487 8722 10513
rect 8694 10481 8722 10487
rect 8862 10513 8890 11270
rect 9142 11185 9170 11191
rect 9142 11159 9143 11185
rect 9169 11159 9170 11185
rect 9142 11130 9170 11159
rect 9142 11097 9170 11102
rect 8862 10487 8863 10513
rect 8889 10487 8890 10513
rect 8862 10481 8890 10487
rect 8974 10514 9002 10519
rect 8974 10457 9002 10486
rect 8974 10431 8975 10457
rect 9001 10431 9002 10457
rect 8974 10425 9002 10431
rect 8470 10345 8554 10346
rect 8470 10319 8471 10345
rect 8497 10319 8554 10345
rect 8470 10318 8554 10319
rect 9198 10346 9226 11662
rect 9254 11643 9282 11662
rect 9478 11634 9506 12670
rect 9478 11601 9506 11606
rect 9534 12586 9562 12591
rect 9534 12361 9562 12558
rect 9534 12335 9535 12361
rect 9561 12335 9562 12361
rect 9534 12306 9562 12335
rect 9534 11521 9562 12278
rect 9590 12362 9618 12367
rect 9814 12362 9842 13119
rect 9982 13146 10010 13151
rect 10262 13146 10290 13151
rect 9982 13145 10290 13146
rect 9982 13119 9983 13145
rect 10009 13119 10263 13145
rect 10289 13119 10290 13145
rect 9982 13118 10290 13119
rect 9982 13113 10010 13118
rect 10262 13113 10290 13118
rect 10094 13033 10122 13039
rect 10094 13007 10095 13033
rect 10121 13007 10122 13033
rect 9918 12558 10050 12563
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 9918 12525 10050 12530
rect 10094 12474 10122 13007
rect 10374 12642 10402 13175
rect 10374 12609 10402 12614
rect 10430 13145 10458 13151
rect 10430 13119 10431 13145
rect 10457 13119 10458 13145
rect 9618 12334 9842 12362
rect 10038 12446 10122 12474
rect 9590 11970 9618 12334
rect 9870 12306 9898 12311
rect 9646 12305 9898 12306
rect 9646 12279 9871 12305
rect 9897 12279 9898 12305
rect 9646 12278 9898 12279
rect 9646 12025 9674 12278
rect 9870 12273 9898 12278
rect 9646 11999 9647 12025
rect 9673 11999 9674 12025
rect 9646 11993 9674 11999
rect 9814 11970 9842 11975
rect 9590 11923 9618 11942
rect 9758 11969 9842 11970
rect 9758 11943 9815 11969
rect 9841 11943 9842 11969
rect 9758 11942 9842 11943
rect 9702 11914 9730 11919
rect 9702 11867 9730 11886
rect 9758 11578 9786 11942
rect 9814 11937 9842 11942
rect 9870 11970 9898 11975
rect 10038 11970 10066 12446
rect 10430 12250 10458 13119
rect 10822 13146 10850 13151
rect 10822 13099 10850 13118
rect 9870 11969 10066 11970
rect 9870 11943 9871 11969
rect 9897 11943 10066 11969
rect 9870 11942 10066 11943
rect 10150 12222 10458 12250
rect 10934 12305 10962 12311
rect 10934 12279 10935 12305
rect 10961 12279 10962 12305
rect 9870 11858 9898 11942
rect 9534 11495 9535 11521
rect 9561 11495 9562 11521
rect 9310 11410 9338 11415
rect 9534 11410 9562 11495
rect 9310 11297 9338 11382
rect 9310 11271 9311 11297
rect 9337 11271 9338 11297
rect 9310 11265 9338 11271
rect 9366 11382 9562 11410
rect 9646 11550 9786 11578
rect 9814 11830 9898 11858
rect 9366 11130 9394 11382
rect 9478 11186 9506 11191
rect 9478 11185 9562 11186
rect 9478 11159 9479 11185
rect 9505 11159 9562 11185
rect 9478 11158 9562 11159
rect 9478 11153 9506 11158
rect 9366 10738 9394 11102
rect 9478 10738 9506 10743
rect 9366 10737 9506 10738
rect 9366 10711 9479 10737
rect 9505 10711 9506 10737
rect 9366 10710 9506 10711
rect 8470 10313 8498 10318
rect 9198 10122 9226 10318
rect 9254 10457 9282 10463
rect 9254 10431 9255 10457
rect 9281 10431 9282 10457
rect 9254 10290 9282 10431
rect 9254 10257 9282 10262
rect 9310 10401 9338 10407
rect 9310 10375 9311 10401
rect 9337 10375 9338 10401
rect 9254 10122 9282 10127
rect 9198 10121 9282 10122
rect 9198 10095 9255 10121
rect 9281 10095 9282 10121
rect 9198 10094 9282 10095
rect 9254 10089 9282 10094
rect 8862 10066 8890 10071
rect 8862 10019 8890 10038
rect 8918 10010 8946 10015
rect 9086 10010 9114 10015
rect 8442 9982 8498 10010
rect 8414 9977 8442 9982
rect 7182 9927 7183 9953
rect 7209 9927 7210 9953
rect 7182 9226 7210 9927
rect 8246 9953 8274 9959
rect 8246 9927 8247 9953
rect 8273 9927 8274 9953
rect 8246 9562 8274 9927
rect 7798 9282 7826 9287
rect 8246 9282 8274 9534
rect 8358 9506 8386 9511
rect 8358 9459 8386 9478
rect 8302 9282 8330 9287
rect 7798 9281 7882 9282
rect 7798 9255 7799 9281
rect 7825 9255 7882 9281
rect 7798 9254 7882 9255
rect 8246 9281 8386 9282
rect 8246 9255 8303 9281
rect 8329 9255 8386 9281
rect 8246 9254 8386 9255
rect 7798 9249 7826 9254
rect 7406 9226 7434 9231
rect 7182 9225 7434 9226
rect 7182 9199 7407 9225
rect 7433 9199 7434 9225
rect 7182 9198 7434 9199
rect 7126 9170 7154 9198
rect 7406 9193 7434 9198
rect 7742 9226 7770 9231
rect 7126 9142 7266 9170
rect 7238 9113 7266 9142
rect 7238 9087 7239 9113
rect 7265 9087 7266 9113
rect 7238 9081 7266 9087
rect 6958 8890 6986 8895
rect 6958 8843 6986 8862
rect 7126 8890 7154 8895
rect 6902 8801 6930 8806
rect 7126 8833 7154 8862
rect 7742 8890 7770 9198
rect 7126 8807 7127 8833
rect 7153 8807 7154 8833
rect 7126 8801 7154 8807
rect 7462 8834 7490 8839
rect 7462 8787 7490 8806
rect 7014 8778 7042 8783
rect 7014 8731 7042 8750
rect 7238 8778 7266 8783
rect 7238 8731 7266 8750
rect 7742 8778 7770 8862
rect 7742 8745 7770 8750
rect 7798 9002 7826 9007
rect 6958 8721 6986 8727
rect 6958 8695 6959 8721
rect 6985 8695 6986 8721
rect 6958 8554 6986 8695
rect 7406 8721 7434 8727
rect 7406 8695 7407 8721
rect 7433 8695 7434 8721
rect 7406 8666 7434 8695
rect 7182 8638 7434 8666
rect 7630 8722 7658 8727
rect 7182 8554 7210 8638
rect 6958 8526 7210 8554
rect 7462 8498 7490 8503
rect 7462 8451 7490 8470
rect 7014 8442 7042 8447
rect 7238 8442 7266 8447
rect 6678 8441 7266 8442
rect 6678 8415 7015 8441
rect 7041 8415 7239 8441
rect 7265 8415 7266 8441
rect 6678 8414 7266 8415
rect 5558 8359 5559 8385
rect 5585 8359 5586 8385
rect 5558 8353 5586 8359
rect 2238 8246 2370 8251
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2238 8213 2370 8218
rect 6790 7657 6818 7663
rect 6790 7631 6791 7657
rect 6817 7631 6818 7657
rect 6790 7602 6818 7631
rect 6846 7602 6874 7607
rect 6790 7574 6846 7602
rect 6846 7569 6874 7574
rect 7014 7602 7042 8414
rect 7238 8409 7266 8414
rect 7518 8442 7546 8447
rect 7518 8049 7546 8414
rect 7630 8441 7658 8694
rect 7630 8415 7631 8441
rect 7657 8415 7658 8441
rect 7630 8409 7658 8415
rect 7798 8441 7826 8974
rect 7798 8415 7799 8441
rect 7825 8415 7826 8441
rect 7798 8409 7826 8415
rect 7854 8945 7882 9254
rect 8302 9249 8330 9254
rect 8246 9113 8274 9119
rect 8246 9087 8247 9113
rect 8273 9087 8274 9113
rect 7854 8919 7855 8945
rect 7881 8919 7882 8945
rect 7854 8442 7882 8919
rect 8022 9058 8050 9063
rect 8022 8945 8050 9030
rect 8022 8919 8023 8945
rect 8049 8919 8050 8945
rect 8022 8913 8050 8919
rect 8246 8890 8274 9087
rect 8078 8862 8274 8890
rect 7910 8721 7938 8727
rect 7910 8695 7911 8721
rect 7937 8695 7938 8721
rect 7910 8666 7938 8695
rect 8078 8666 8106 8862
rect 8246 8833 8274 8862
rect 8246 8807 8247 8833
rect 8273 8807 8274 8833
rect 8246 8801 8274 8807
rect 7910 8638 8106 8666
rect 8134 8778 8162 8783
rect 7910 8442 7938 8447
rect 7854 8441 7938 8442
rect 7854 8415 7911 8441
rect 7937 8415 7938 8441
rect 7854 8414 7938 8415
rect 7910 8409 7938 8414
rect 8134 8441 8162 8750
rect 8134 8415 8135 8441
rect 8161 8415 8162 8441
rect 8134 8409 8162 8415
rect 8190 8498 8218 8503
rect 7686 8385 7714 8391
rect 7686 8359 7687 8385
rect 7713 8359 7714 8385
rect 7686 8330 7714 8359
rect 8022 8330 8050 8335
rect 7686 8329 8050 8330
rect 7686 8303 8023 8329
rect 8049 8303 8050 8329
rect 7686 8302 8050 8303
rect 8022 8297 8050 8302
rect 7518 8023 7519 8049
rect 7545 8023 7546 8049
rect 7518 8017 7546 8023
rect 7350 7938 7378 7943
rect 7126 7937 7378 7938
rect 7126 7911 7351 7937
rect 7377 7911 7378 7937
rect 7126 7910 7378 7911
rect 7126 7713 7154 7910
rect 7350 7905 7378 7910
rect 7126 7687 7127 7713
rect 7153 7687 7154 7713
rect 7126 7681 7154 7687
rect 7014 7569 7042 7574
rect 8190 7601 8218 8470
rect 8302 8442 8330 8447
rect 8302 8395 8330 8414
rect 8246 8386 8274 8391
rect 8246 8339 8274 8358
rect 8358 8049 8386 9254
rect 8414 9114 8442 9119
rect 8414 9067 8442 9086
rect 8470 9002 8498 9982
rect 8918 10009 9170 10010
rect 8918 9983 8919 10009
rect 8945 9983 9087 10009
rect 9113 9983 9170 10009
rect 8918 9982 9170 9983
rect 8918 9977 8946 9982
rect 9086 9977 9114 9982
rect 8918 9898 8946 9903
rect 8862 9618 8890 9623
rect 8806 9590 8862 9618
rect 8750 9505 8778 9511
rect 8750 9479 8751 9505
rect 8777 9479 8778 9505
rect 8750 9338 8778 9479
rect 8750 9305 8778 9310
rect 8638 9226 8666 9231
rect 8638 9179 8666 9198
rect 8806 9225 8834 9590
rect 8862 9585 8890 9590
rect 8918 9617 8946 9870
rect 8918 9591 8919 9617
rect 8945 9591 8946 9617
rect 8918 9585 8946 9591
rect 9142 9561 9170 9982
rect 9142 9535 9143 9561
rect 9169 9535 9170 9561
rect 8862 9505 8890 9511
rect 8862 9479 8863 9505
rect 8889 9479 8890 9505
rect 8862 9450 8890 9479
rect 8862 9417 8890 9422
rect 8806 9199 8807 9225
rect 8833 9199 8834 9225
rect 8470 8969 8498 8974
rect 8414 8890 8442 8895
rect 8414 8722 8442 8862
rect 8750 8834 8778 8839
rect 8806 8834 8834 9199
rect 9030 9226 9058 9231
rect 9142 9226 9170 9535
rect 9030 9225 9170 9226
rect 9030 9199 9031 9225
rect 9057 9199 9170 9225
rect 9030 9198 9170 9199
rect 9198 9954 9226 9959
rect 9030 9193 9058 9198
rect 8750 8833 8834 8834
rect 8750 8807 8751 8833
rect 8777 8807 8834 8833
rect 8750 8806 8834 8807
rect 8918 9169 8946 9175
rect 8918 9143 8919 9169
rect 8945 9143 8946 9169
rect 8918 9114 8946 9143
rect 8918 8833 8946 9086
rect 8918 8807 8919 8833
rect 8945 8807 8946 8833
rect 8750 8801 8778 8806
rect 8414 8689 8442 8694
rect 8694 8722 8722 8727
rect 8694 8675 8722 8694
rect 8918 8442 8946 8807
rect 8358 8023 8359 8049
rect 8385 8023 8386 8049
rect 8358 8017 8386 8023
rect 8638 8441 8946 8442
rect 8638 8415 8919 8441
rect 8945 8415 8946 8441
rect 8638 8414 8946 8415
rect 8638 8049 8666 8414
rect 8918 8409 8946 8414
rect 8974 9002 9002 9007
rect 8638 8023 8639 8049
rect 8665 8023 8666 8049
rect 8638 8017 8666 8023
rect 8694 7993 8722 7999
rect 8694 7967 8695 7993
rect 8721 7967 8722 7993
rect 8694 7713 8722 7967
rect 8694 7687 8695 7713
rect 8721 7687 8722 7713
rect 8694 7681 8722 7687
rect 8862 7713 8890 7719
rect 8862 7687 8863 7713
rect 8889 7687 8890 7713
rect 8190 7575 8191 7601
rect 8217 7575 8218 7601
rect 8190 7574 8218 7575
rect 8414 7602 8442 7621
rect 8190 7546 8386 7574
rect 8414 7569 8442 7574
rect 8358 7490 8386 7546
rect 2238 7462 2370 7467
rect 8358 7462 8442 7490
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2238 7429 2370 7434
rect 2238 6678 2370 6683
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2238 6645 2370 6650
rect 8134 6538 8162 6543
rect 8134 6481 8162 6510
rect 8134 6455 8135 6481
rect 8161 6455 8162 6481
rect 8134 6449 8162 6455
rect 2238 5894 2370 5899
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2238 5861 2370 5866
rect 2238 5110 2370 5115
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2238 5077 2370 5082
rect 2238 4326 2370 4331
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2238 4293 2370 4298
rect 8414 4214 8442 7462
rect 8470 6538 8498 6543
rect 8862 6538 8890 7687
rect 8974 7322 9002 8974
rect 9198 8777 9226 9926
rect 9310 9674 9338 10375
rect 9422 9954 9450 9959
rect 9254 9646 9338 9674
rect 9366 9953 9450 9954
rect 9366 9927 9423 9953
rect 9449 9927 9450 9953
rect 9366 9926 9450 9927
rect 9254 9170 9282 9646
rect 9366 9618 9394 9926
rect 9422 9921 9450 9926
rect 9310 9590 9366 9618
rect 9310 9282 9338 9590
rect 9366 9585 9394 9590
rect 9366 9505 9394 9511
rect 9366 9479 9367 9505
rect 9393 9479 9394 9505
rect 9366 9450 9394 9479
rect 9422 9506 9450 9511
rect 9478 9506 9506 10710
rect 9534 9898 9562 11158
rect 9590 11129 9618 11135
rect 9590 11103 9591 11129
rect 9617 11103 9618 11129
rect 9590 10570 9618 11103
rect 9590 10537 9618 10542
rect 9534 9865 9562 9870
rect 9590 10401 9618 10407
rect 9590 10375 9591 10401
rect 9617 10375 9618 10401
rect 9450 9478 9506 9506
rect 9422 9473 9450 9478
rect 9366 9338 9394 9422
rect 9366 9310 9506 9338
rect 9478 9282 9506 9310
rect 9310 9254 9450 9282
rect 9254 9137 9282 9142
rect 9422 8833 9450 9254
rect 9478 9249 9506 9254
rect 9534 9226 9562 9231
rect 9590 9226 9618 10375
rect 9646 10178 9674 11550
rect 9758 11466 9786 11471
rect 9814 11466 9842 11830
rect 10094 11802 10122 11807
rect 9918 11774 10050 11779
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 9918 11741 10050 11746
rect 10094 11690 10122 11774
rect 10094 11643 10122 11662
rect 9758 11465 9842 11466
rect 9758 11439 9759 11465
rect 9785 11439 9842 11465
rect 9758 11438 9842 11439
rect 9870 11634 9898 11639
rect 9758 10514 9786 11438
rect 9870 11074 9898 11606
rect 9926 11466 9954 11471
rect 9926 11419 9954 11438
rect 9814 11046 9898 11074
rect 9982 11129 10010 11135
rect 9982 11103 9983 11129
rect 10009 11103 10010 11129
rect 9982 11074 10010 11103
rect 10150 11130 10178 12222
rect 10654 11970 10682 11975
rect 10654 11913 10682 11942
rect 10654 11887 10655 11913
rect 10681 11887 10682 11913
rect 10654 11881 10682 11887
rect 10710 11914 10738 11919
rect 10654 11690 10682 11695
rect 10710 11690 10738 11886
rect 10934 11914 10962 12279
rect 11102 11970 11130 13510
rect 11214 13505 11242 13510
rect 11718 13537 11746 13543
rect 11718 13511 11719 13537
rect 11745 13511 11746 13537
rect 11494 13482 11522 13487
rect 11494 13435 11522 13454
rect 11382 13426 11410 13431
rect 11382 13379 11410 13398
rect 11550 13425 11578 13431
rect 11550 13399 11551 13425
rect 11577 13399 11578 13425
rect 11158 13090 11186 13095
rect 11158 13089 11354 13090
rect 11158 13063 11159 13089
rect 11185 13063 11354 13089
rect 11158 13062 11354 13063
rect 11158 13057 11186 13062
rect 11326 12753 11354 13062
rect 11326 12727 11327 12753
rect 11353 12727 11354 12753
rect 11326 12721 11354 12727
rect 11494 12754 11522 12759
rect 11550 12754 11578 13399
rect 11718 13146 11746 13511
rect 12222 13482 12250 15946
rect 12670 13986 12698 13991
rect 12670 13985 12810 13986
rect 12670 13959 12671 13985
rect 12697 13959 12810 13985
rect 12670 13958 12810 13959
rect 12670 13953 12698 13958
rect 12614 13930 12642 13935
rect 11718 13113 11746 13118
rect 12110 13426 12138 13431
rect 11494 12753 11578 12754
rect 11494 12727 11495 12753
rect 11521 12727 11578 12753
rect 11494 12726 11578 12727
rect 12110 12754 12138 13398
rect 12166 13146 12194 13151
rect 12166 12810 12194 13118
rect 12222 13089 12250 13454
rect 12222 13063 12223 13089
rect 12249 13063 12250 13089
rect 12222 13057 12250 13063
rect 12558 13929 12642 13930
rect 12558 13903 12615 13929
rect 12641 13903 12642 13929
rect 12558 13902 12642 13903
rect 12222 12810 12250 12815
rect 12166 12809 12250 12810
rect 12166 12783 12223 12809
rect 12249 12783 12250 12809
rect 12166 12782 12250 12783
rect 12222 12777 12250 12782
rect 12558 12809 12586 13902
rect 12614 13897 12642 13902
rect 12782 13874 12810 13958
rect 12782 13846 12978 13874
rect 12670 13818 12698 13823
rect 12670 13771 12698 13790
rect 12670 13594 12698 13599
rect 12670 13454 12698 13566
rect 12558 12783 12559 12809
rect 12585 12783 12586 12809
rect 12558 12777 12586 12783
rect 12614 13426 12698 13454
rect 11494 12721 11522 12726
rect 11438 12642 11466 12647
rect 11158 12306 11186 12311
rect 11158 12259 11186 12278
rect 11438 11970 11466 12614
rect 12110 12473 12138 12726
rect 12502 12754 12530 12759
rect 12502 12707 12530 12726
rect 12110 12447 12111 12473
rect 12137 12447 12138 12473
rect 12110 12441 12138 12447
rect 12390 12697 12418 12703
rect 12390 12671 12391 12697
rect 12417 12671 12418 12697
rect 11102 11937 11130 11942
rect 11326 11942 11466 11970
rect 12222 12361 12250 12367
rect 12222 12335 12223 12361
rect 12249 12335 12250 12361
rect 10934 11881 10962 11886
rect 11214 11914 11242 11919
rect 11214 11867 11242 11886
rect 10822 11858 10850 11863
rect 10822 11857 10906 11858
rect 10822 11831 10823 11857
rect 10849 11831 10906 11857
rect 10822 11830 10906 11831
rect 10822 11825 10850 11830
rect 10654 11689 10738 11690
rect 10654 11663 10655 11689
rect 10681 11663 10738 11689
rect 10654 11662 10738 11663
rect 10878 11802 10906 11830
rect 10654 11657 10682 11662
rect 10486 11634 10514 11639
rect 10318 11633 10514 11634
rect 10318 11607 10487 11633
rect 10513 11607 10514 11633
rect 10318 11606 10514 11607
rect 10262 11577 10290 11583
rect 10262 11551 10263 11577
rect 10289 11551 10290 11577
rect 9982 11046 10122 11074
rect 9814 10906 9842 11046
rect 9918 10990 10050 10995
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 9918 10957 10050 10962
rect 10094 10906 10122 11046
rect 10150 11073 10178 11102
rect 10150 11047 10151 11073
rect 10177 11047 10178 11073
rect 10150 11041 10178 11047
rect 10206 11129 10234 11135
rect 10206 11103 10207 11129
rect 10233 11103 10234 11129
rect 9814 10878 9954 10906
rect 9870 10514 9898 10519
rect 9758 10513 9898 10514
rect 9758 10487 9871 10513
rect 9897 10487 9898 10513
rect 9758 10486 9898 10487
rect 9870 10481 9898 10486
rect 9702 10401 9730 10407
rect 9814 10402 9842 10407
rect 9702 10375 9703 10401
rect 9729 10375 9730 10401
rect 9702 10290 9730 10375
rect 9758 10401 9842 10402
rect 9758 10375 9815 10401
rect 9841 10375 9842 10401
rect 9758 10374 9842 10375
rect 9758 10346 9786 10374
rect 9814 10369 9842 10374
rect 9758 10313 9786 10318
rect 9926 10290 9954 10878
rect 9702 10257 9730 10262
rect 9814 10262 9954 10290
rect 10038 10878 10122 10906
rect 10038 10290 10066 10878
rect 10206 10290 10234 11103
rect 10038 10262 10122 10290
rect 9646 10150 9786 10178
rect 9702 10009 9730 10015
rect 9702 9983 9703 10009
rect 9729 9983 9730 10009
rect 9702 9730 9730 9983
rect 9702 9697 9730 9702
rect 9758 9674 9786 10150
rect 9758 9627 9786 9646
rect 9534 9225 9590 9226
rect 9534 9199 9535 9225
rect 9561 9199 9590 9225
rect 9534 9198 9590 9199
rect 9534 9193 9562 9198
rect 9590 9179 9618 9198
rect 9646 9617 9674 9623
rect 9646 9591 9647 9617
rect 9673 9591 9674 9617
rect 9422 8807 9423 8833
rect 9449 8807 9450 8833
rect 9422 8801 9450 8807
rect 9478 9169 9506 9175
rect 9478 9143 9479 9169
rect 9505 9143 9506 9169
rect 9478 9114 9506 9143
rect 9646 9114 9674 9591
rect 9702 9562 9730 9567
rect 9702 9337 9730 9534
rect 9702 9311 9703 9337
rect 9729 9311 9730 9337
rect 9702 9305 9730 9311
rect 9478 9086 9674 9114
rect 9198 8751 9199 8777
rect 9225 8751 9226 8777
rect 9198 8745 9226 8751
rect 9198 8442 9226 8447
rect 9198 8395 9226 8414
rect 9478 8442 9506 9086
rect 9478 8409 9506 8414
rect 9590 8722 9618 8727
rect 9814 8722 9842 10262
rect 9918 10206 10050 10211
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 9918 10173 10050 10178
rect 9926 9954 9954 9959
rect 9926 9907 9954 9926
rect 10094 9842 10122 10262
rect 10206 10257 10234 10262
rect 10262 10178 10290 11551
rect 10094 9809 10122 9814
rect 10150 10150 10290 10178
rect 10150 9730 10178 10150
rect 10150 9697 10178 9702
rect 10206 10066 10234 10071
rect 10318 10066 10346 11606
rect 10486 11601 10514 11606
rect 10878 11578 10906 11774
rect 10878 11550 10962 11578
rect 10822 11521 10850 11527
rect 10822 11495 10823 11521
rect 10849 11495 10850 11521
rect 10822 11241 10850 11495
rect 10822 11215 10823 11241
rect 10849 11215 10850 11241
rect 10374 11186 10402 11191
rect 10766 11186 10794 11191
rect 10374 11185 10626 11186
rect 10374 11159 10375 11185
rect 10401 11159 10626 11185
rect 10374 11158 10626 11159
rect 10374 11153 10402 11158
rect 10430 10402 10458 10407
rect 10430 10355 10458 10374
rect 10234 10038 10346 10066
rect 10206 9618 10234 10038
rect 10598 10010 10626 11158
rect 10766 11139 10794 11158
rect 10654 10402 10682 10407
rect 10654 10355 10682 10374
rect 10206 9571 10234 9590
rect 10262 9842 10290 9847
rect 9918 9422 10050 9427
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 9918 9389 10050 9394
rect 9870 9281 9898 9287
rect 9870 9255 9871 9281
rect 9897 9255 9898 9281
rect 9870 9170 9898 9255
rect 10150 9226 10178 9231
rect 10150 9179 10178 9198
rect 9870 9137 9898 9142
rect 10262 9114 10290 9814
rect 10598 9730 10626 9982
rect 10654 10009 10682 10015
rect 10654 9983 10655 10009
rect 10681 9983 10682 10009
rect 10654 9842 10682 9983
rect 10654 9809 10682 9814
rect 10766 10009 10794 10015
rect 10766 9983 10767 10009
rect 10793 9983 10794 10009
rect 10654 9730 10682 9735
rect 10598 9729 10682 9730
rect 10598 9703 10655 9729
rect 10681 9703 10682 9729
rect 10598 9702 10682 9703
rect 10654 9697 10682 9702
rect 10654 9618 10682 9623
rect 10654 9571 10682 9590
rect 10766 9562 10794 9983
rect 10822 9953 10850 11215
rect 10878 11465 10906 11471
rect 10878 11439 10879 11465
rect 10905 11439 10906 11465
rect 10878 10850 10906 11439
rect 10878 10817 10906 10822
rect 10934 10738 10962 11550
rect 11046 11522 11074 11527
rect 11326 11522 11354 11942
rect 11382 11858 11410 11863
rect 11382 11578 11410 11830
rect 11550 11857 11578 11863
rect 11550 11831 11551 11857
rect 11577 11831 11578 11857
rect 11550 11802 11578 11831
rect 11718 11857 11746 11863
rect 11718 11831 11719 11857
rect 11745 11831 11746 11857
rect 11718 11802 11746 11831
rect 12222 11858 12250 12335
rect 12222 11825 12250 11830
rect 11998 11802 12026 11807
rect 11718 11774 11998 11802
rect 11550 11769 11578 11774
rect 11662 11634 11690 11639
rect 11606 11633 11690 11634
rect 11606 11607 11663 11633
rect 11689 11607 11690 11633
rect 11606 11606 11690 11607
rect 11494 11578 11522 11583
rect 11382 11577 11522 11578
rect 11382 11551 11495 11577
rect 11521 11551 11522 11577
rect 11382 11550 11522 11551
rect 11326 11494 11410 11522
rect 11046 11129 11074 11494
rect 11046 11103 11047 11129
rect 11073 11103 11074 11129
rect 11046 11018 11074 11103
rect 11046 10985 11074 10990
rect 11102 11242 11130 11247
rect 10878 10710 10962 10738
rect 10878 10121 10906 10710
rect 10878 10095 10879 10121
rect 10905 10095 10906 10121
rect 10878 10089 10906 10095
rect 10822 9927 10823 9953
rect 10849 9927 10850 9953
rect 10822 9921 10850 9927
rect 11046 10066 11074 10071
rect 10822 9730 10850 9735
rect 10822 9683 10850 9702
rect 9590 8721 9842 8722
rect 9590 8695 9591 8721
rect 9617 8695 9842 8721
rect 9590 8694 9842 8695
rect 10150 9086 10290 9114
rect 10318 9281 10346 9287
rect 10318 9255 10319 9281
rect 10345 9255 10346 9281
rect 9590 8050 9618 8694
rect 9918 8638 10050 8643
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 9918 8605 10050 8610
rect 9590 8017 9618 8022
rect 9814 8442 9842 8447
rect 9702 7938 9730 7943
rect 9702 7713 9730 7910
rect 9702 7687 9703 7713
rect 9729 7687 9730 7713
rect 9702 7681 9730 7687
rect 9366 7657 9394 7663
rect 9366 7631 9367 7657
rect 9393 7631 9394 7657
rect 9366 7602 9394 7631
rect 9030 7322 9058 7327
rect 8974 7321 9058 7322
rect 8974 7295 9031 7321
rect 9057 7295 9058 7321
rect 8974 7294 9058 7295
rect 9030 7289 9058 7294
rect 9142 7265 9170 7271
rect 9142 7239 9143 7265
rect 9169 7239 9170 7265
rect 9142 6538 9170 7239
rect 9310 7154 9338 7159
rect 9310 7107 9338 7126
rect 8470 6537 9170 6538
rect 8470 6511 8471 6537
rect 8497 6511 9170 6537
rect 8470 6510 9170 6511
rect 9366 6538 9394 7574
rect 9814 7266 9842 8414
rect 10094 8050 10122 8055
rect 10094 8003 10122 8022
rect 9918 7854 10050 7859
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 9918 7821 10050 7826
rect 10150 7546 10178 9086
rect 10318 8946 10346 9255
rect 10318 8913 10346 8918
rect 10374 9170 10402 9175
rect 10374 8833 10402 9142
rect 10766 9170 10794 9534
rect 10990 9562 11018 9567
rect 10990 9515 11018 9534
rect 10766 9137 10794 9142
rect 10710 8946 10738 8951
rect 10738 8918 10794 8946
rect 10710 8913 10738 8918
rect 10374 8807 10375 8833
rect 10401 8807 10402 8833
rect 10374 8801 10402 8807
rect 10710 8834 10738 8839
rect 10710 8787 10738 8806
rect 10766 8777 10794 8918
rect 11046 8834 11074 10038
rect 11046 8801 11074 8806
rect 10766 8751 10767 8777
rect 10793 8751 10794 8777
rect 10766 8745 10794 8751
rect 10934 8777 10962 8783
rect 10934 8751 10935 8777
rect 10961 8751 10962 8777
rect 10206 8722 10234 8727
rect 10206 8675 10234 8694
rect 10710 8722 10738 8727
rect 10262 8050 10290 8055
rect 10262 8003 10290 8022
rect 10710 8049 10738 8694
rect 10934 8722 10962 8751
rect 10934 8689 10962 8694
rect 11102 8554 11130 11214
rect 11270 11186 11298 11191
rect 11270 11139 11298 11158
rect 11326 10793 11354 10799
rect 11326 10767 11327 10793
rect 11353 10767 11354 10793
rect 11158 10570 11186 10575
rect 11158 9562 11186 10542
rect 11326 10346 11354 10767
rect 11382 10626 11410 11494
rect 11382 10593 11410 10598
rect 11326 10313 11354 10318
rect 11438 10066 11466 11550
rect 11494 11545 11522 11550
rect 11606 11242 11634 11606
rect 11662 11601 11690 11606
rect 11606 11209 11634 11214
rect 11662 11466 11690 11471
rect 11606 11130 11634 11135
rect 11550 11129 11634 11130
rect 11550 11103 11607 11129
rect 11633 11103 11634 11129
rect 11550 11102 11634 11103
rect 11550 10905 11578 11102
rect 11606 11097 11634 11102
rect 11550 10879 11551 10905
rect 11577 10879 11578 10905
rect 11550 10873 11578 10879
rect 11494 10850 11522 10855
rect 11494 10803 11522 10822
rect 11662 10793 11690 11438
rect 11662 10767 11663 10793
rect 11689 10767 11690 10793
rect 11438 10033 11466 10038
rect 11550 10626 11578 10631
rect 11214 10010 11242 10015
rect 11214 9963 11242 9982
rect 11158 9561 11410 9562
rect 11158 9535 11159 9561
rect 11185 9535 11410 9561
rect 11158 9534 11410 9535
rect 11158 9529 11186 9534
rect 11158 9225 11186 9231
rect 11158 9199 11159 9225
rect 11185 9199 11186 9225
rect 11158 9058 11186 9199
rect 11158 9025 11186 9030
rect 10710 8023 10711 8049
rect 10737 8023 10738 8049
rect 10710 8017 10738 8023
rect 10878 8526 11130 8554
rect 11158 8946 11186 8951
rect 10878 8050 10906 8526
rect 11158 8498 11186 8918
rect 11214 8553 11242 9534
rect 11382 9225 11410 9534
rect 11438 9282 11466 9287
rect 11438 9235 11466 9254
rect 11550 9281 11578 10598
rect 11662 10122 11690 10767
rect 11662 10089 11690 10094
rect 11550 9255 11551 9281
rect 11577 9255 11578 9281
rect 11550 9249 11578 9255
rect 11718 10010 11746 10015
rect 11718 9898 11746 9982
rect 11718 9505 11746 9870
rect 11718 9479 11719 9505
rect 11745 9479 11746 9505
rect 11382 9199 11383 9225
rect 11409 9199 11410 9225
rect 11382 9193 11410 9199
rect 11606 9170 11634 9175
rect 11718 9170 11746 9479
rect 11774 9954 11802 9959
rect 11774 9561 11802 9926
rect 11774 9535 11775 9561
rect 11801 9535 11802 9561
rect 11774 9338 11802 9535
rect 11774 9281 11802 9310
rect 11774 9255 11775 9281
rect 11801 9255 11802 9281
rect 11774 9249 11802 9255
rect 11718 9142 11970 9170
rect 11270 9113 11298 9119
rect 11270 9087 11271 9113
rect 11297 9087 11298 9113
rect 11270 8946 11298 9087
rect 11270 8913 11298 8918
rect 11606 8833 11634 9142
rect 11606 8807 11607 8833
rect 11633 8807 11634 8833
rect 11606 8801 11634 8807
rect 11270 8777 11298 8783
rect 11270 8751 11271 8777
rect 11297 8751 11298 8777
rect 11270 8666 11298 8751
rect 11942 8777 11970 9142
rect 11942 8751 11943 8777
rect 11969 8751 11970 8777
rect 11942 8745 11970 8751
rect 11270 8633 11298 8638
rect 11326 8722 11354 8727
rect 11326 8554 11354 8694
rect 11214 8527 11215 8553
rect 11241 8527 11242 8553
rect 11214 8521 11242 8527
rect 11270 8526 11354 8554
rect 11438 8722 11466 8727
rect 10934 8497 11186 8498
rect 10934 8471 11159 8497
rect 11185 8471 11186 8497
rect 10934 8470 11186 8471
rect 10934 8161 10962 8470
rect 11158 8465 11186 8470
rect 10934 8135 10935 8161
rect 10961 8135 10962 8161
rect 10934 8129 10962 8135
rect 10878 8017 10906 8022
rect 11046 8049 11074 8055
rect 11046 8023 11047 8049
rect 11073 8023 11074 8049
rect 10430 7994 10458 7999
rect 10654 7994 10682 7999
rect 10430 7993 10682 7994
rect 10430 7967 10431 7993
rect 10457 7967 10655 7993
rect 10681 7967 10682 7993
rect 10430 7966 10682 7967
rect 10430 7961 10458 7966
rect 10654 7961 10682 7966
rect 10822 7993 10850 7999
rect 10822 7967 10823 7993
rect 10849 7967 10850 7993
rect 10374 7937 10402 7943
rect 10374 7911 10375 7937
rect 10401 7911 10402 7937
rect 10374 7574 10402 7911
rect 10822 7938 10850 7967
rect 10822 7905 10850 7910
rect 10934 7770 10962 7775
rect 10822 7769 10962 7770
rect 10822 7743 10935 7769
rect 10961 7743 10962 7769
rect 10822 7742 10962 7743
rect 10766 7601 10794 7607
rect 10766 7575 10767 7601
rect 10793 7575 10794 7601
rect 10766 7574 10794 7575
rect 10206 7546 10234 7551
rect 10374 7546 10794 7574
rect 10150 7518 10206 7546
rect 10206 7321 10234 7518
rect 10206 7295 10207 7321
rect 10233 7295 10234 7321
rect 10206 7289 10234 7295
rect 9926 7266 9954 7271
rect 8470 6505 8498 6510
rect 9366 6505 9394 6510
rect 9534 7265 9954 7266
rect 9534 7239 9927 7265
rect 9953 7239 9954 7265
rect 9534 7238 9954 7239
rect 9534 6537 9562 7238
rect 9926 7233 9954 7238
rect 9918 7070 10050 7075
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 10766 7042 10794 7546
rect 9918 7037 10050 7042
rect 10654 7014 10794 7042
rect 10374 6873 10402 6879
rect 10374 6847 10375 6873
rect 10401 6847 10402 6873
rect 10374 6762 10402 6847
rect 10374 6729 10402 6734
rect 9534 6511 9535 6537
rect 9561 6511 9562 6537
rect 9534 6505 9562 6511
rect 9814 6538 9842 6543
rect 9814 6491 9842 6510
rect 9918 6286 10050 6291
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 9918 6253 10050 6258
rect 9918 5502 10050 5507
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 9918 5469 10050 5474
rect 9918 4718 10050 4723
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 9918 4685 10050 4690
rect 10654 4214 10682 7014
rect 10710 6930 10738 6935
rect 10822 6930 10850 7742
rect 10934 7737 10962 7742
rect 10990 7770 11018 7775
rect 11046 7770 11074 8023
rect 11018 7742 11074 7770
rect 10990 7657 11018 7742
rect 11270 7713 11298 8526
rect 11326 8442 11354 8447
rect 11326 8395 11354 8414
rect 11438 7770 11466 8694
rect 11774 8721 11802 8727
rect 11774 8695 11775 8721
rect 11801 8695 11802 8721
rect 11774 8442 11802 8695
rect 11774 8409 11802 8414
rect 11830 8721 11858 8727
rect 11830 8695 11831 8721
rect 11857 8695 11858 8721
rect 11830 8162 11858 8695
rect 11886 8722 11914 8727
rect 11998 8722 12026 11774
rect 12390 11802 12418 12671
rect 12614 12697 12642 13426
rect 12782 13146 12810 13151
rect 12782 13099 12810 13118
rect 12614 12671 12615 12697
rect 12641 12671 12642 12697
rect 12614 12665 12642 12671
rect 12838 12697 12866 12703
rect 12838 12671 12839 12697
rect 12865 12671 12866 12697
rect 12502 12250 12530 12255
rect 12502 11913 12530 12222
rect 12838 12250 12866 12671
rect 12950 12642 12978 13846
rect 13062 13818 13090 13823
rect 13062 12753 13090 13790
rect 13118 13594 13146 15946
rect 17598 15302 17730 15307
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17598 15269 17730 15274
rect 17598 14518 17730 14523
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17598 14485 17730 14490
rect 18830 13930 18858 13935
rect 18830 13883 18858 13902
rect 13734 13874 13762 13879
rect 13734 13827 13762 13846
rect 14238 13874 14266 13879
rect 13678 13818 13706 13823
rect 13678 13771 13706 13790
rect 13118 13547 13146 13566
rect 13342 13425 13370 13431
rect 13342 13399 13343 13425
rect 13369 13399 13370 13425
rect 13342 13146 13370 13399
rect 13174 13089 13202 13095
rect 13174 13063 13175 13089
rect 13201 13063 13202 13089
rect 13118 12810 13146 12815
rect 13174 12810 13202 13063
rect 13342 12866 13370 13118
rect 14238 13089 14266 13846
rect 20006 13818 20034 13823
rect 20006 13771 20034 13790
rect 17598 13734 17730 13739
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17598 13701 17730 13706
rect 14238 13063 14239 13089
rect 14265 13063 14266 13089
rect 14238 13057 14266 13063
rect 14462 13089 14490 13095
rect 14462 13063 14463 13089
rect 14489 13063 14490 13089
rect 13342 12833 13370 12838
rect 13622 12866 13650 12871
rect 13118 12809 13202 12810
rect 13118 12783 13119 12809
rect 13145 12783 13202 12809
rect 13118 12782 13202 12783
rect 13118 12777 13146 12782
rect 13062 12727 13063 12753
rect 13089 12727 13090 12753
rect 13062 12721 13090 12727
rect 13118 12698 13146 12703
rect 13118 12651 13146 12670
rect 12838 12217 12866 12222
rect 12894 12641 12978 12642
rect 12894 12615 12951 12641
rect 12977 12615 12978 12641
rect 12894 12614 12978 12615
rect 12502 11887 12503 11913
rect 12529 11887 12530 11913
rect 12502 11881 12530 11887
rect 12670 11858 12698 11863
rect 12670 11857 12810 11858
rect 12670 11831 12671 11857
rect 12697 11831 12810 11857
rect 12670 11830 12810 11831
rect 12670 11825 12698 11830
rect 12390 11769 12418 11774
rect 12670 11242 12698 11247
rect 12670 11241 12754 11242
rect 12670 11215 12671 11241
rect 12697 11215 12754 11241
rect 12670 11214 12754 11215
rect 12670 11209 12698 11214
rect 12614 10849 12642 10855
rect 12614 10823 12615 10849
rect 12641 10823 12642 10849
rect 12614 10402 12642 10823
rect 12726 10793 12754 11214
rect 12782 11074 12810 11830
rect 12782 11041 12810 11046
rect 12838 11129 12866 11135
rect 12838 11103 12839 11129
rect 12865 11103 12866 11129
rect 12726 10767 12727 10793
rect 12753 10767 12754 10793
rect 12726 10738 12754 10767
rect 12726 10705 12754 10710
rect 12614 10374 12754 10402
rect 12558 10346 12586 10351
rect 12586 10318 12642 10346
rect 12558 10299 12586 10318
rect 12278 10066 12306 10071
rect 12278 10019 12306 10038
rect 12222 10009 12250 10015
rect 12222 9983 12223 10009
rect 12249 9983 12250 10009
rect 12222 9954 12250 9983
rect 12614 10009 12642 10318
rect 12614 9983 12615 10009
rect 12641 9983 12642 10009
rect 12614 9977 12642 9983
rect 12054 9926 12222 9954
rect 12054 9561 12082 9926
rect 12222 9921 12250 9926
rect 12670 9954 12698 9959
rect 12278 9898 12306 9903
rect 12278 9851 12306 9870
rect 12110 9842 12138 9847
rect 12110 9617 12138 9814
rect 12614 9674 12642 9679
rect 12670 9674 12698 9926
rect 12726 9730 12754 10374
rect 12782 10122 12810 10127
rect 12782 9898 12810 10094
rect 12838 10010 12866 11103
rect 12894 11130 12922 12614
rect 12950 12609 12978 12614
rect 13622 12362 13650 12838
rect 14462 12866 14490 13063
rect 17598 12950 17730 12955
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17598 12917 17730 12922
rect 14490 12838 15106 12866
rect 14462 12819 14490 12838
rect 13846 12754 13874 12759
rect 13790 12698 13818 12703
rect 13790 12651 13818 12670
rect 13846 12697 13874 12726
rect 13846 12671 13847 12697
rect 13873 12671 13874 12697
rect 13846 12665 13874 12671
rect 14910 12754 14938 12759
rect 13958 12642 13986 12647
rect 13958 12641 14098 12642
rect 13958 12615 13959 12641
rect 13985 12615 14098 12641
rect 13958 12614 14098 12615
rect 13958 12609 13986 12614
rect 13454 12361 13650 12362
rect 13454 12335 13623 12361
rect 13649 12335 13650 12361
rect 13454 12334 13650 12335
rect 13398 11578 13426 11583
rect 13454 11578 13482 12334
rect 13622 12329 13650 12334
rect 13958 12305 13986 12311
rect 13958 12279 13959 12305
rect 13985 12279 13986 12305
rect 13398 11577 13482 11578
rect 13398 11551 13399 11577
rect 13425 11551 13482 11577
rect 13398 11550 13482 11551
rect 13790 11913 13818 11919
rect 13790 11887 13791 11913
rect 13817 11887 13818 11913
rect 13398 11545 13426 11550
rect 13734 11522 13762 11527
rect 13454 11521 13762 11522
rect 13454 11495 13735 11521
rect 13761 11495 13762 11521
rect 13454 11494 13762 11495
rect 13174 11186 13202 11191
rect 13174 11139 13202 11158
rect 13398 11185 13426 11191
rect 13398 11159 13399 11185
rect 13425 11159 13426 11185
rect 12894 11083 12922 11102
rect 13006 11130 13034 11135
rect 13006 11083 13034 11102
rect 13398 11130 13426 11159
rect 13398 11097 13426 11102
rect 13454 11073 13482 11494
rect 13734 11489 13762 11494
rect 13566 11242 13594 11247
rect 13510 11214 13566 11242
rect 13510 11185 13538 11214
rect 13566 11209 13594 11214
rect 13510 11159 13511 11185
rect 13537 11159 13538 11185
rect 13510 11153 13538 11159
rect 13622 11186 13650 11191
rect 13622 11185 13762 11186
rect 13622 11159 13623 11185
rect 13649 11159 13762 11185
rect 13622 11158 13762 11159
rect 13622 11153 13650 11158
rect 13454 11047 13455 11073
rect 13481 11047 13482 11073
rect 13454 11041 13482 11047
rect 13734 11018 13762 11158
rect 12950 10849 12978 10855
rect 12950 10823 12951 10849
rect 12977 10823 12978 10849
rect 12950 10402 12978 10823
rect 13118 10850 13146 10855
rect 13342 10850 13370 10855
rect 13118 10849 13370 10850
rect 13118 10823 13119 10849
rect 13145 10823 13343 10849
rect 13369 10823 13370 10849
rect 13118 10822 13370 10823
rect 13118 10817 13146 10822
rect 13286 10738 13314 10743
rect 13286 10691 13314 10710
rect 13342 10402 13370 10822
rect 13622 10682 13650 10687
rect 13622 10635 13650 10654
rect 13678 10681 13706 10687
rect 13678 10655 13679 10681
rect 13705 10655 13706 10681
rect 13566 10402 13594 10407
rect 12978 10374 13034 10402
rect 13342 10401 13594 10402
rect 13342 10375 13567 10401
rect 13593 10375 13594 10401
rect 13342 10374 13594 10375
rect 12950 10369 12978 10374
rect 12838 9977 12866 9982
rect 12782 9870 12866 9898
rect 12726 9697 12754 9702
rect 12614 9673 12698 9674
rect 12614 9647 12615 9673
rect 12641 9647 12698 9673
rect 12614 9646 12698 9647
rect 12782 9674 12810 9679
rect 12614 9641 12642 9646
rect 12110 9591 12111 9617
rect 12137 9591 12138 9617
rect 12110 9585 12138 9591
rect 12726 9618 12754 9623
rect 12782 9618 12810 9646
rect 12726 9617 12810 9618
rect 12726 9591 12727 9617
rect 12753 9591 12810 9617
rect 12726 9590 12810 9591
rect 12726 9585 12754 9590
rect 12054 9535 12055 9561
rect 12081 9535 12082 9561
rect 12054 9281 12082 9535
rect 12054 9255 12055 9281
rect 12081 9255 12082 9281
rect 12054 9249 12082 9255
rect 12166 9506 12194 9511
rect 12110 9226 12138 9231
rect 12054 8890 12082 8895
rect 12110 8890 12138 9198
rect 12082 8862 12138 8890
rect 12054 8857 12082 8862
rect 12166 8833 12194 9478
rect 12166 8807 12167 8833
rect 12193 8807 12194 8833
rect 12166 8801 12194 8807
rect 11998 8694 12194 8722
rect 11886 8675 11914 8694
rect 11438 7737 11466 7742
rect 11606 8134 11858 8162
rect 11998 8442 12026 8447
rect 11270 7687 11271 7713
rect 11297 7687 11298 7713
rect 11270 7681 11298 7687
rect 11550 7714 11578 7719
rect 11550 7667 11578 7686
rect 10990 7631 10991 7657
rect 11017 7631 11018 7657
rect 10990 7625 11018 7631
rect 10878 7602 10906 7607
rect 10878 7321 10906 7574
rect 11102 7602 11130 7621
rect 11102 7569 11130 7574
rect 11382 7546 11410 7551
rect 11494 7546 11522 7551
rect 11382 7545 11522 7546
rect 11382 7519 11383 7545
rect 11409 7519 11495 7545
rect 11521 7519 11522 7545
rect 11382 7518 11522 7519
rect 11382 7513 11410 7518
rect 11494 7513 11522 7518
rect 11606 7434 11634 8134
rect 11662 8050 11690 8055
rect 11662 8003 11690 8022
rect 11830 7938 11858 7943
rect 11830 7937 11914 7938
rect 11830 7911 11831 7937
rect 11857 7911 11914 7937
rect 11830 7910 11914 7911
rect 11830 7905 11858 7910
rect 11830 7714 11858 7719
rect 11662 7658 11690 7663
rect 11662 7611 11690 7630
rect 11774 7657 11802 7663
rect 11774 7631 11775 7657
rect 11801 7631 11802 7657
rect 11774 7546 11802 7631
rect 11774 7513 11802 7518
rect 10878 7295 10879 7321
rect 10905 7295 10906 7321
rect 10878 7289 10906 7295
rect 11438 7406 11634 7434
rect 11438 7265 11466 7406
rect 11438 7239 11439 7265
rect 11465 7239 11466 7265
rect 11438 7233 11466 7239
rect 11774 7265 11802 7271
rect 11774 7239 11775 7265
rect 11801 7239 11802 7265
rect 10710 6929 10850 6930
rect 10710 6903 10711 6929
rect 10737 6903 10850 6929
rect 10710 6902 10850 6903
rect 11494 7153 11522 7159
rect 11494 7127 11495 7153
rect 11521 7127 11522 7153
rect 10710 6897 10738 6902
rect 11102 6706 11130 6711
rect 11102 6481 11130 6678
rect 11494 6537 11522 7127
rect 11550 7154 11578 7159
rect 11550 7107 11578 7126
rect 11774 7154 11802 7239
rect 11774 7121 11802 7126
rect 11494 6511 11495 6537
rect 11521 6511 11522 6537
rect 11494 6505 11522 6511
rect 11774 6818 11802 6823
rect 11830 6818 11858 7686
rect 11886 7658 11914 7910
rect 11998 7769 12026 8414
rect 11998 7743 11999 7769
rect 12025 7743 12026 7769
rect 11998 7737 12026 7743
rect 12110 7770 12138 7775
rect 12110 7723 12138 7742
rect 11886 7625 11914 7630
rect 12054 7601 12082 7607
rect 12054 7575 12055 7601
rect 12081 7575 12082 7601
rect 11998 7546 12026 7551
rect 11774 6817 11858 6818
rect 11774 6791 11775 6817
rect 11801 6791 11858 6817
rect 11774 6790 11858 6791
rect 11942 7265 11970 7271
rect 11942 7239 11943 7265
rect 11969 7239 11970 7265
rect 11102 6455 11103 6481
rect 11129 6455 11130 6481
rect 11102 6449 11130 6455
rect 11774 4214 11802 6790
rect 11942 6706 11970 7239
rect 11998 6930 12026 7518
rect 12054 7378 12082 7575
rect 12166 7546 12194 8694
rect 12166 7513 12194 7518
rect 12334 7657 12362 7663
rect 12334 7631 12335 7657
rect 12361 7631 12362 7657
rect 12054 7350 12306 7378
rect 12278 7321 12306 7350
rect 12278 7295 12279 7321
rect 12305 7295 12306 7321
rect 12278 7289 12306 7295
rect 11998 6873 12026 6902
rect 11998 6847 11999 6873
rect 12025 6847 12026 6873
rect 11998 6841 12026 6847
rect 12110 7154 12138 7159
rect 12110 6817 12138 7126
rect 12222 6986 12250 6991
rect 12166 6958 12222 6986
rect 12166 6929 12194 6958
rect 12222 6953 12250 6958
rect 12166 6903 12167 6929
rect 12193 6903 12194 6929
rect 12166 6897 12194 6903
rect 12278 6929 12306 6935
rect 12278 6903 12279 6929
rect 12305 6903 12306 6929
rect 12110 6791 12111 6817
rect 12137 6791 12138 6817
rect 12110 6785 12138 6791
rect 11942 6201 11970 6678
rect 12278 6538 12306 6903
rect 12334 6818 12362 7631
rect 12726 7658 12754 7663
rect 12838 7658 12866 9870
rect 12894 9786 12922 9791
rect 12894 9506 12922 9758
rect 12894 9459 12922 9478
rect 13006 9506 13034 10374
rect 13566 10369 13594 10374
rect 13454 10289 13482 10295
rect 13454 10263 13455 10289
rect 13481 10263 13482 10289
rect 13062 10066 13090 10071
rect 13062 9673 13090 10038
rect 13454 9954 13482 10263
rect 13678 10178 13706 10655
rect 13454 9921 13482 9926
rect 13622 10150 13706 10178
rect 13734 10178 13762 10990
rect 13510 9898 13538 9903
rect 13174 9730 13202 9735
rect 13174 9683 13202 9702
rect 13062 9647 13063 9673
rect 13089 9647 13090 9673
rect 13062 9641 13090 9647
rect 13510 9617 13538 9870
rect 13622 9730 13650 10150
rect 13734 10145 13762 10150
rect 13790 10793 13818 11887
rect 13902 11913 13930 11919
rect 13902 11887 13903 11913
rect 13929 11887 13930 11913
rect 13902 11634 13930 11887
rect 13958 11857 13986 12279
rect 14070 11969 14098 12614
rect 14910 12306 14938 12726
rect 15078 12586 15106 12838
rect 20006 12809 20034 12815
rect 20006 12783 20007 12809
rect 20033 12783 20034 12809
rect 18830 12754 18858 12759
rect 18830 12707 18858 12726
rect 15078 12558 15162 12586
rect 15022 12306 15050 12311
rect 14910 12305 15050 12306
rect 14910 12279 15023 12305
rect 15049 12279 15050 12305
rect 14910 12278 15050 12279
rect 15134 12306 15162 12558
rect 20006 12474 20034 12783
rect 20006 12441 20034 12446
rect 15246 12306 15274 12311
rect 15134 12305 15274 12306
rect 15134 12279 15247 12305
rect 15273 12279 15274 12305
rect 15134 12278 15274 12279
rect 15022 12273 15050 12278
rect 14070 11943 14071 11969
rect 14097 11943 14098 11969
rect 14070 11937 14098 11943
rect 13958 11831 13959 11857
rect 13985 11831 13986 11857
rect 13958 11825 13986 11831
rect 13902 11606 14210 11634
rect 14014 11522 14042 11527
rect 13958 11494 14014 11522
rect 13902 11242 13930 11247
rect 13902 11195 13930 11214
rect 13846 11129 13874 11135
rect 13846 11103 13847 11129
rect 13873 11103 13874 11129
rect 13846 11074 13874 11103
rect 13958 11129 13986 11494
rect 14014 11489 14042 11494
rect 13958 11103 13959 11129
rect 13985 11103 13986 11129
rect 13958 11097 13986 11103
rect 14014 11186 14042 11191
rect 13874 11046 13930 11074
rect 13846 11041 13874 11046
rect 13790 10767 13791 10793
rect 13817 10767 13818 10793
rect 13790 10094 13818 10767
rect 13846 10738 13874 10743
rect 13846 10691 13874 10710
rect 13622 9697 13650 9702
rect 13678 10066 13818 10094
rect 13510 9591 13511 9617
rect 13537 9591 13538 9617
rect 13006 9478 13146 9506
rect 12894 9338 12922 9343
rect 12894 8834 12922 9310
rect 13006 9281 13034 9478
rect 13006 9255 13007 9281
rect 13033 9255 13034 9281
rect 13006 9249 13034 9255
rect 13062 9394 13090 9399
rect 12950 9226 12978 9231
rect 12950 9179 12978 9198
rect 13062 9169 13090 9366
rect 13062 9143 13063 9169
rect 13089 9143 13090 9169
rect 13006 8834 13034 8839
rect 12894 8833 13034 8834
rect 12894 8807 13007 8833
rect 13033 8807 13034 8833
rect 12894 8806 13034 8807
rect 13006 8801 13034 8806
rect 13006 8386 13034 8391
rect 13062 8386 13090 9143
rect 13034 8358 13090 8386
rect 13118 8833 13146 9478
rect 13342 9505 13370 9511
rect 13342 9479 13343 9505
rect 13369 9479 13370 9505
rect 13118 8807 13119 8833
rect 13145 8807 13146 8833
rect 13118 8386 13146 8807
rect 13174 9226 13202 9231
rect 13174 8833 13202 9198
rect 13342 9170 13370 9479
rect 13510 9225 13538 9591
rect 13510 9199 13511 9225
rect 13537 9199 13538 9225
rect 13398 9170 13426 9175
rect 13342 9142 13398 9170
rect 13398 9137 13426 9142
rect 13174 8807 13175 8833
rect 13201 8807 13202 8833
rect 13174 8801 13202 8807
rect 13398 8834 13426 8839
rect 13510 8834 13538 9199
rect 13566 9281 13594 9287
rect 13566 9255 13567 9281
rect 13593 9255 13594 9281
rect 13566 9226 13594 9255
rect 13566 9193 13594 9198
rect 13622 8946 13650 8951
rect 13678 8946 13706 10066
rect 13902 9786 13930 11046
rect 14014 10793 14042 11158
rect 14014 10767 14015 10793
rect 14041 10767 14042 10793
rect 14014 9954 14042 10767
rect 14070 10682 14098 10687
rect 14098 10654 14154 10682
rect 14070 10649 14098 10654
rect 14126 10457 14154 10654
rect 14126 10431 14127 10457
rect 14153 10431 14154 10457
rect 14126 10425 14154 10431
rect 14070 10402 14098 10407
rect 14070 10355 14098 10374
rect 14182 10234 14210 11606
rect 14798 11522 14826 11527
rect 14798 11475 14826 11494
rect 15022 11521 15050 11527
rect 15022 11495 15023 11521
rect 15049 11495 15050 11521
rect 15022 11466 15050 11495
rect 15246 11466 15274 12278
rect 17598 12166 17730 12171
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17598 12133 17730 12138
rect 20006 12025 20034 12031
rect 20006 11999 20007 12025
rect 20033 11999 20034 12025
rect 18830 11969 18858 11975
rect 18830 11943 18831 11969
rect 18857 11943 18858 11969
rect 18830 11522 18858 11943
rect 20006 11802 20034 11999
rect 20006 11769 20034 11774
rect 18830 11489 18858 11494
rect 15022 11438 15554 11466
rect 14406 10738 14434 10743
rect 14406 10691 14434 10710
rect 15470 10738 15498 10743
rect 15526 10738 15554 11438
rect 17598 11382 17730 11387
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17598 11349 17730 11354
rect 20006 11241 20034 11247
rect 20006 11215 20007 11241
rect 20033 11215 20034 11241
rect 18830 11185 18858 11191
rect 18830 11159 18831 11185
rect 18857 11159 18858 11185
rect 15694 10738 15722 10743
rect 15526 10737 15722 10738
rect 15526 10711 15695 10737
rect 15721 10711 15722 10737
rect 15526 10710 15722 10711
rect 14238 10402 14266 10407
rect 14238 10355 14266 10374
rect 15470 10402 15498 10710
rect 15470 10369 15498 10374
rect 14014 9921 14042 9926
rect 14070 10206 14210 10234
rect 13846 9618 13874 9623
rect 13902 9618 13930 9758
rect 13846 9617 13930 9618
rect 13846 9591 13847 9617
rect 13873 9591 13930 9617
rect 13846 9590 13930 9591
rect 14014 9617 14042 9623
rect 14014 9591 14015 9617
rect 14041 9591 14042 9617
rect 13846 9585 13874 9590
rect 13734 9506 13762 9511
rect 13734 9459 13762 9478
rect 13790 9506 13818 9511
rect 14014 9506 14042 9591
rect 13790 9505 14042 9506
rect 13790 9479 13791 9505
rect 13817 9479 14042 9505
rect 13790 9478 14042 9479
rect 13790 9473 13818 9478
rect 13846 9338 13874 9343
rect 13622 8945 13706 8946
rect 13622 8919 13623 8945
rect 13649 8919 13706 8945
rect 13622 8918 13706 8919
rect 13734 9226 13762 9231
rect 13622 8913 13650 8918
rect 13566 8834 13594 8839
rect 13510 8833 13594 8834
rect 13510 8807 13567 8833
rect 13593 8807 13594 8833
rect 13510 8806 13594 8807
rect 13398 8787 13426 8806
rect 13566 8801 13594 8806
rect 13622 8778 13650 8783
rect 13734 8778 13762 9198
rect 13846 8833 13874 9310
rect 14014 9282 14042 9287
rect 14014 9226 14042 9254
rect 13846 8807 13847 8833
rect 13873 8807 13874 8833
rect 13846 8801 13874 8807
rect 13958 9225 14042 9226
rect 13958 9199 14015 9225
rect 14041 9199 14042 9225
rect 13958 9198 14042 9199
rect 13622 8777 13762 8778
rect 13622 8751 13623 8777
rect 13649 8751 13762 8777
rect 13622 8750 13762 8751
rect 13622 8745 13650 8750
rect 13902 8442 13930 8447
rect 13958 8442 13986 9198
rect 14014 9193 14042 9198
rect 14014 8834 14042 8839
rect 14014 8787 14042 8806
rect 14070 8666 14098 10206
rect 14182 10122 14210 10127
rect 14126 9730 14154 9735
rect 14182 9730 14210 10094
rect 14126 9729 14210 9730
rect 14126 9703 14127 9729
rect 14153 9703 14210 9729
rect 14126 9702 14210 9703
rect 14462 9954 14490 9959
rect 14126 9697 14154 9702
rect 14238 9617 14266 9623
rect 14238 9591 14239 9617
rect 14265 9591 14266 9617
rect 14182 9562 14210 9567
rect 14126 8890 14154 8895
rect 14126 8833 14154 8862
rect 14182 8889 14210 9534
rect 14238 9338 14266 9591
rect 14294 9562 14322 9567
rect 14294 9561 14434 9562
rect 14294 9535 14295 9561
rect 14321 9535 14434 9561
rect 14294 9534 14434 9535
rect 14294 9529 14322 9534
rect 14238 9305 14266 9310
rect 14406 9281 14434 9534
rect 14406 9255 14407 9281
rect 14433 9255 14434 9281
rect 14406 9249 14434 9255
rect 14462 9282 14490 9926
rect 14574 9562 14602 9567
rect 14574 9515 14602 9534
rect 14462 9249 14490 9254
rect 14630 9505 14658 9511
rect 14630 9479 14631 9505
rect 14657 9479 14658 9505
rect 14182 8863 14183 8889
rect 14209 8863 14210 8889
rect 14182 8857 14210 8863
rect 14238 9170 14266 9175
rect 14126 8807 14127 8833
rect 14153 8807 14154 8833
rect 14126 8801 14154 8807
rect 14238 8833 14266 9142
rect 14238 8807 14239 8833
rect 14265 8807 14266 8833
rect 14238 8722 14266 8807
rect 14574 8834 14602 8839
rect 14574 8787 14602 8806
rect 14238 8689 14266 8694
rect 14070 8633 14098 8638
rect 14630 8554 14658 9479
rect 14686 9505 14714 9511
rect 14686 9479 14687 9505
rect 14713 9479 14714 9505
rect 14686 9394 14714 9479
rect 15470 9506 15498 9511
rect 14686 9361 14714 9366
rect 15246 9394 15274 9399
rect 15274 9366 15330 9394
rect 15246 9361 15274 9366
rect 14798 8890 14826 8895
rect 14798 8889 14994 8890
rect 14798 8863 14799 8889
rect 14825 8863 14994 8889
rect 14798 8862 14994 8863
rect 14798 8857 14826 8862
rect 14966 8833 14994 8862
rect 14966 8807 14967 8833
rect 14993 8807 14994 8833
rect 14966 8801 14994 8807
rect 15134 8833 15162 8839
rect 15134 8807 15135 8833
rect 15161 8807 15162 8833
rect 14686 8778 14714 8783
rect 14686 8731 14714 8750
rect 14854 8777 14882 8783
rect 14854 8751 14855 8777
rect 14881 8751 14882 8777
rect 14854 8722 14882 8751
rect 14854 8689 14882 8694
rect 15078 8721 15106 8727
rect 15078 8695 15079 8721
rect 15105 8695 15106 8721
rect 14406 8526 14658 8554
rect 14238 8498 14266 8503
rect 14238 8451 14266 8470
rect 13902 8441 13986 8442
rect 13902 8415 13903 8441
rect 13929 8415 13986 8441
rect 13902 8414 13986 8415
rect 13006 8353 13034 8358
rect 13118 8353 13146 8358
rect 13510 8386 13538 8391
rect 13342 7770 13370 7775
rect 13118 7769 13370 7770
rect 13118 7743 13343 7769
rect 13369 7743 13370 7769
rect 13118 7742 13370 7743
rect 13118 7713 13146 7742
rect 13342 7737 13370 7742
rect 13118 7687 13119 7713
rect 13145 7687 13146 7713
rect 13118 7681 13146 7687
rect 12950 7658 12978 7663
rect 12838 7657 12978 7658
rect 12838 7631 12951 7657
rect 12977 7631 12978 7657
rect 12838 7630 12978 7631
rect 12726 6986 12754 7630
rect 12950 7625 12978 7630
rect 13230 7658 13258 7663
rect 13230 7611 13258 7630
rect 13398 7658 13426 7663
rect 13398 7611 13426 7630
rect 13510 7657 13538 8358
rect 13510 7631 13511 7657
rect 13537 7631 13538 7657
rect 13510 7625 13538 7631
rect 13902 7658 13930 8414
rect 14406 7713 14434 8526
rect 15078 8498 15106 8695
rect 15134 8666 15162 8807
rect 15302 8833 15330 9366
rect 15470 9169 15498 9478
rect 15470 9143 15471 9169
rect 15497 9143 15498 9169
rect 15470 9137 15498 9143
rect 15526 9282 15554 9287
rect 15526 9170 15554 9254
rect 15694 9170 15722 10710
rect 18830 10738 18858 11159
rect 20006 10794 20034 11215
rect 20006 10761 20034 10766
rect 18830 10705 18858 10710
rect 17598 10598 17730 10603
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17598 10565 17730 10570
rect 20006 10457 20034 10463
rect 20006 10431 20007 10457
rect 20033 10431 20034 10457
rect 18830 10401 18858 10407
rect 18830 10375 18831 10401
rect 18857 10375 18858 10401
rect 17598 9814 17730 9819
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17598 9781 17730 9786
rect 18830 9506 18858 10375
rect 20006 10122 20034 10431
rect 20006 10089 20034 10094
rect 18830 9473 18858 9478
rect 15526 9169 15722 9170
rect 15526 9143 15695 9169
rect 15721 9143 15722 9169
rect 15526 9142 15722 9143
rect 15302 8807 15303 8833
rect 15329 8807 15330 8833
rect 15302 8801 15330 8807
rect 15470 8890 15498 8895
rect 15134 8633 15162 8638
rect 15246 8778 15274 8783
rect 15078 8465 15106 8470
rect 15246 8442 15274 8750
rect 15246 8386 15274 8414
rect 15302 8386 15330 8391
rect 15246 8385 15330 8386
rect 15246 8359 15303 8385
rect 15329 8359 15330 8385
rect 15246 8358 15330 8359
rect 15302 8353 15330 8358
rect 14406 7687 14407 7713
rect 14433 7687 14434 7713
rect 14406 7681 14434 7687
rect 14014 7658 14042 7663
rect 13902 7657 14042 7658
rect 13902 7631 14015 7657
rect 14041 7631 14042 7657
rect 13902 7630 14042 7631
rect 13062 7601 13090 7607
rect 13062 7575 13063 7601
rect 13089 7575 13090 7601
rect 13062 7154 13090 7575
rect 13062 7121 13090 7126
rect 13342 7321 13370 7327
rect 13342 7295 13343 7321
rect 13369 7295 13370 7321
rect 13342 6986 13370 7295
rect 12726 6939 12754 6958
rect 13062 6958 13370 6986
rect 13454 7154 13482 7159
rect 12558 6930 12586 6935
rect 12558 6873 12586 6902
rect 12558 6847 12559 6873
rect 12585 6847 12586 6873
rect 12558 6841 12586 6847
rect 12838 6930 12866 6935
rect 13062 6930 13090 6958
rect 12838 6929 13090 6930
rect 12838 6903 12839 6929
rect 12865 6903 13090 6929
rect 12838 6902 13090 6903
rect 13454 6929 13482 7126
rect 13454 6903 13455 6929
rect 13481 6903 13482 6929
rect 12334 6785 12362 6790
rect 12670 6818 12698 6823
rect 12670 6771 12698 6790
rect 12782 6706 12810 6711
rect 12558 6538 12586 6543
rect 12278 6537 12586 6538
rect 12278 6511 12559 6537
rect 12585 6511 12586 6537
rect 12278 6510 12586 6511
rect 11942 6175 11943 6201
rect 11969 6175 11970 6201
rect 11942 6169 11970 6175
rect 12558 5866 12586 6510
rect 12782 6537 12810 6678
rect 12782 6511 12783 6537
rect 12809 6511 12810 6537
rect 12782 6505 12810 6511
rect 12558 5838 12642 5866
rect 8414 4186 8554 4214
rect 10654 4186 10850 4214
rect 11774 4186 12306 4214
rect 2238 3542 2370 3547
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2238 3509 2370 3514
rect 2238 2758 2370 2763
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2238 2725 2370 2730
rect 2238 1974 2370 1979
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2238 1941 2370 1946
rect 8526 1777 8554 4186
rect 9918 3934 10050 3939
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 9918 3901 10050 3906
rect 9918 3150 10050 3155
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 9918 3117 10050 3122
rect 9918 2366 10050 2371
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 9918 2333 10050 2338
rect 8526 1751 8527 1777
rect 8553 1751 8554 1777
rect 8526 1745 8554 1751
rect 10766 1834 10794 1839
rect 8414 1722 8442 1727
rect 8414 400 8442 1694
rect 9030 1722 9058 1727
rect 9030 1665 9058 1694
rect 9030 1639 9031 1665
rect 9057 1639 9058 1665
rect 9030 1633 9058 1639
rect 9918 1582 10050 1587
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 9918 1549 10050 1554
rect 10766 400 10794 1806
rect 10822 1777 10850 4186
rect 11214 1834 11242 1839
rect 11214 1787 11242 1806
rect 11774 1834 11802 1839
rect 10822 1751 10823 1777
rect 10849 1751 10850 1777
rect 10822 1745 10850 1751
rect 11774 400 11802 1806
rect 12278 1777 12306 4186
rect 12614 2169 12642 5838
rect 12838 4214 12866 6902
rect 13454 6897 13482 6903
rect 13566 7154 13594 7159
rect 13118 6873 13146 6879
rect 13118 6847 13119 6873
rect 13145 6847 13146 6873
rect 13062 6762 13090 6767
rect 13118 6762 13146 6847
rect 13090 6734 13146 6762
rect 13566 6762 13594 7126
rect 14014 7154 14042 7630
rect 14014 7121 14042 7126
rect 14518 7658 14546 7663
rect 14518 6817 14546 7630
rect 15470 7601 15498 8862
rect 15526 8554 15554 9142
rect 15694 9137 15722 9142
rect 17598 9030 17730 9035
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17598 8997 17730 9002
rect 20006 8889 20034 8895
rect 20006 8863 20007 8889
rect 20033 8863 20034 8889
rect 18830 8834 18858 8839
rect 18830 8787 18858 8806
rect 20006 8778 20034 8863
rect 20006 8745 20034 8750
rect 15526 8553 15722 8554
rect 15526 8527 15527 8553
rect 15553 8527 15722 8553
rect 15526 8526 15722 8527
rect 15526 8521 15554 8526
rect 15694 7769 15722 8526
rect 18830 8442 18858 8447
rect 18830 8395 18858 8414
rect 20006 8442 20034 8447
rect 20006 8385 20034 8414
rect 20006 8359 20007 8385
rect 20033 8359 20034 8385
rect 20006 8353 20034 8359
rect 17598 8246 17730 8251
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17598 8213 17730 8218
rect 15694 7743 15695 7769
rect 15721 7743 15722 7769
rect 15694 7737 15722 7743
rect 18830 7658 18858 7663
rect 18830 7611 18858 7630
rect 15470 7575 15471 7601
rect 15497 7575 15498 7601
rect 15470 7569 15498 7575
rect 20006 7601 20034 7607
rect 20006 7575 20007 7601
rect 20033 7575 20034 7601
rect 17598 7462 17730 7467
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17598 7429 17730 7434
rect 20006 7434 20034 7575
rect 20006 7401 20034 7406
rect 14742 7154 14770 7159
rect 14742 6985 14770 7126
rect 14742 6959 14743 6985
rect 14769 6959 14770 6985
rect 14742 6953 14770 6959
rect 14518 6791 14519 6817
rect 14545 6791 14546 6817
rect 14518 6785 14546 6791
rect 13062 6729 13090 6734
rect 13566 6729 13594 6734
rect 17598 6678 17730 6683
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17598 6645 17730 6650
rect 17598 5894 17730 5899
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17598 5861 17730 5866
rect 17598 5110 17730 5115
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17598 5077 17730 5082
rect 17598 4326 17730 4331
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17598 4293 17730 4298
rect 12838 4186 12922 4214
rect 12614 2143 12615 2169
rect 12641 2143 12642 2169
rect 12614 2137 12642 2143
rect 12838 2618 12866 2623
rect 12278 1751 12279 1777
rect 12305 1751 12306 1777
rect 12278 1745 12306 1751
rect 12446 2058 12474 2063
rect 12446 400 12474 2030
rect 12782 1834 12810 1839
rect 12782 1787 12810 1806
rect 12838 1218 12866 2590
rect 12894 2561 12922 4186
rect 17598 3542 17730 3547
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17598 3509 17730 3514
rect 17598 2758 17730 2763
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17598 2725 17730 2730
rect 13398 2618 13426 2623
rect 13398 2571 13426 2590
rect 12894 2535 12895 2561
rect 12921 2535 12922 2561
rect 12894 2529 12922 2535
rect 13118 2058 13146 2063
rect 13118 2011 13146 2030
rect 17598 1974 17730 1979
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17598 1941 17730 1946
rect 12782 1190 12866 1218
rect 12782 400 12810 1190
rect 8400 0 8456 400
rect 10752 0 10808 400
rect 11760 0 11816 400
rect 12432 0 12488 400
rect 12768 0 12824 400
<< via2 >>
rect 2238 19221 2266 19222
rect 2238 19195 2239 19221
rect 2239 19195 2265 19221
rect 2265 19195 2266 19221
rect 2238 19194 2266 19195
rect 2290 19221 2318 19222
rect 2290 19195 2291 19221
rect 2291 19195 2317 19221
rect 2317 19195 2318 19221
rect 2290 19194 2318 19195
rect 2342 19221 2370 19222
rect 2342 19195 2343 19221
rect 2343 19195 2369 19221
rect 2369 19195 2370 19221
rect 2342 19194 2370 19195
rect 2238 18437 2266 18438
rect 2238 18411 2239 18437
rect 2239 18411 2265 18437
rect 2265 18411 2266 18437
rect 2238 18410 2266 18411
rect 2290 18437 2318 18438
rect 2290 18411 2291 18437
rect 2291 18411 2317 18437
rect 2317 18411 2318 18437
rect 2290 18410 2318 18411
rect 2342 18437 2370 18438
rect 2342 18411 2343 18437
rect 2343 18411 2369 18437
rect 2369 18411 2370 18437
rect 2342 18410 2370 18411
rect 8078 19110 8106 19138
rect 8974 19137 9002 19138
rect 8974 19111 8975 19137
rect 8975 19111 9001 19137
rect 9001 19111 9002 19137
rect 8974 19110 9002 19111
rect 7742 18326 7770 18354
rect 8358 18353 8386 18354
rect 8358 18327 8359 18353
rect 8359 18327 8385 18353
rect 8385 18327 8386 18353
rect 8358 18326 8386 18327
rect 2238 17653 2266 17654
rect 2238 17627 2239 17653
rect 2239 17627 2265 17653
rect 2265 17627 2266 17653
rect 2238 17626 2266 17627
rect 2290 17653 2318 17654
rect 2290 17627 2291 17653
rect 2291 17627 2317 17653
rect 2317 17627 2318 17653
rect 2290 17626 2318 17627
rect 2342 17653 2370 17654
rect 2342 17627 2343 17653
rect 2343 17627 2369 17653
rect 2369 17627 2370 17653
rect 2342 17626 2370 17627
rect 2238 16869 2266 16870
rect 2238 16843 2239 16869
rect 2239 16843 2265 16869
rect 2265 16843 2266 16869
rect 2238 16842 2266 16843
rect 2290 16869 2318 16870
rect 2290 16843 2291 16869
rect 2291 16843 2317 16869
rect 2317 16843 2318 16869
rect 2290 16842 2318 16843
rect 2342 16869 2370 16870
rect 2342 16843 2343 16869
rect 2343 16843 2369 16869
rect 2369 16843 2370 16869
rect 2342 16842 2370 16843
rect 2238 16085 2266 16086
rect 2238 16059 2239 16085
rect 2239 16059 2265 16085
rect 2265 16059 2266 16085
rect 2238 16058 2266 16059
rect 2290 16085 2318 16086
rect 2290 16059 2291 16085
rect 2291 16059 2317 16085
rect 2317 16059 2318 16085
rect 2290 16058 2318 16059
rect 2342 16085 2370 16086
rect 2342 16059 2343 16085
rect 2343 16059 2369 16085
rect 2369 16059 2370 16085
rect 2342 16058 2370 16059
rect 2238 15301 2266 15302
rect 2238 15275 2239 15301
rect 2239 15275 2265 15301
rect 2265 15275 2266 15301
rect 2238 15274 2266 15275
rect 2290 15301 2318 15302
rect 2290 15275 2291 15301
rect 2291 15275 2317 15301
rect 2317 15275 2318 15301
rect 2290 15274 2318 15275
rect 2342 15301 2370 15302
rect 2342 15275 2343 15301
rect 2343 15275 2369 15301
rect 2369 15275 2370 15301
rect 2342 15274 2370 15275
rect 2238 14517 2266 14518
rect 2238 14491 2239 14517
rect 2239 14491 2265 14517
rect 2265 14491 2266 14517
rect 2238 14490 2266 14491
rect 2290 14517 2318 14518
rect 2290 14491 2291 14517
rect 2291 14491 2317 14517
rect 2317 14491 2318 14517
rect 2290 14490 2318 14491
rect 2342 14517 2370 14518
rect 2342 14491 2343 14517
rect 2343 14491 2369 14517
rect 2369 14491 2370 14517
rect 2342 14490 2370 14491
rect 10430 19110 10458 19138
rect 11046 19137 11074 19138
rect 11046 19111 11047 19137
rect 11047 19111 11073 19137
rect 11073 19111 11074 19137
rect 11046 19110 11074 19111
rect 12110 19110 12138 19138
rect 12782 19137 12810 19138
rect 12782 19111 12783 19137
rect 12783 19111 12809 19137
rect 12809 19111 12810 19137
rect 12782 19110 12810 19111
rect 9918 18829 9946 18830
rect 9918 18803 9919 18829
rect 9919 18803 9945 18829
rect 9945 18803 9946 18829
rect 9918 18802 9946 18803
rect 9970 18829 9998 18830
rect 9970 18803 9971 18829
rect 9971 18803 9997 18829
rect 9997 18803 9998 18829
rect 9970 18802 9998 18803
rect 10022 18829 10050 18830
rect 10022 18803 10023 18829
rect 10023 18803 10049 18829
rect 10049 18803 10050 18829
rect 10022 18802 10050 18803
rect 9422 18718 9450 18746
rect 10038 18745 10066 18746
rect 10038 18719 10039 18745
rect 10039 18719 10065 18745
rect 10065 18719 10066 18745
rect 10038 18718 10066 18719
rect 6678 13929 6706 13930
rect 6678 13903 6679 13929
rect 6679 13903 6705 13929
rect 6705 13903 6706 13929
rect 6678 13902 6706 13903
rect 2238 13733 2266 13734
rect 2238 13707 2239 13733
rect 2239 13707 2265 13733
rect 2265 13707 2266 13733
rect 2238 13706 2266 13707
rect 2290 13733 2318 13734
rect 2290 13707 2291 13733
rect 2291 13707 2317 13733
rect 2317 13707 2318 13733
rect 2290 13706 2318 13707
rect 2342 13733 2370 13734
rect 2342 13707 2343 13733
rect 2343 13707 2369 13733
rect 2369 13707 2370 13733
rect 2342 13706 2370 13707
rect 2086 13454 2114 13482
rect 966 12446 994 12474
rect 966 12249 994 12250
rect 966 12223 967 12249
rect 967 12223 993 12249
rect 993 12223 994 12249
rect 966 12222 994 12223
rect 966 11774 994 11802
rect 2030 11494 2058 11522
rect 966 11465 994 11466
rect 966 11439 967 11465
rect 967 11439 993 11465
rect 993 11439 994 11465
rect 966 11438 994 11439
rect 966 10430 994 10458
rect 2238 12949 2266 12950
rect 2238 12923 2239 12949
rect 2239 12923 2265 12949
rect 2265 12923 2266 12949
rect 2238 12922 2266 12923
rect 2290 12949 2318 12950
rect 2290 12923 2291 12949
rect 2291 12923 2317 12949
rect 2317 12923 2318 12949
rect 2290 12922 2318 12923
rect 2342 12949 2370 12950
rect 2342 12923 2343 12949
rect 2343 12923 2369 12949
rect 2369 12923 2370 12949
rect 2342 12922 2370 12923
rect 2142 12753 2170 12754
rect 2142 12727 2143 12753
rect 2143 12727 2169 12753
rect 2169 12727 2170 12753
rect 2142 12726 2170 12727
rect 6734 12726 6762 12754
rect 7294 12670 7322 12698
rect 2142 12361 2170 12362
rect 2142 12335 2143 12361
rect 2143 12335 2169 12361
rect 2169 12335 2170 12361
rect 2142 12334 2170 12335
rect 6902 12334 6930 12362
rect 2238 12165 2266 12166
rect 2238 12139 2239 12165
rect 2239 12139 2265 12165
rect 2265 12139 2266 12165
rect 2238 12138 2266 12139
rect 2290 12165 2318 12166
rect 2290 12139 2291 12165
rect 2291 12139 2317 12165
rect 2317 12139 2318 12165
rect 2290 12138 2318 12139
rect 2342 12165 2370 12166
rect 2342 12139 2343 12165
rect 2343 12139 2369 12165
rect 2369 12139 2370 12165
rect 2342 12138 2370 12139
rect 7126 12222 7154 12250
rect 2142 11718 2170 11746
rect 7014 11606 7042 11634
rect 6902 11577 6930 11578
rect 6902 11551 6903 11577
rect 6903 11551 6929 11577
rect 6929 11551 6930 11577
rect 6902 11550 6930 11551
rect 5502 11521 5530 11522
rect 5502 11495 5503 11521
rect 5503 11495 5529 11521
rect 5529 11495 5530 11521
rect 5502 11494 5530 11495
rect 6566 11521 6594 11522
rect 6566 11495 6567 11521
rect 6567 11495 6593 11521
rect 6593 11495 6594 11521
rect 6566 11494 6594 11495
rect 2238 11381 2266 11382
rect 2238 11355 2239 11381
rect 2239 11355 2265 11381
rect 2265 11355 2266 11381
rect 2238 11354 2266 11355
rect 2290 11381 2318 11382
rect 2290 11355 2291 11381
rect 2291 11355 2317 11381
rect 2317 11355 2318 11381
rect 2290 11354 2318 11355
rect 2342 11381 2370 11382
rect 2342 11355 2343 11381
rect 2343 11355 2369 11381
rect 2369 11355 2370 11381
rect 2342 11354 2370 11355
rect 7126 11438 7154 11466
rect 2142 10793 2170 10794
rect 2142 10767 2143 10793
rect 2143 10767 2169 10793
rect 2169 10767 2170 10793
rect 2142 10766 2170 10767
rect 4998 10766 5026 10794
rect 2238 10597 2266 10598
rect 2238 10571 2239 10597
rect 2239 10571 2265 10597
rect 2265 10571 2266 10597
rect 2238 10570 2266 10571
rect 2290 10597 2318 10598
rect 2290 10571 2291 10597
rect 2291 10571 2317 10597
rect 2317 10571 2318 10597
rect 2290 10570 2318 10571
rect 2342 10597 2370 10598
rect 2342 10571 2343 10597
rect 2343 10571 2369 10597
rect 2369 10571 2370 10597
rect 2342 10570 2370 10571
rect 2086 10374 2114 10402
rect 4998 10318 5026 10346
rect 2142 10009 2170 10010
rect 2142 9983 2143 10009
rect 2143 9983 2169 10009
rect 2169 9983 2170 10009
rect 2142 9982 2170 9983
rect 4942 9982 4970 10010
rect 966 9897 994 9898
rect 966 9871 967 9897
rect 967 9871 993 9897
rect 993 9871 994 9897
rect 966 9870 994 9871
rect 2238 9813 2266 9814
rect 2238 9787 2239 9813
rect 2239 9787 2265 9813
rect 2265 9787 2266 9813
rect 2238 9786 2266 9787
rect 2290 9813 2318 9814
rect 2290 9787 2291 9813
rect 2291 9787 2317 9813
rect 2317 9787 2318 9813
rect 2290 9786 2318 9787
rect 2342 9813 2370 9814
rect 2342 9787 2343 9813
rect 2343 9787 2369 9813
rect 2369 9787 2370 9813
rect 2342 9786 2370 9787
rect 6230 10262 6258 10290
rect 4942 9590 4970 9618
rect 6846 10598 6874 10626
rect 7350 12278 7378 12306
rect 8134 13902 8162 13930
rect 8750 13902 8778 13930
rect 7966 13481 7994 13482
rect 7966 13455 7967 13481
rect 7967 13455 7993 13481
rect 7993 13455 7994 13481
rect 7966 13454 7994 13455
rect 7742 13033 7770 13034
rect 7742 13007 7743 13033
rect 7743 13007 7769 13033
rect 7769 13007 7770 13033
rect 7742 13006 7770 13007
rect 7630 12726 7658 12754
rect 8470 13454 8498 13482
rect 8358 13006 8386 13034
rect 8358 12753 8386 12754
rect 8358 12727 8359 12753
rect 8359 12727 8385 12753
rect 8385 12727 8386 12753
rect 8358 12726 8386 12727
rect 7798 12697 7826 12698
rect 7798 12671 7799 12697
rect 7799 12671 7825 12697
rect 7825 12671 7826 12697
rect 7798 12670 7826 12671
rect 8526 13230 8554 13258
rect 8974 13929 9002 13930
rect 8974 13903 8975 13929
rect 8975 13903 9001 13929
rect 9001 13903 9002 13929
rect 8974 13902 9002 13903
rect 9086 13454 9114 13482
rect 9918 18045 9946 18046
rect 9918 18019 9919 18045
rect 9919 18019 9945 18045
rect 9945 18019 9946 18045
rect 9918 18018 9946 18019
rect 9970 18045 9998 18046
rect 9970 18019 9971 18045
rect 9971 18019 9997 18045
rect 9997 18019 9998 18045
rect 9970 18018 9998 18019
rect 10022 18045 10050 18046
rect 10022 18019 10023 18045
rect 10023 18019 10049 18045
rect 10049 18019 10050 18045
rect 10022 18018 10050 18019
rect 9918 17261 9946 17262
rect 9918 17235 9919 17261
rect 9919 17235 9945 17261
rect 9945 17235 9946 17261
rect 9918 17234 9946 17235
rect 9970 17261 9998 17262
rect 9970 17235 9971 17261
rect 9971 17235 9997 17261
rect 9997 17235 9998 17261
rect 9970 17234 9998 17235
rect 10022 17261 10050 17262
rect 10022 17235 10023 17261
rect 10023 17235 10049 17261
rect 10049 17235 10050 17261
rect 10022 17234 10050 17235
rect 9918 16477 9946 16478
rect 9918 16451 9919 16477
rect 9919 16451 9945 16477
rect 9945 16451 9946 16477
rect 9918 16450 9946 16451
rect 9970 16477 9998 16478
rect 9970 16451 9971 16477
rect 9971 16451 9997 16477
rect 9997 16451 9998 16477
rect 9970 16450 9998 16451
rect 10022 16477 10050 16478
rect 10022 16451 10023 16477
rect 10023 16451 10049 16477
rect 10049 16451 10050 16477
rect 10022 16450 10050 16451
rect 17598 19221 17626 19222
rect 17598 19195 17599 19221
rect 17599 19195 17625 19221
rect 17625 19195 17626 19221
rect 17598 19194 17626 19195
rect 17650 19221 17678 19222
rect 17650 19195 17651 19221
rect 17651 19195 17677 19221
rect 17677 19195 17678 19221
rect 17650 19194 17678 19195
rect 17702 19221 17730 19222
rect 17702 19195 17703 19221
rect 17703 19195 17729 19221
rect 17729 19195 17730 19221
rect 17702 19194 17730 19195
rect 13118 18718 13146 18746
rect 13734 18745 13762 18746
rect 13734 18719 13735 18745
rect 13735 18719 13761 18745
rect 13761 18719 13762 18745
rect 13734 18718 13762 18719
rect 17598 18437 17626 18438
rect 17598 18411 17599 18437
rect 17599 18411 17625 18437
rect 17625 18411 17626 18437
rect 17598 18410 17626 18411
rect 17650 18437 17678 18438
rect 17650 18411 17651 18437
rect 17651 18411 17677 18437
rect 17677 18411 17678 18437
rect 17650 18410 17678 18411
rect 17702 18437 17730 18438
rect 17702 18411 17703 18437
rect 17703 18411 17729 18437
rect 17729 18411 17730 18437
rect 17702 18410 17730 18411
rect 17598 17653 17626 17654
rect 17598 17627 17599 17653
rect 17599 17627 17625 17653
rect 17625 17627 17626 17653
rect 17598 17626 17626 17627
rect 17650 17653 17678 17654
rect 17650 17627 17651 17653
rect 17651 17627 17677 17653
rect 17677 17627 17678 17653
rect 17650 17626 17678 17627
rect 17702 17653 17730 17654
rect 17702 17627 17703 17653
rect 17703 17627 17729 17653
rect 17729 17627 17730 17653
rect 17702 17626 17730 17627
rect 17598 16869 17626 16870
rect 17598 16843 17599 16869
rect 17599 16843 17625 16869
rect 17625 16843 17626 16869
rect 17598 16842 17626 16843
rect 17650 16869 17678 16870
rect 17650 16843 17651 16869
rect 17651 16843 17677 16869
rect 17677 16843 17678 16869
rect 17650 16842 17678 16843
rect 17702 16869 17730 16870
rect 17702 16843 17703 16869
rect 17703 16843 17729 16869
rect 17729 16843 17730 16869
rect 17702 16842 17730 16843
rect 17598 16085 17626 16086
rect 17598 16059 17599 16085
rect 17599 16059 17625 16085
rect 17625 16059 17626 16085
rect 17598 16058 17626 16059
rect 17650 16085 17678 16086
rect 17650 16059 17651 16085
rect 17651 16059 17677 16085
rect 17677 16059 17678 16085
rect 17650 16058 17678 16059
rect 17702 16085 17730 16086
rect 17702 16059 17703 16085
rect 17703 16059 17729 16085
rect 17729 16059 17730 16085
rect 17702 16058 17730 16059
rect 9918 15693 9946 15694
rect 9918 15667 9919 15693
rect 9919 15667 9945 15693
rect 9945 15667 9946 15693
rect 9918 15666 9946 15667
rect 9970 15693 9998 15694
rect 9970 15667 9971 15693
rect 9971 15667 9997 15693
rect 9997 15667 9998 15693
rect 9970 15666 9998 15667
rect 10022 15693 10050 15694
rect 10022 15667 10023 15693
rect 10023 15667 10049 15693
rect 10049 15667 10050 15693
rect 10022 15666 10050 15667
rect 9918 14909 9946 14910
rect 9918 14883 9919 14909
rect 9919 14883 9945 14909
rect 9945 14883 9946 14909
rect 9918 14882 9946 14883
rect 9970 14909 9998 14910
rect 9970 14883 9971 14909
rect 9971 14883 9997 14909
rect 9997 14883 9998 14909
rect 9970 14882 9998 14883
rect 10022 14909 10050 14910
rect 10022 14883 10023 14909
rect 10023 14883 10049 14909
rect 10049 14883 10050 14909
rect 10022 14882 10050 14883
rect 9918 14125 9946 14126
rect 9918 14099 9919 14125
rect 9919 14099 9945 14125
rect 9945 14099 9946 14125
rect 9918 14098 9946 14099
rect 9970 14125 9998 14126
rect 9970 14099 9971 14125
rect 9971 14099 9997 14125
rect 9997 14099 9998 14125
rect 9970 14098 9998 14099
rect 10022 14125 10050 14126
rect 10022 14099 10023 14125
rect 10023 14099 10049 14125
rect 10049 14099 10050 14125
rect 10022 14098 10050 14099
rect 10262 13846 10290 13874
rect 8974 13257 9002 13258
rect 8974 13231 8975 13257
rect 8975 13231 9001 13257
rect 9001 13231 9002 13257
rect 8974 13230 9002 13231
rect 8750 12641 8778 12642
rect 8750 12615 8751 12641
rect 8751 12615 8777 12641
rect 8777 12615 8778 12641
rect 8750 12614 8778 12615
rect 7462 12222 7490 12250
rect 9030 13145 9058 13146
rect 9030 13119 9031 13145
rect 9031 13119 9057 13145
rect 9057 13119 9058 13145
rect 9030 13118 9058 13119
rect 7238 11633 7266 11634
rect 7238 11607 7239 11633
rect 7239 11607 7265 11633
rect 7265 11607 7266 11633
rect 7238 11606 7266 11607
rect 7350 11633 7378 11634
rect 7350 11607 7351 11633
rect 7351 11607 7377 11633
rect 7377 11607 7378 11633
rect 7350 11606 7378 11607
rect 7686 11633 7714 11634
rect 7686 11607 7687 11633
rect 7687 11607 7713 11633
rect 7713 11607 7714 11633
rect 7686 11606 7714 11607
rect 7294 11550 7322 11578
rect 6958 10486 6986 10514
rect 6846 10345 6874 10346
rect 6846 10319 6847 10345
rect 6847 10319 6873 10345
rect 6873 10319 6874 10345
rect 6846 10318 6874 10319
rect 6790 10289 6818 10290
rect 6790 10263 6791 10289
rect 6791 10263 6817 10289
rect 6817 10263 6818 10289
rect 6790 10262 6818 10263
rect 7014 10542 7042 10570
rect 7630 11521 7658 11522
rect 7630 11495 7631 11521
rect 7631 11495 7657 11521
rect 7657 11495 7658 11521
rect 7630 11494 7658 11495
rect 7574 11465 7602 11466
rect 7574 11439 7575 11465
rect 7575 11439 7601 11465
rect 7601 11439 7602 11465
rect 7574 11438 7602 11439
rect 7686 11438 7714 11466
rect 7462 11102 7490 11130
rect 8526 10542 8554 10570
rect 8470 10513 8498 10514
rect 8470 10487 8471 10513
rect 8471 10487 8497 10513
rect 8497 10487 8498 10513
rect 8470 10486 8498 10487
rect 7182 10262 7210 10290
rect 6734 9617 6762 9618
rect 6734 9591 6735 9617
rect 6735 9591 6761 9617
rect 6761 9591 6762 9617
rect 6734 9590 6762 9591
rect 6398 9478 6426 9506
rect 6678 9478 6706 9506
rect 6230 9310 6258 9338
rect 6342 9254 6370 9282
rect 2238 9029 2266 9030
rect 2238 9003 2239 9029
rect 2239 9003 2265 9029
rect 2265 9003 2266 9029
rect 2238 9002 2266 9003
rect 2290 9029 2318 9030
rect 2290 9003 2291 9029
rect 2291 9003 2317 9029
rect 2317 9003 2318 9029
rect 2290 9002 2318 9003
rect 2342 9029 2370 9030
rect 2342 9003 2343 9029
rect 2343 9003 2369 9029
rect 2369 9003 2370 9029
rect 2342 9002 2370 9003
rect 6454 9225 6482 9226
rect 6454 9199 6455 9225
rect 6455 9199 6481 9225
rect 6481 9199 6482 9225
rect 6454 9198 6482 9199
rect 6846 9254 6874 9282
rect 6398 8862 6426 8890
rect 2142 8833 2170 8834
rect 2142 8807 2143 8833
rect 2143 8807 2169 8833
rect 2169 8807 2170 8833
rect 2142 8806 2170 8807
rect 5558 8806 5586 8834
rect 966 8414 994 8442
rect 7126 9198 7154 9226
rect 9030 12726 9058 12754
rect 9366 13145 9394 13146
rect 9366 13119 9367 13145
rect 9367 13119 9393 13145
rect 9393 13119 9394 13145
rect 9366 13118 9394 13119
rect 9870 13790 9898 13818
rect 10654 13873 10682 13874
rect 10654 13847 10655 13873
rect 10655 13847 10681 13873
rect 10681 13847 10682 13873
rect 10654 13846 10682 13847
rect 10430 13790 10458 13818
rect 12054 13790 12082 13818
rect 9758 13481 9786 13482
rect 9758 13455 9759 13481
rect 9759 13455 9785 13481
rect 9785 13455 9786 13481
rect 9758 13454 9786 13455
rect 9534 13398 9562 13426
rect 9422 13006 9450 13034
rect 9870 13398 9898 13426
rect 9918 13341 9946 13342
rect 9918 13315 9919 13341
rect 9919 13315 9945 13341
rect 9945 13315 9946 13341
rect 9918 13314 9946 13315
rect 9970 13341 9998 13342
rect 9970 13315 9971 13341
rect 9971 13315 9997 13341
rect 9997 13315 9998 13341
rect 9970 13314 9998 13315
rect 10022 13341 10050 13342
rect 10022 13315 10023 13341
rect 10023 13315 10049 13341
rect 10049 13315 10050 13341
rect 10022 13314 10050 13315
rect 9758 13033 9786 13034
rect 9758 13007 9759 13033
rect 9759 13007 9785 13033
rect 9785 13007 9786 13033
rect 9758 13006 9786 13007
rect 9142 11886 9170 11914
rect 8974 11494 9002 11522
rect 8862 11382 8890 11410
rect 9142 11438 9170 11466
rect 9142 11102 9170 11130
rect 8974 10486 9002 10514
rect 9254 11689 9282 11690
rect 9254 11663 9255 11689
rect 9255 11663 9281 11689
rect 9281 11663 9282 11689
rect 9254 11662 9282 11663
rect 9478 11606 9506 11634
rect 9534 12558 9562 12586
rect 9534 12278 9562 12306
rect 9918 12557 9946 12558
rect 9918 12531 9919 12557
rect 9919 12531 9945 12557
rect 9945 12531 9946 12557
rect 9918 12530 9946 12531
rect 9970 12557 9998 12558
rect 9970 12531 9971 12557
rect 9971 12531 9997 12557
rect 9997 12531 9998 12557
rect 9970 12530 9998 12531
rect 10022 12557 10050 12558
rect 10022 12531 10023 12557
rect 10023 12531 10049 12557
rect 10049 12531 10050 12557
rect 10022 12530 10050 12531
rect 10374 12614 10402 12642
rect 9590 12334 9618 12362
rect 9590 11969 9618 11970
rect 9590 11943 9591 11969
rect 9591 11943 9617 11969
rect 9617 11943 9618 11969
rect 9590 11942 9618 11943
rect 9702 11913 9730 11914
rect 9702 11887 9703 11913
rect 9703 11887 9729 11913
rect 9729 11887 9730 11913
rect 9702 11886 9730 11887
rect 10822 13145 10850 13146
rect 10822 13119 10823 13145
rect 10823 13119 10849 13145
rect 10849 13119 10850 13145
rect 10822 13118 10850 13119
rect 9310 11382 9338 11410
rect 9366 11102 9394 11130
rect 9198 10318 9226 10346
rect 9254 10262 9282 10290
rect 8862 10065 8890 10066
rect 8862 10039 8863 10065
rect 8863 10039 8889 10065
rect 8889 10039 8890 10065
rect 8862 10038 8890 10039
rect 8414 9982 8442 10010
rect 8246 9534 8274 9562
rect 8358 9505 8386 9506
rect 8358 9479 8359 9505
rect 8359 9479 8385 9505
rect 8385 9479 8386 9505
rect 8358 9478 8386 9479
rect 7742 9225 7770 9226
rect 7742 9199 7743 9225
rect 7743 9199 7769 9225
rect 7769 9199 7770 9225
rect 7742 9198 7770 9199
rect 6958 8889 6986 8890
rect 6958 8863 6959 8889
rect 6959 8863 6985 8889
rect 6985 8863 6986 8889
rect 6958 8862 6986 8863
rect 7126 8862 7154 8890
rect 6902 8806 6930 8834
rect 7742 8862 7770 8890
rect 7462 8833 7490 8834
rect 7462 8807 7463 8833
rect 7463 8807 7489 8833
rect 7489 8807 7490 8833
rect 7462 8806 7490 8807
rect 7014 8777 7042 8778
rect 7014 8751 7015 8777
rect 7015 8751 7041 8777
rect 7041 8751 7042 8777
rect 7014 8750 7042 8751
rect 7238 8777 7266 8778
rect 7238 8751 7239 8777
rect 7239 8751 7265 8777
rect 7265 8751 7266 8777
rect 7238 8750 7266 8751
rect 7742 8750 7770 8778
rect 7798 8974 7826 9002
rect 7630 8694 7658 8722
rect 7462 8497 7490 8498
rect 7462 8471 7463 8497
rect 7463 8471 7489 8497
rect 7489 8471 7490 8497
rect 7462 8470 7490 8471
rect 2238 8245 2266 8246
rect 2238 8219 2239 8245
rect 2239 8219 2265 8245
rect 2265 8219 2266 8245
rect 2238 8218 2266 8219
rect 2290 8245 2318 8246
rect 2290 8219 2291 8245
rect 2291 8219 2317 8245
rect 2317 8219 2318 8245
rect 2290 8218 2318 8219
rect 2342 8245 2370 8246
rect 2342 8219 2343 8245
rect 2343 8219 2369 8245
rect 2369 8219 2370 8245
rect 2342 8218 2370 8219
rect 6846 7574 6874 7602
rect 7518 8414 7546 8442
rect 8022 9030 8050 9058
rect 8134 8750 8162 8778
rect 8190 8470 8218 8498
rect 7014 7574 7042 7602
rect 8302 8441 8330 8442
rect 8302 8415 8303 8441
rect 8303 8415 8329 8441
rect 8329 8415 8330 8441
rect 8302 8414 8330 8415
rect 8246 8385 8274 8386
rect 8246 8359 8247 8385
rect 8247 8359 8273 8385
rect 8273 8359 8274 8385
rect 8246 8358 8274 8359
rect 8414 9113 8442 9114
rect 8414 9087 8415 9113
rect 8415 9087 8441 9113
rect 8441 9087 8442 9113
rect 8414 9086 8442 9087
rect 8918 9870 8946 9898
rect 8862 9590 8890 9618
rect 8750 9310 8778 9338
rect 8638 9225 8666 9226
rect 8638 9199 8639 9225
rect 8639 9199 8665 9225
rect 8665 9199 8666 9225
rect 8638 9198 8666 9199
rect 8862 9422 8890 9450
rect 8470 8974 8498 9002
rect 8414 8889 8442 8890
rect 8414 8863 8415 8889
rect 8415 8863 8441 8889
rect 8441 8863 8442 8889
rect 8414 8862 8442 8863
rect 9198 9926 9226 9954
rect 8918 9086 8946 9114
rect 8414 8694 8442 8722
rect 8694 8721 8722 8722
rect 8694 8695 8695 8721
rect 8695 8695 8721 8721
rect 8721 8695 8722 8721
rect 8694 8694 8722 8695
rect 8974 8974 9002 9002
rect 8414 7601 8442 7602
rect 8414 7575 8415 7601
rect 8415 7575 8441 7601
rect 8441 7575 8442 7601
rect 8414 7574 8442 7575
rect 2238 7461 2266 7462
rect 2238 7435 2239 7461
rect 2239 7435 2265 7461
rect 2265 7435 2266 7461
rect 2238 7434 2266 7435
rect 2290 7461 2318 7462
rect 2290 7435 2291 7461
rect 2291 7435 2317 7461
rect 2317 7435 2318 7461
rect 2290 7434 2318 7435
rect 2342 7461 2370 7462
rect 2342 7435 2343 7461
rect 2343 7435 2369 7461
rect 2369 7435 2370 7461
rect 2342 7434 2370 7435
rect 2238 6677 2266 6678
rect 2238 6651 2239 6677
rect 2239 6651 2265 6677
rect 2265 6651 2266 6677
rect 2238 6650 2266 6651
rect 2290 6677 2318 6678
rect 2290 6651 2291 6677
rect 2291 6651 2317 6677
rect 2317 6651 2318 6677
rect 2290 6650 2318 6651
rect 2342 6677 2370 6678
rect 2342 6651 2343 6677
rect 2343 6651 2369 6677
rect 2369 6651 2370 6677
rect 2342 6650 2370 6651
rect 8134 6510 8162 6538
rect 2238 5893 2266 5894
rect 2238 5867 2239 5893
rect 2239 5867 2265 5893
rect 2265 5867 2266 5893
rect 2238 5866 2266 5867
rect 2290 5893 2318 5894
rect 2290 5867 2291 5893
rect 2291 5867 2317 5893
rect 2317 5867 2318 5893
rect 2290 5866 2318 5867
rect 2342 5893 2370 5894
rect 2342 5867 2343 5893
rect 2343 5867 2369 5893
rect 2369 5867 2370 5893
rect 2342 5866 2370 5867
rect 2238 5109 2266 5110
rect 2238 5083 2239 5109
rect 2239 5083 2265 5109
rect 2265 5083 2266 5109
rect 2238 5082 2266 5083
rect 2290 5109 2318 5110
rect 2290 5083 2291 5109
rect 2291 5083 2317 5109
rect 2317 5083 2318 5109
rect 2290 5082 2318 5083
rect 2342 5109 2370 5110
rect 2342 5083 2343 5109
rect 2343 5083 2369 5109
rect 2369 5083 2370 5109
rect 2342 5082 2370 5083
rect 2238 4325 2266 4326
rect 2238 4299 2239 4325
rect 2239 4299 2265 4325
rect 2265 4299 2266 4325
rect 2238 4298 2266 4299
rect 2290 4325 2318 4326
rect 2290 4299 2291 4325
rect 2291 4299 2317 4325
rect 2317 4299 2318 4325
rect 2290 4298 2318 4299
rect 2342 4325 2370 4326
rect 2342 4299 2343 4325
rect 2343 4299 2369 4325
rect 2369 4299 2370 4325
rect 2342 4298 2370 4299
rect 9366 9617 9394 9618
rect 9366 9591 9367 9617
rect 9367 9591 9393 9617
rect 9393 9591 9394 9617
rect 9366 9590 9394 9591
rect 9590 10542 9618 10570
rect 9534 9870 9562 9898
rect 9422 9478 9450 9506
rect 9366 9422 9394 9450
rect 9254 9142 9282 9170
rect 9478 9254 9506 9282
rect 9918 11773 9946 11774
rect 9918 11747 9919 11773
rect 9919 11747 9945 11773
rect 9945 11747 9946 11773
rect 9918 11746 9946 11747
rect 9970 11773 9998 11774
rect 9970 11747 9971 11773
rect 9971 11747 9997 11773
rect 9997 11747 9998 11773
rect 9970 11746 9998 11747
rect 10022 11773 10050 11774
rect 10022 11747 10023 11773
rect 10023 11747 10049 11773
rect 10049 11747 10050 11773
rect 10022 11746 10050 11747
rect 10094 11774 10122 11802
rect 10094 11689 10122 11690
rect 10094 11663 10095 11689
rect 10095 11663 10121 11689
rect 10121 11663 10122 11689
rect 10094 11662 10122 11663
rect 9870 11633 9898 11634
rect 9870 11607 9871 11633
rect 9871 11607 9897 11633
rect 9897 11607 9898 11633
rect 9870 11606 9898 11607
rect 9926 11465 9954 11466
rect 9926 11439 9927 11465
rect 9927 11439 9953 11465
rect 9953 11439 9954 11465
rect 9926 11438 9954 11439
rect 10654 11942 10682 11970
rect 10710 11886 10738 11914
rect 11494 13481 11522 13482
rect 11494 13455 11495 13481
rect 11495 13455 11521 13481
rect 11521 13455 11522 13481
rect 11494 13454 11522 13455
rect 11382 13425 11410 13426
rect 11382 13399 11383 13425
rect 11383 13399 11409 13425
rect 11409 13399 11410 13425
rect 11382 13398 11410 13399
rect 12222 13454 12250 13482
rect 11718 13118 11746 13146
rect 12110 13398 12138 13426
rect 12166 13118 12194 13146
rect 12670 13817 12698 13818
rect 12670 13791 12671 13817
rect 12671 13791 12697 13817
rect 12697 13791 12698 13817
rect 12670 13790 12698 13791
rect 12670 13566 12698 13594
rect 12110 12726 12138 12754
rect 11438 12641 11466 12642
rect 11438 12615 11439 12641
rect 11439 12615 11465 12641
rect 11465 12615 11466 12641
rect 11438 12614 11466 12615
rect 11158 12305 11186 12306
rect 11158 12279 11159 12305
rect 11159 12279 11185 12305
rect 11185 12279 11186 12305
rect 11158 12278 11186 12279
rect 12502 12753 12530 12754
rect 12502 12727 12503 12753
rect 12503 12727 12529 12753
rect 12529 12727 12530 12753
rect 12502 12726 12530 12727
rect 11102 11942 11130 11970
rect 10934 11886 10962 11914
rect 11214 11913 11242 11914
rect 11214 11887 11215 11913
rect 11215 11887 11241 11913
rect 11241 11887 11242 11913
rect 11214 11886 11242 11887
rect 10878 11774 10906 11802
rect 10150 11102 10178 11130
rect 9918 10989 9946 10990
rect 9918 10963 9919 10989
rect 9919 10963 9945 10989
rect 9945 10963 9946 10989
rect 9918 10962 9946 10963
rect 9970 10989 9998 10990
rect 9970 10963 9971 10989
rect 9971 10963 9997 10989
rect 9997 10963 9998 10989
rect 9970 10962 9998 10963
rect 10022 10989 10050 10990
rect 10022 10963 10023 10989
rect 10023 10963 10049 10989
rect 10049 10963 10050 10989
rect 10022 10962 10050 10963
rect 9758 10318 9786 10346
rect 9702 10262 9730 10290
rect 9702 9702 9730 9730
rect 9758 9673 9786 9674
rect 9758 9647 9759 9673
rect 9759 9647 9785 9673
rect 9785 9647 9786 9673
rect 9758 9646 9786 9647
rect 9590 9198 9618 9226
rect 9702 9561 9730 9562
rect 9702 9535 9703 9561
rect 9703 9535 9729 9561
rect 9729 9535 9730 9561
rect 9702 9534 9730 9535
rect 9198 8441 9226 8442
rect 9198 8415 9199 8441
rect 9199 8415 9225 8441
rect 9225 8415 9226 8441
rect 9198 8414 9226 8415
rect 9478 8414 9506 8442
rect 9918 10205 9946 10206
rect 9918 10179 9919 10205
rect 9919 10179 9945 10205
rect 9945 10179 9946 10205
rect 9918 10178 9946 10179
rect 9970 10205 9998 10206
rect 9970 10179 9971 10205
rect 9971 10179 9997 10205
rect 9997 10179 9998 10205
rect 9970 10178 9998 10179
rect 10022 10205 10050 10206
rect 10022 10179 10023 10205
rect 10023 10179 10049 10205
rect 10049 10179 10050 10205
rect 10022 10178 10050 10179
rect 9926 9953 9954 9954
rect 9926 9927 9927 9953
rect 9927 9927 9953 9953
rect 9953 9927 9954 9953
rect 9926 9926 9954 9927
rect 10206 10262 10234 10290
rect 10094 9814 10122 9842
rect 10150 9702 10178 9730
rect 10430 10401 10458 10402
rect 10430 10375 10431 10401
rect 10431 10375 10457 10401
rect 10457 10375 10458 10401
rect 10430 10374 10458 10375
rect 10206 10065 10234 10066
rect 10206 10039 10207 10065
rect 10207 10039 10233 10065
rect 10233 10039 10234 10065
rect 10206 10038 10234 10039
rect 10766 11185 10794 11186
rect 10766 11159 10767 11185
rect 10767 11159 10793 11185
rect 10793 11159 10794 11185
rect 10766 11158 10794 11159
rect 10654 10401 10682 10402
rect 10654 10375 10655 10401
rect 10655 10375 10681 10401
rect 10681 10375 10682 10401
rect 10654 10374 10682 10375
rect 10598 9982 10626 10010
rect 10206 9617 10234 9618
rect 10206 9591 10207 9617
rect 10207 9591 10233 9617
rect 10233 9591 10234 9617
rect 10206 9590 10234 9591
rect 10262 9814 10290 9842
rect 9918 9421 9946 9422
rect 9918 9395 9919 9421
rect 9919 9395 9945 9421
rect 9945 9395 9946 9421
rect 9918 9394 9946 9395
rect 9970 9421 9998 9422
rect 9970 9395 9971 9421
rect 9971 9395 9997 9421
rect 9997 9395 9998 9421
rect 9970 9394 9998 9395
rect 10022 9421 10050 9422
rect 10022 9395 10023 9421
rect 10023 9395 10049 9421
rect 10049 9395 10050 9421
rect 10022 9394 10050 9395
rect 10150 9225 10178 9226
rect 10150 9199 10151 9225
rect 10151 9199 10177 9225
rect 10177 9199 10178 9225
rect 10150 9198 10178 9199
rect 9870 9142 9898 9170
rect 10654 9814 10682 9842
rect 10654 9617 10682 9618
rect 10654 9591 10655 9617
rect 10655 9591 10681 9617
rect 10681 9591 10682 9617
rect 10654 9590 10682 9591
rect 10878 10822 10906 10850
rect 11046 11494 11074 11522
rect 11382 11857 11410 11858
rect 11382 11831 11383 11857
rect 11383 11831 11409 11857
rect 11409 11831 11410 11857
rect 11382 11830 11410 11831
rect 11550 11774 11578 11802
rect 12222 11830 12250 11858
rect 11998 11774 12026 11802
rect 11046 10990 11074 11018
rect 11102 11214 11130 11242
rect 11046 10065 11074 10066
rect 11046 10039 11047 10065
rect 11047 10039 11073 10065
rect 11073 10039 11074 10065
rect 11046 10038 11074 10039
rect 10822 9729 10850 9730
rect 10822 9703 10823 9729
rect 10823 9703 10849 9729
rect 10849 9703 10850 9729
rect 10822 9702 10850 9703
rect 10766 9534 10794 9562
rect 9918 8637 9946 8638
rect 9918 8611 9919 8637
rect 9919 8611 9945 8637
rect 9945 8611 9946 8637
rect 9918 8610 9946 8611
rect 9970 8637 9998 8638
rect 9970 8611 9971 8637
rect 9971 8611 9997 8637
rect 9997 8611 9998 8637
rect 9970 8610 9998 8611
rect 10022 8637 10050 8638
rect 10022 8611 10023 8637
rect 10023 8611 10049 8637
rect 10049 8611 10050 8637
rect 10022 8610 10050 8611
rect 9590 8022 9618 8050
rect 9814 8414 9842 8442
rect 9702 7910 9730 7938
rect 9366 7574 9394 7602
rect 9310 7153 9338 7154
rect 9310 7127 9311 7153
rect 9311 7127 9337 7153
rect 9337 7127 9338 7153
rect 9310 7126 9338 7127
rect 10094 8049 10122 8050
rect 10094 8023 10095 8049
rect 10095 8023 10121 8049
rect 10121 8023 10122 8049
rect 10094 8022 10122 8023
rect 9918 7853 9946 7854
rect 9918 7827 9919 7853
rect 9919 7827 9945 7853
rect 9945 7827 9946 7853
rect 9918 7826 9946 7827
rect 9970 7853 9998 7854
rect 9970 7827 9971 7853
rect 9971 7827 9997 7853
rect 9997 7827 9998 7853
rect 9970 7826 9998 7827
rect 10022 7853 10050 7854
rect 10022 7827 10023 7853
rect 10023 7827 10049 7853
rect 10049 7827 10050 7853
rect 10022 7826 10050 7827
rect 10318 8918 10346 8946
rect 10374 9142 10402 9170
rect 10990 9561 11018 9562
rect 10990 9535 10991 9561
rect 10991 9535 11017 9561
rect 11017 9535 11018 9561
rect 10990 9534 11018 9535
rect 10766 9142 10794 9170
rect 10710 8918 10738 8946
rect 10710 8833 10738 8834
rect 10710 8807 10711 8833
rect 10711 8807 10737 8833
rect 10737 8807 10738 8833
rect 10710 8806 10738 8807
rect 11046 8806 11074 8834
rect 10206 8721 10234 8722
rect 10206 8695 10207 8721
rect 10207 8695 10233 8721
rect 10233 8695 10234 8721
rect 10206 8694 10234 8695
rect 10710 8694 10738 8722
rect 10262 8049 10290 8050
rect 10262 8023 10263 8049
rect 10263 8023 10289 8049
rect 10289 8023 10290 8049
rect 10262 8022 10290 8023
rect 10934 8694 10962 8722
rect 11270 11185 11298 11186
rect 11270 11159 11271 11185
rect 11271 11159 11297 11185
rect 11297 11159 11298 11185
rect 11270 11158 11298 11159
rect 11158 10542 11186 10570
rect 11382 10598 11410 10626
rect 11326 10318 11354 10346
rect 11606 11214 11634 11242
rect 11662 11438 11690 11466
rect 11494 10849 11522 10850
rect 11494 10823 11495 10849
rect 11495 10823 11521 10849
rect 11521 10823 11522 10849
rect 11494 10822 11522 10823
rect 11438 10038 11466 10066
rect 11550 10598 11578 10626
rect 11214 10009 11242 10010
rect 11214 9983 11215 10009
rect 11215 9983 11241 10009
rect 11241 9983 11242 10009
rect 11214 9982 11242 9983
rect 11158 9030 11186 9058
rect 11158 8918 11186 8946
rect 11438 9281 11466 9282
rect 11438 9255 11439 9281
rect 11439 9255 11465 9281
rect 11465 9255 11466 9281
rect 11438 9254 11466 9255
rect 11662 10094 11690 10122
rect 11718 9982 11746 10010
rect 11718 9870 11746 9898
rect 11606 9142 11634 9170
rect 11774 9926 11802 9954
rect 11774 9310 11802 9338
rect 11270 8918 11298 8946
rect 11270 8638 11298 8666
rect 11326 8694 11354 8722
rect 11438 8721 11466 8722
rect 11438 8695 11439 8721
rect 11439 8695 11465 8721
rect 11465 8695 11466 8721
rect 11438 8694 11466 8695
rect 10878 8022 10906 8050
rect 10822 7910 10850 7938
rect 10206 7518 10234 7546
rect 9366 6510 9394 6538
rect 9918 7069 9946 7070
rect 9918 7043 9919 7069
rect 9919 7043 9945 7069
rect 9945 7043 9946 7069
rect 9918 7042 9946 7043
rect 9970 7069 9998 7070
rect 9970 7043 9971 7069
rect 9971 7043 9997 7069
rect 9997 7043 9998 7069
rect 9970 7042 9998 7043
rect 10022 7069 10050 7070
rect 10022 7043 10023 7069
rect 10023 7043 10049 7069
rect 10049 7043 10050 7069
rect 10022 7042 10050 7043
rect 10374 6734 10402 6762
rect 9814 6537 9842 6538
rect 9814 6511 9815 6537
rect 9815 6511 9841 6537
rect 9841 6511 9842 6537
rect 9814 6510 9842 6511
rect 9918 6285 9946 6286
rect 9918 6259 9919 6285
rect 9919 6259 9945 6285
rect 9945 6259 9946 6285
rect 9918 6258 9946 6259
rect 9970 6285 9998 6286
rect 9970 6259 9971 6285
rect 9971 6259 9997 6285
rect 9997 6259 9998 6285
rect 9970 6258 9998 6259
rect 10022 6285 10050 6286
rect 10022 6259 10023 6285
rect 10023 6259 10049 6285
rect 10049 6259 10050 6285
rect 10022 6258 10050 6259
rect 9918 5501 9946 5502
rect 9918 5475 9919 5501
rect 9919 5475 9945 5501
rect 9945 5475 9946 5501
rect 9918 5474 9946 5475
rect 9970 5501 9998 5502
rect 9970 5475 9971 5501
rect 9971 5475 9997 5501
rect 9997 5475 9998 5501
rect 9970 5474 9998 5475
rect 10022 5501 10050 5502
rect 10022 5475 10023 5501
rect 10023 5475 10049 5501
rect 10049 5475 10050 5501
rect 10022 5474 10050 5475
rect 9918 4717 9946 4718
rect 9918 4691 9919 4717
rect 9919 4691 9945 4717
rect 9945 4691 9946 4717
rect 9918 4690 9946 4691
rect 9970 4717 9998 4718
rect 9970 4691 9971 4717
rect 9971 4691 9997 4717
rect 9997 4691 9998 4717
rect 9970 4690 9998 4691
rect 10022 4717 10050 4718
rect 10022 4691 10023 4717
rect 10023 4691 10049 4717
rect 10049 4691 10050 4717
rect 10022 4690 10050 4691
rect 10990 7742 11018 7770
rect 11326 8441 11354 8442
rect 11326 8415 11327 8441
rect 11327 8415 11353 8441
rect 11353 8415 11354 8441
rect 11326 8414 11354 8415
rect 11774 8414 11802 8442
rect 11886 8721 11914 8722
rect 11886 8695 11887 8721
rect 11887 8695 11913 8721
rect 11913 8695 11914 8721
rect 11886 8694 11914 8695
rect 12782 13145 12810 13146
rect 12782 13119 12783 13145
rect 12783 13119 12809 13145
rect 12809 13119 12810 13145
rect 12782 13118 12810 13119
rect 12502 12222 12530 12250
rect 13062 13790 13090 13818
rect 17598 15301 17626 15302
rect 17598 15275 17599 15301
rect 17599 15275 17625 15301
rect 17625 15275 17626 15301
rect 17598 15274 17626 15275
rect 17650 15301 17678 15302
rect 17650 15275 17651 15301
rect 17651 15275 17677 15301
rect 17677 15275 17678 15301
rect 17650 15274 17678 15275
rect 17702 15301 17730 15302
rect 17702 15275 17703 15301
rect 17703 15275 17729 15301
rect 17729 15275 17730 15301
rect 17702 15274 17730 15275
rect 17598 14517 17626 14518
rect 17598 14491 17599 14517
rect 17599 14491 17625 14517
rect 17625 14491 17626 14517
rect 17598 14490 17626 14491
rect 17650 14517 17678 14518
rect 17650 14491 17651 14517
rect 17651 14491 17677 14517
rect 17677 14491 17678 14517
rect 17650 14490 17678 14491
rect 17702 14517 17730 14518
rect 17702 14491 17703 14517
rect 17703 14491 17729 14517
rect 17729 14491 17730 14517
rect 17702 14490 17730 14491
rect 18830 13929 18858 13930
rect 18830 13903 18831 13929
rect 18831 13903 18857 13929
rect 18857 13903 18858 13929
rect 18830 13902 18858 13903
rect 13734 13873 13762 13874
rect 13734 13847 13735 13873
rect 13735 13847 13761 13873
rect 13761 13847 13762 13873
rect 13734 13846 13762 13847
rect 14238 13846 14266 13874
rect 13678 13817 13706 13818
rect 13678 13791 13679 13817
rect 13679 13791 13705 13817
rect 13705 13791 13706 13817
rect 13678 13790 13706 13791
rect 13118 13593 13146 13594
rect 13118 13567 13119 13593
rect 13119 13567 13145 13593
rect 13145 13567 13146 13593
rect 13118 13566 13146 13567
rect 13342 13118 13370 13146
rect 20006 13817 20034 13818
rect 20006 13791 20007 13817
rect 20007 13791 20033 13817
rect 20033 13791 20034 13817
rect 20006 13790 20034 13791
rect 17598 13733 17626 13734
rect 17598 13707 17599 13733
rect 17599 13707 17625 13733
rect 17625 13707 17626 13733
rect 17598 13706 17626 13707
rect 17650 13733 17678 13734
rect 17650 13707 17651 13733
rect 17651 13707 17677 13733
rect 17677 13707 17678 13733
rect 17650 13706 17678 13707
rect 17702 13733 17730 13734
rect 17702 13707 17703 13733
rect 17703 13707 17729 13733
rect 17729 13707 17730 13733
rect 17702 13706 17730 13707
rect 13342 12838 13370 12866
rect 13622 12838 13650 12866
rect 13118 12697 13146 12698
rect 13118 12671 13119 12697
rect 13119 12671 13145 12697
rect 13145 12671 13146 12697
rect 13118 12670 13146 12671
rect 12838 12222 12866 12250
rect 12390 11774 12418 11802
rect 12782 11046 12810 11074
rect 12726 10710 12754 10738
rect 12558 10345 12586 10346
rect 12558 10319 12559 10345
rect 12559 10319 12585 10345
rect 12585 10319 12586 10345
rect 12558 10318 12586 10319
rect 12278 10065 12306 10066
rect 12278 10039 12279 10065
rect 12279 10039 12305 10065
rect 12305 10039 12306 10065
rect 12278 10038 12306 10039
rect 12222 9926 12250 9954
rect 12670 9926 12698 9954
rect 12278 9897 12306 9898
rect 12278 9871 12279 9897
rect 12279 9871 12305 9897
rect 12305 9871 12306 9897
rect 12278 9870 12306 9871
rect 12110 9814 12138 9842
rect 12782 10094 12810 10122
rect 17598 12949 17626 12950
rect 17598 12923 17599 12949
rect 17599 12923 17625 12949
rect 17625 12923 17626 12949
rect 17598 12922 17626 12923
rect 17650 12949 17678 12950
rect 17650 12923 17651 12949
rect 17651 12923 17677 12949
rect 17677 12923 17678 12949
rect 17650 12922 17678 12923
rect 17702 12949 17730 12950
rect 17702 12923 17703 12949
rect 17703 12923 17729 12949
rect 17729 12923 17730 12949
rect 17702 12922 17730 12923
rect 14462 12838 14490 12866
rect 13846 12726 13874 12754
rect 13790 12697 13818 12698
rect 13790 12671 13791 12697
rect 13791 12671 13817 12697
rect 13817 12671 13818 12697
rect 13790 12670 13818 12671
rect 14910 12726 14938 12754
rect 13174 11185 13202 11186
rect 13174 11159 13175 11185
rect 13175 11159 13201 11185
rect 13201 11159 13202 11185
rect 13174 11158 13202 11159
rect 12894 11129 12922 11130
rect 12894 11103 12895 11129
rect 12895 11103 12921 11129
rect 12921 11103 12922 11129
rect 12894 11102 12922 11103
rect 13006 11129 13034 11130
rect 13006 11103 13007 11129
rect 13007 11103 13033 11129
rect 13033 11103 13034 11129
rect 13006 11102 13034 11103
rect 13398 11102 13426 11130
rect 13566 11214 13594 11242
rect 13734 10990 13762 11018
rect 13286 10737 13314 10738
rect 13286 10711 13287 10737
rect 13287 10711 13313 10737
rect 13313 10711 13314 10737
rect 13286 10710 13314 10711
rect 13622 10681 13650 10682
rect 13622 10655 13623 10681
rect 13623 10655 13649 10681
rect 13649 10655 13650 10681
rect 13622 10654 13650 10655
rect 12950 10374 12978 10402
rect 12838 9982 12866 10010
rect 12726 9702 12754 9730
rect 12782 9646 12810 9674
rect 12166 9478 12194 9506
rect 12110 9225 12138 9226
rect 12110 9199 12111 9225
rect 12111 9199 12137 9225
rect 12137 9199 12138 9225
rect 12110 9198 12138 9199
rect 12054 8862 12082 8890
rect 11438 7742 11466 7770
rect 11998 8414 12026 8442
rect 11550 7713 11578 7714
rect 11550 7687 11551 7713
rect 11551 7687 11577 7713
rect 11577 7687 11578 7713
rect 11550 7686 11578 7687
rect 10878 7574 10906 7602
rect 11102 7601 11130 7602
rect 11102 7575 11103 7601
rect 11103 7575 11129 7601
rect 11129 7575 11130 7601
rect 11102 7574 11130 7575
rect 11662 8049 11690 8050
rect 11662 8023 11663 8049
rect 11663 8023 11689 8049
rect 11689 8023 11690 8049
rect 11662 8022 11690 8023
rect 11830 7686 11858 7714
rect 11662 7657 11690 7658
rect 11662 7631 11663 7657
rect 11663 7631 11689 7657
rect 11689 7631 11690 7657
rect 11662 7630 11690 7631
rect 11774 7518 11802 7546
rect 11102 6678 11130 6706
rect 11550 7153 11578 7154
rect 11550 7127 11551 7153
rect 11551 7127 11577 7153
rect 11577 7127 11578 7153
rect 11550 7126 11578 7127
rect 11774 7126 11802 7154
rect 12110 7769 12138 7770
rect 12110 7743 12111 7769
rect 12111 7743 12137 7769
rect 12137 7743 12138 7769
rect 12110 7742 12138 7743
rect 11886 7630 11914 7658
rect 11998 7518 12026 7546
rect 12166 7518 12194 7546
rect 11998 6902 12026 6930
rect 12110 7126 12138 7154
rect 12222 6958 12250 6986
rect 11942 6678 11970 6706
rect 12726 7630 12754 7658
rect 12894 9758 12922 9786
rect 12894 9505 12922 9506
rect 12894 9479 12895 9505
rect 12895 9479 12921 9505
rect 12921 9479 12922 9505
rect 12894 9478 12922 9479
rect 13062 10038 13090 10066
rect 13454 9926 13482 9954
rect 13734 10150 13762 10178
rect 13510 9870 13538 9898
rect 13174 9729 13202 9730
rect 13174 9703 13175 9729
rect 13175 9703 13201 9729
rect 13201 9703 13202 9729
rect 13174 9702 13202 9703
rect 18830 12753 18858 12754
rect 18830 12727 18831 12753
rect 18831 12727 18857 12753
rect 18857 12727 18858 12753
rect 18830 12726 18858 12727
rect 20006 12446 20034 12474
rect 14014 11494 14042 11522
rect 13902 11241 13930 11242
rect 13902 11215 13903 11241
rect 13903 11215 13929 11241
rect 13929 11215 13930 11241
rect 13902 11214 13930 11215
rect 14014 11158 14042 11186
rect 13846 11046 13874 11074
rect 13846 10737 13874 10738
rect 13846 10711 13847 10737
rect 13847 10711 13873 10737
rect 13873 10711 13874 10737
rect 13846 10710 13874 10711
rect 13622 9702 13650 9730
rect 12894 9310 12922 9338
rect 13062 9366 13090 9394
rect 12950 9225 12978 9226
rect 12950 9199 12951 9225
rect 12951 9199 12977 9225
rect 12977 9199 12978 9225
rect 12950 9198 12978 9199
rect 13006 8358 13034 8386
rect 13174 9198 13202 9226
rect 13398 9142 13426 9170
rect 13398 8833 13426 8834
rect 13398 8807 13399 8833
rect 13399 8807 13425 8833
rect 13425 8807 13426 8833
rect 13398 8806 13426 8807
rect 13566 9198 13594 9226
rect 14070 10654 14098 10682
rect 14070 10401 14098 10402
rect 14070 10375 14071 10401
rect 14071 10375 14097 10401
rect 14097 10375 14098 10401
rect 14070 10374 14098 10375
rect 14798 11521 14826 11522
rect 14798 11495 14799 11521
rect 14799 11495 14825 11521
rect 14825 11495 14826 11521
rect 14798 11494 14826 11495
rect 17598 12165 17626 12166
rect 17598 12139 17599 12165
rect 17599 12139 17625 12165
rect 17625 12139 17626 12165
rect 17598 12138 17626 12139
rect 17650 12165 17678 12166
rect 17650 12139 17651 12165
rect 17651 12139 17677 12165
rect 17677 12139 17678 12165
rect 17650 12138 17678 12139
rect 17702 12165 17730 12166
rect 17702 12139 17703 12165
rect 17703 12139 17729 12165
rect 17729 12139 17730 12165
rect 17702 12138 17730 12139
rect 20006 11774 20034 11802
rect 18830 11494 18858 11522
rect 14406 10737 14434 10738
rect 14406 10711 14407 10737
rect 14407 10711 14433 10737
rect 14433 10711 14434 10737
rect 14406 10710 14434 10711
rect 15470 10737 15498 10738
rect 15470 10711 15471 10737
rect 15471 10711 15497 10737
rect 15497 10711 15498 10737
rect 15470 10710 15498 10711
rect 17598 11381 17626 11382
rect 17598 11355 17599 11381
rect 17599 11355 17625 11381
rect 17625 11355 17626 11381
rect 17598 11354 17626 11355
rect 17650 11381 17678 11382
rect 17650 11355 17651 11381
rect 17651 11355 17677 11381
rect 17677 11355 17678 11381
rect 17650 11354 17678 11355
rect 17702 11381 17730 11382
rect 17702 11355 17703 11381
rect 17703 11355 17729 11381
rect 17729 11355 17730 11381
rect 17702 11354 17730 11355
rect 14238 10401 14266 10402
rect 14238 10375 14239 10401
rect 14239 10375 14265 10401
rect 14265 10375 14266 10401
rect 14238 10374 14266 10375
rect 15470 10374 15498 10402
rect 14014 9926 14042 9954
rect 13902 9758 13930 9786
rect 13734 9505 13762 9506
rect 13734 9479 13735 9505
rect 13735 9479 13761 9505
rect 13761 9479 13762 9505
rect 13734 9478 13762 9479
rect 13846 9310 13874 9338
rect 13734 9198 13762 9226
rect 14014 9254 14042 9282
rect 14014 8833 14042 8834
rect 14014 8807 14015 8833
rect 14015 8807 14041 8833
rect 14041 8807 14042 8833
rect 14014 8806 14042 8807
rect 14182 10094 14210 10122
rect 14462 9953 14490 9954
rect 14462 9927 14463 9953
rect 14463 9927 14489 9953
rect 14489 9927 14490 9953
rect 14462 9926 14490 9927
rect 14182 9534 14210 9562
rect 14126 8862 14154 8890
rect 14238 9310 14266 9338
rect 14574 9561 14602 9562
rect 14574 9535 14575 9561
rect 14575 9535 14601 9561
rect 14601 9535 14602 9561
rect 14574 9534 14602 9535
rect 14462 9254 14490 9282
rect 14238 9142 14266 9170
rect 14574 8833 14602 8834
rect 14574 8807 14575 8833
rect 14575 8807 14601 8833
rect 14601 8807 14602 8833
rect 14574 8806 14602 8807
rect 14238 8694 14266 8722
rect 14070 8638 14098 8666
rect 15470 9478 15498 9506
rect 14686 9366 14714 9394
rect 15246 9366 15274 9394
rect 14686 8777 14714 8778
rect 14686 8751 14687 8777
rect 14687 8751 14713 8777
rect 14713 8751 14714 8777
rect 14686 8750 14714 8751
rect 14854 8694 14882 8722
rect 14238 8497 14266 8498
rect 14238 8471 14239 8497
rect 14239 8471 14265 8497
rect 14265 8471 14266 8497
rect 14238 8470 14266 8471
rect 13118 8358 13146 8386
rect 13510 8358 13538 8386
rect 13230 7657 13258 7658
rect 13230 7631 13231 7657
rect 13231 7631 13257 7657
rect 13257 7631 13258 7657
rect 13230 7630 13258 7631
rect 13398 7657 13426 7658
rect 13398 7631 13399 7657
rect 13399 7631 13425 7657
rect 13425 7631 13426 7657
rect 13398 7630 13426 7631
rect 15526 9254 15554 9282
rect 20006 10766 20034 10794
rect 18830 10710 18858 10738
rect 17598 10597 17626 10598
rect 17598 10571 17599 10597
rect 17599 10571 17625 10597
rect 17625 10571 17626 10597
rect 17598 10570 17626 10571
rect 17650 10597 17678 10598
rect 17650 10571 17651 10597
rect 17651 10571 17677 10597
rect 17677 10571 17678 10597
rect 17650 10570 17678 10571
rect 17702 10597 17730 10598
rect 17702 10571 17703 10597
rect 17703 10571 17729 10597
rect 17729 10571 17730 10597
rect 17702 10570 17730 10571
rect 17598 9813 17626 9814
rect 17598 9787 17599 9813
rect 17599 9787 17625 9813
rect 17625 9787 17626 9813
rect 17598 9786 17626 9787
rect 17650 9813 17678 9814
rect 17650 9787 17651 9813
rect 17651 9787 17677 9813
rect 17677 9787 17678 9813
rect 17650 9786 17678 9787
rect 17702 9813 17730 9814
rect 17702 9787 17703 9813
rect 17703 9787 17729 9813
rect 17729 9787 17730 9813
rect 17702 9786 17730 9787
rect 20006 10094 20034 10122
rect 18830 9478 18858 9506
rect 15470 8862 15498 8890
rect 15134 8638 15162 8666
rect 15246 8750 15274 8778
rect 15078 8470 15106 8498
rect 15246 8414 15274 8442
rect 13062 7126 13090 7154
rect 12726 6985 12754 6986
rect 12726 6959 12727 6985
rect 12727 6959 12753 6985
rect 12753 6959 12754 6985
rect 12726 6958 12754 6959
rect 13454 7126 13482 7154
rect 12558 6902 12586 6930
rect 12334 6790 12362 6818
rect 12670 6817 12698 6818
rect 12670 6791 12671 6817
rect 12671 6791 12697 6817
rect 12697 6791 12698 6817
rect 12670 6790 12698 6791
rect 12782 6678 12810 6706
rect 2238 3541 2266 3542
rect 2238 3515 2239 3541
rect 2239 3515 2265 3541
rect 2265 3515 2266 3541
rect 2238 3514 2266 3515
rect 2290 3541 2318 3542
rect 2290 3515 2291 3541
rect 2291 3515 2317 3541
rect 2317 3515 2318 3541
rect 2290 3514 2318 3515
rect 2342 3541 2370 3542
rect 2342 3515 2343 3541
rect 2343 3515 2369 3541
rect 2369 3515 2370 3541
rect 2342 3514 2370 3515
rect 2238 2757 2266 2758
rect 2238 2731 2239 2757
rect 2239 2731 2265 2757
rect 2265 2731 2266 2757
rect 2238 2730 2266 2731
rect 2290 2757 2318 2758
rect 2290 2731 2291 2757
rect 2291 2731 2317 2757
rect 2317 2731 2318 2757
rect 2290 2730 2318 2731
rect 2342 2757 2370 2758
rect 2342 2731 2343 2757
rect 2343 2731 2369 2757
rect 2369 2731 2370 2757
rect 2342 2730 2370 2731
rect 2238 1973 2266 1974
rect 2238 1947 2239 1973
rect 2239 1947 2265 1973
rect 2265 1947 2266 1973
rect 2238 1946 2266 1947
rect 2290 1973 2318 1974
rect 2290 1947 2291 1973
rect 2291 1947 2317 1973
rect 2317 1947 2318 1973
rect 2290 1946 2318 1947
rect 2342 1973 2370 1974
rect 2342 1947 2343 1973
rect 2343 1947 2369 1973
rect 2369 1947 2370 1973
rect 2342 1946 2370 1947
rect 9918 3933 9946 3934
rect 9918 3907 9919 3933
rect 9919 3907 9945 3933
rect 9945 3907 9946 3933
rect 9918 3906 9946 3907
rect 9970 3933 9998 3934
rect 9970 3907 9971 3933
rect 9971 3907 9997 3933
rect 9997 3907 9998 3933
rect 9970 3906 9998 3907
rect 10022 3933 10050 3934
rect 10022 3907 10023 3933
rect 10023 3907 10049 3933
rect 10049 3907 10050 3933
rect 10022 3906 10050 3907
rect 9918 3149 9946 3150
rect 9918 3123 9919 3149
rect 9919 3123 9945 3149
rect 9945 3123 9946 3149
rect 9918 3122 9946 3123
rect 9970 3149 9998 3150
rect 9970 3123 9971 3149
rect 9971 3123 9997 3149
rect 9997 3123 9998 3149
rect 9970 3122 9998 3123
rect 10022 3149 10050 3150
rect 10022 3123 10023 3149
rect 10023 3123 10049 3149
rect 10049 3123 10050 3149
rect 10022 3122 10050 3123
rect 9918 2365 9946 2366
rect 9918 2339 9919 2365
rect 9919 2339 9945 2365
rect 9945 2339 9946 2365
rect 9918 2338 9946 2339
rect 9970 2365 9998 2366
rect 9970 2339 9971 2365
rect 9971 2339 9997 2365
rect 9997 2339 9998 2365
rect 9970 2338 9998 2339
rect 10022 2365 10050 2366
rect 10022 2339 10023 2365
rect 10023 2339 10049 2365
rect 10049 2339 10050 2365
rect 10022 2338 10050 2339
rect 10766 1806 10794 1834
rect 8414 1694 8442 1722
rect 9030 1694 9058 1722
rect 9918 1581 9946 1582
rect 9918 1555 9919 1581
rect 9919 1555 9945 1581
rect 9945 1555 9946 1581
rect 9918 1554 9946 1555
rect 9970 1581 9998 1582
rect 9970 1555 9971 1581
rect 9971 1555 9997 1581
rect 9997 1555 9998 1581
rect 9970 1554 9998 1555
rect 10022 1581 10050 1582
rect 10022 1555 10023 1581
rect 10023 1555 10049 1581
rect 10049 1555 10050 1581
rect 10022 1554 10050 1555
rect 11214 1833 11242 1834
rect 11214 1807 11215 1833
rect 11215 1807 11241 1833
rect 11241 1807 11242 1833
rect 11214 1806 11242 1807
rect 11774 1806 11802 1834
rect 13566 7153 13594 7154
rect 13566 7127 13567 7153
rect 13567 7127 13593 7153
rect 13593 7127 13594 7153
rect 13566 7126 13594 7127
rect 13062 6734 13090 6762
rect 14014 7126 14042 7154
rect 14518 7630 14546 7658
rect 17598 9029 17626 9030
rect 17598 9003 17599 9029
rect 17599 9003 17625 9029
rect 17625 9003 17626 9029
rect 17598 9002 17626 9003
rect 17650 9029 17678 9030
rect 17650 9003 17651 9029
rect 17651 9003 17677 9029
rect 17677 9003 17678 9029
rect 17650 9002 17678 9003
rect 17702 9029 17730 9030
rect 17702 9003 17703 9029
rect 17703 9003 17729 9029
rect 17729 9003 17730 9029
rect 17702 9002 17730 9003
rect 18830 8833 18858 8834
rect 18830 8807 18831 8833
rect 18831 8807 18857 8833
rect 18857 8807 18858 8833
rect 18830 8806 18858 8807
rect 20006 8750 20034 8778
rect 18830 8441 18858 8442
rect 18830 8415 18831 8441
rect 18831 8415 18857 8441
rect 18857 8415 18858 8441
rect 18830 8414 18858 8415
rect 20006 8414 20034 8442
rect 17598 8245 17626 8246
rect 17598 8219 17599 8245
rect 17599 8219 17625 8245
rect 17625 8219 17626 8245
rect 17598 8218 17626 8219
rect 17650 8245 17678 8246
rect 17650 8219 17651 8245
rect 17651 8219 17677 8245
rect 17677 8219 17678 8245
rect 17650 8218 17678 8219
rect 17702 8245 17730 8246
rect 17702 8219 17703 8245
rect 17703 8219 17729 8245
rect 17729 8219 17730 8245
rect 17702 8218 17730 8219
rect 18830 7657 18858 7658
rect 18830 7631 18831 7657
rect 18831 7631 18857 7657
rect 18857 7631 18858 7657
rect 18830 7630 18858 7631
rect 17598 7461 17626 7462
rect 17598 7435 17599 7461
rect 17599 7435 17625 7461
rect 17625 7435 17626 7461
rect 17598 7434 17626 7435
rect 17650 7461 17678 7462
rect 17650 7435 17651 7461
rect 17651 7435 17677 7461
rect 17677 7435 17678 7461
rect 17650 7434 17678 7435
rect 17702 7461 17730 7462
rect 17702 7435 17703 7461
rect 17703 7435 17729 7461
rect 17729 7435 17730 7461
rect 17702 7434 17730 7435
rect 20006 7406 20034 7434
rect 14742 7126 14770 7154
rect 13566 6734 13594 6762
rect 17598 6677 17626 6678
rect 17598 6651 17599 6677
rect 17599 6651 17625 6677
rect 17625 6651 17626 6677
rect 17598 6650 17626 6651
rect 17650 6677 17678 6678
rect 17650 6651 17651 6677
rect 17651 6651 17677 6677
rect 17677 6651 17678 6677
rect 17650 6650 17678 6651
rect 17702 6677 17730 6678
rect 17702 6651 17703 6677
rect 17703 6651 17729 6677
rect 17729 6651 17730 6677
rect 17702 6650 17730 6651
rect 17598 5893 17626 5894
rect 17598 5867 17599 5893
rect 17599 5867 17625 5893
rect 17625 5867 17626 5893
rect 17598 5866 17626 5867
rect 17650 5893 17678 5894
rect 17650 5867 17651 5893
rect 17651 5867 17677 5893
rect 17677 5867 17678 5893
rect 17650 5866 17678 5867
rect 17702 5893 17730 5894
rect 17702 5867 17703 5893
rect 17703 5867 17729 5893
rect 17729 5867 17730 5893
rect 17702 5866 17730 5867
rect 17598 5109 17626 5110
rect 17598 5083 17599 5109
rect 17599 5083 17625 5109
rect 17625 5083 17626 5109
rect 17598 5082 17626 5083
rect 17650 5109 17678 5110
rect 17650 5083 17651 5109
rect 17651 5083 17677 5109
rect 17677 5083 17678 5109
rect 17650 5082 17678 5083
rect 17702 5109 17730 5110
rect 17702 5083 17703 5109
rect 17703 5083 17729 5109
rect 17729 5083 17730 5109
rect 17702 5082 17730 5083
rect 17598 4325 17626 4326
rect 17598 4299 17599 4325
rect 17599 4299 17625 4325
rect 17625 4299 17626 4325
rect 17598 4298 17626 4299
rect 17650 4325 17678 4326
rect 17650 4299 17651 4325
rect 17651 4299 17677 4325
rect 17677 4299 17678 4325
rect 17650 4298 17678 4299
rect 17702 4325 17730 4326
rect 17702 4299 17703 4325
rect 17703 4299 17729 4325
rect 17729 4299 17730 4325
rect 17702 4298 17730 4299
rect 12838 2590 12866 2618
rect 12446 2030 12474 2058
rect 12782 1833 12810 1834
rect 12782 1807 12783 1833
rect 12783 1807 12809 1833
rect 12809 1807 12810 1833
rect 12782 1806 12810 1807
rect 17598 3541 17626 3542
rect 17598 3515 17599 3541
rect 17599 3515 17625 3541
rect 17625 3515 17626 3541
rect 17598 3514 17626 3515
rect 17650 3541 17678 3542
rect 17650 3515 17651 3541
rect 17651 3515 17677 3541
rect 17677 3515 17678 3541
rect 17650 3514 17678 3515
rect 17702 3541 17730 3542
rect 17702 3515 17703 3541
rect 17703 3515 17729 3541
rect 17729 3515 17730 3541
rect 17702 3514 17730 3515
rect 17598 2757 17626 2758
rect 17598 2731 17599 2757
rect 17599 2731 17625 2757
rect 17625 2731 17626 2757
rect 17598 2730 17626 2731
rect 17650 2757 17678 2758
rect 17650 2731 17651 2757
rect 17651 2731 17677 2757
rect 17677 2731 17678 2757
rect 17650 2730 17678 2731
rect 17702 2757 17730 2758
rect 17702 2731 17703 2757
rect 17703 2731 17729 2757
rect 17729 2731 17730 2757
rect 17702 2730 17730 2731
rect 13398 2617 13426 2618
rect 13398 2591 13399 2617
rect 13399 2591 13425 2617
rect 13425 2591 13426 2617
rect 13398 2590 13426 2591
rect 13118 2057 13146 2058
rect 13118 2031 13119 2057
rect 13119 2031 13145 2057
rect 13145 2031 13146 2057
rect 13118 2030 13146 2031
rect 17598 1973 17626 1974
rect 17598 1947 17599 1973
rect 17599 1947 17625 1973
rect 17625 1947 17626 1973
rect 17598 1946 17626 1947
rect 17650 1973 17678 1974
rect 17650 1947 17651 1973
rect 17651 1947 17677 1973
rect 17677 1947 17678 1973
rect 17650 1946 17678 1947
rect 17702 1973 17730 1974
rect 17702 1947 17703 1973
rect 17703 1947 17729 1973
rect 17729 1947 17730 1973
rect 17702 1946 17730 1947
<< metal3 >>
rect 2233 19194 2238 19222
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2370 19194 2375 19222
rect 17593 19194 17598 19222
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17730 19194 17735 19222
rect 8073 19110 8078 19138
rect 8106 19110 8974 19138
rect 9002 19110 9007 19138
rect 10425 19110 10430 19138
rect 10458 19110 11046 19138
rect 11074 19110 11079 19138
rect 12105 19110 12110 19138
rect 12138 19110 12782 19138
rect 12810 19110 12815 19138
rect 9913 18802 9918 18830
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 10050 18802 10055 18830
rect 9417 18718 9422 18746
rect 9450 18718 10038 18746
rect 10066 18718 10071 18746
rect 13113 18718 13118 18746
rect 13146 18718 13734 18746
rect 13762 18718 13767 18746
rect 2233 18410 2238 18438
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2370 18410 2375 18438
rect 17593 18410 17598 18438
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17730 18410 17735 18438
rect 7737 18326 7742 18354
rect 7770 18326 8358 18354
rect 8386 18326 8391 18354
rect 9913 18018 9918 18046
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 10050 18018 10055 18046
rect 2233 17626 2238 17654
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2370 17626 2375 17654
rect 17593 17626 17598 17654
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17730 17626 17735 17654
rect 9913 17234 9918 17262
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 10050 17234 10055 17262
rect 2233 16842 2238 16870
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2370 16842 2375 16870
rect 17593 16842 17598 16870
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17730 16842 17735 16870
rect 9913 16450 9918 16478
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 10050 16450 10055 16478
rect 2233 16058 2238 16086
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2370 16058 2375 16086
rect 17593 16058 17598 16086
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17730 16058 17735 16086
rect 9913 15666 9918 15694
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 10050 15666 10055 15694
rect 2233 15274 2238 15302
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2370 15274 2375 15302
rect 17593 15274 17598 15302
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17730 15274 17735 15302
rect 9913 14882 9918 14910
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 10050 14882 10055 14910
rect 2233 14490 2238 14518
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2370 14490 2375 14518
rect 17593 14490 17598 14518
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17730 14490 17735 14518
rect 9913 14098 9918 14126
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 10050 14098 10055 14126
rect 6673 13902 6678 13930
rect 6706 13902 8134 13930
rect 8162 13902 8750 13930
rect 8778 13902 8974 13930
rect 9002 13902 10290 13930
rect 10262 13874 10290 13902
rect 15946 13902 18830 13930
rect 18858 13902 18863 13930
rect 15946 13874 15974 13902
rect 10257 13846 10262 13874
rect 10290 13846 10654 13874
rect 10682 13846 10687 13874
rect 13729 13846 13734 13874
rect 13762 13846 14238 13874
rect 14266 13846 15974 13874
rect 20600 13818 21000 13832
rect 9865 13790 9870 13818
rect 9898 13790 10430 13818
rect 10458 13790 10463 13818
rect 12049 13790 12054 13818
rect 12082 13790 12670 13818
rect 12698 13790 12703 13818
rect 13057 13790 13062 13818
rect 13090 13790 13678 13818
rect 13706 13790 13711 13818
rect 20001 13790 20006 13818
rect 20034 13790 21000 13818
rect 20600 13776 21000 13790
rect 2233 13706 2238 13734
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2370 13706 2375 13734
rect 17593 13706 17598 13734
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17730 13706 17735 13734
rect 12665 13566 12670 13594
rect 12698 13566 13118 13594
rect 13146 13566 13151 13594
rect 0 13482 400 13496
rect 0 13454 2086 13482
rect 2114 13454 2119 13482
rect 7961 13454 7966 13482
rect 7994 13454 8470 13482
rect 8498 13454 9086 13482
rect 9114 13454 9758 13482
rect 9786 13454 9791 13482
rect 11489 13454 11494 13482
rect 11522 13454 12222 13482
rect 12250 13454 12255 13482
rect 0 13440 400 13454
rect 9529 13398 9534 13426
rect 9562 13398 9870 13426
rect 9898 13398 9903 13426
rect 11377 13398 11382 13426
rect 11410 13398 12110 13426
rect 12138 13398 12143 13426
rect 9913 13314 9918 13342
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 10050 13314 10055 13342
rect 8521 13230 8526 13258
rect 8554 13230 8974 13258
rect 9002 13230 9007 13258
rect 9025 13118 9030 13146
rect 9058 13118 9366 13146
rect 9394 13118 9399 13146
rect 10817 13118 10822 13146
rect 10850 13118 11718 13146
rect 11746 13118 12166 13146
rect 12194 13118 12782 13146
rect 12810 13118 13342 13146
rect 13370 13118 13375 13146
rect 7737 13006 7742 13034
rect 7770 13006 8358 13034
rect 8386 13006 8391 13034
rect 9417 13006 9422 13034
rect 9450 13006 9758 13034
rect 9786 13006 9791 13034
rect 2233 12922 2238 12950
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2370 12922 2375 12950
rect 17593 12922 17598 12950
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17730 12922 17735 12950
rect 13337 12838 13342 12866
rect 13370 12838 13622 12866
rect 13650 12838 14462 12866
rect 14490 12838 14495 12866
rect 2137 12726 2142 12754
rect 2170 12726 6734 12754
rect 6762 12726 7630 12754
rect 7658 12726 7663 12754
rect 8353 12726 8358 12754
rect 8386 12726 9030 12754
rect 9058 12726 9063 12754
rect 12105 12726 12110 12754
rect 12138 12726 12502 12754
rect 12530 12726 12535 12754
rect 13841 12726 13846 12754
rect 13874 12726 14910 12754
rect 14938 12726 18830 12754
rect 18858 12726 18863 12754
rect 12502 12698 12530 12726
rect 7289 12670 7294 12698
rect 7322 12670 7798 12698
rect 7826 12670 7831 12698
rect 12502 12670 13118 12698
rect 13146 12670 13790 12698
rect 13818 12670 13823 12698
rect 8745 12614 8750 12642
rect 8778 12614 9226 12642
rect 10369 12614 10374 12642
rect 10402 12614 11438 12642
rect 11466 12614 11471 12642
rect 9198 12586 9226 12614
rect 9198 12558 9534 12586
rect 9562 12558 9567 12586
rect 9913 12530 9918 12558
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 10050 12530 10055 12558
rect 0 12474 400 12488
rect 20600 12474 21000 12488
rect 0 12446 966 12474
rect 994 12446 999 12474
rect 20001 12446 20006 12474
rect 20034 12446 21000 12474
rect 0 12432 400 12446
rect 20600 12432 21000 12446
rect 2137 12334 2142 12362
rect 2170 12334 6902 12362
rect 6930 12334 6935 12362
rect 7546 12334 9590 12362
rect 9618 12334 9623 12362
rect 7546 12306 7574 12334
rect 7345 12278 7350 12306
rect 7378 12278 7574 12306
rect 9529 12278 9534 12306
rect 9562 12278 11158 12306
rect 11186 12278 11191 12306
rect 961 12222 966 12250
rect 994 12222 999 12250
rect 7121 12222 7126 12250
rect 7154 12222 7462 12250
rect 7490 12222 12502 12250
rect 12530 12222 12838 12250
rect 12866 12222 12871 12250
rect 0 12138 400 12152
rect 966 12138 994 12222
rect 2233 12138 2238 12166
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2370 12138 2375 12166
rect 17593 12138 17598 12166
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17730 12138 17735 12166
rect 0 12110 994 12138
rect 0 12096 400 12110
rect 9585 11942 9590 11970
rect 9618 11942 10654 11970
rect 10682 11942 11102 11970
rect 11130 11942 11135 11970
rect 9137 11886 9142 11914
rect 9170 11886 9702 11914
rect 9730 11886 9735 11914
rect 10705 11886 10710 11914
rect 10738 11886 10934 11914
rect 10962 11886 11214 11914
rect 11242 11886 11247 11914
rect 11377 11830 11382 11858
rect 11410 11830 12222 11858
rect 12250 11830 12255 11858
rect 0 11802 400 11816
rect 20600 11802 21000 11816
rect 0 11774 966 11802
rect 994 11774 999 11802
rect 10089 11774 10094 11802
rect 10122 11774 10878 11802
rect 10906 11774 11550 11802
rect 11578 11774 11583 11802
rect 11993 11774 11998 11802
rect 12026 11774 12390 11802
rect 12418 11774 12423 11802
rect 20001 11774 20006 11802
rect 20034 11774 21000 11802
rect 0 11760 400 11774
rect 9913 11746 9918 11774
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 10050 11746 10055 11774
rect 20600 11760 21000 11774
rect 2137 11718 2142 11746
rect 2170 11718 7826 11746
rect 5502 11606 7014 11634
rect 7042 11606 7238 11634
rect 7266 11606 7271 11634
rect 7345 11606 7350 11634
rect 7378 11606 7686 11634
rect 7714 11606 7719 11634
rect 5502 11522 5530 11606
rect 6897 11550 6902 11578
rect 6930 11550 7294 11578
rect 7322 11550 7327 11578
rect 2025 11494 2030 11522
rect 2058 11494 5502 11522
rect 5530 11494 5535 11522
rect 6561 11494 6566 11522
rect 6594 11494 7630 11522
rect 7658 11494 7663 11522
rect 0 11466 400 11480
rect 7798 11466 7826 11718
rect 9249 11662 9254 11690
rect 9282 11662 10094 11690
rect 10122 11662 10127 11690
rect 9473 11606 9478 11634
rect 9506 11606 9870 11634
rect 9898 11606 9903 11634
rect 8969 11494 8974 11522
rect 9002 11494 11046 11522
rect 11074 11494 11079 11522
rect 14009 11494 14014 11522
rect 14042 11494 14798 11522
rect 14826 11494 18830 11522
rect 18858 11494 18863 11522
rect 0 11438 966 11466
rect 994 11438 999 11466
rect 7121 11438 7126 11466
rect 7154 11438 7574 11466
rect 7602 11438 7607 11466
rect 7681 11438 7686 11466
rect 7714 11438 9142 11466
rect 9170 11438 9175 11466
rect 9921 11438 9926 11466
rect 9954 11438 11662 11466
rect 11690 11438 11695 11466
rect 0 11424 400 11438
rect 8857 11382 8862 11410
rect 8890 11382 9310 11410
rect 9338 11382 9343 11410
rect 2233 11354 2238 11382
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2370 11354 2375 11382
rect 17593 11354 17598 11382
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17730 11354 17735 11382
rect 10766 11214 11102 11242
rect 11130 11214 11606 11242
rect 11634 11214 11639 11242
rect 13561 11214 13566 11242
rect 13594 11214 13902 11242
rect 13930 11214 13935 11242
rect 10766 11186 10794 11214
rect 7546 11158 10766 11186
rect 10794 11158 10799 11186
rect 11265 11158 11270 11186
rect 11298 11158 13174 11186
rect 13202 11158 14014 11186
rect 14042 11158 14047 11186
rect 7546 11130 7574 11158
rect 7457 11102 7462 11130
rect 7490 11102 7574 11130
rect 9137 11102 9142 11130
rect 9170 11102 9366 11130
rect 9394 11102 9399 11130
rect 10145 11102 10150 11130
rect 10178 11102 12894 11130
rect 12922 11102 12927 11130
rect 13001 11102 13006 11130
rect 13034 11102 13398 11130
rect 13426 11102 13431 11130
rect 12777 11046 12782 11074
rect 12810 11046 13846 11074
rect 13874 11046 13879 11074
rect 11041 10990 11046 11018
rect 11074 10990 13734 11018
rect 13762 10990 13767 11018
rect 9913 10962 9918 10990
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 10050 10962 10055 10990
rect 10873 10822 10878 10850
rect 10906 10822 11494 10850
rect 11522 10822 11527 10850
rect 20600 10794 21000 10808
rect 2137 10766 2142 10794
rect 2170 10766 4998 10794
rect 5026 10766 5031 10794
rect 20001 10766 20006 10794
rect 20034 10766 21000 10794
rect 20600 10752 21000 10766
rect 12721 10710 12726 10738
rect 12754 10710 13286 10738
rect 13314 10710 13319 10738
rect 13841 10710 13846 10738
rect 13874 10710 14406 10738
rect 14434 10710 14439 10738
rect 15465 10710 15470 10738
rect 15498 10710 18830 10738
rect 18858 10710 18863 10738
rect 13617 10654 13622 10682
rect 13650 10654 14070 10682
rect 14098 10654 14103 10682
rect 6841 10598 6846 10626
rect 6874 10598 6879 10626
rect 7546 10598 11382 10626
rect 11410 10598 11550 10626
rect 11578 10598 11583 10626
rect 2233 10570 2238 10598
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2370 10570 2375 10598
rect 6846 10570 6874 10598
rect 7546 10570 7574 10598
rect 17593 10570 17598 10598
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17730 10570 17735 10598
rect 6846 10542 7014 10570
rect 7042 10542 7574 10570
rect 8521 10542 8526 10570
rect 8554 10542 9590 10570
rect 9618 10542 11158 10570
rect 11186 10542 11191 10570
rect 6953 10486 6958 10514
rect 6986 10486 8470 10514
rect 8498 10486 8974 10514
rect 9002 10486 9007 10514
rect 0 10458 400 10472
rect 0 10430 966 10458
rect 994 10430 999 10458
rect 0 10416 400 10430
rect 2081 10374 2086 10402
rect 2114 10374 10430 10402
rect 10458 10374 10654 10402
rect 10682 10374 10687 10402
rect 12945 10374 12950 10402
rect 12978 10374 14070 10402
rect 14098 10374 14103 10402
rect 14233 10374 14238 10402
rect 14266 10374 15470 10402
rect 15498 10374 15503 10402
rect 4993 10318 4998 10346
rect 5026 10318 6846 10346
rect 6874 10318 6879 10346
rect 9193 10318 9198 10346
rect 9226 10318 9758 10346
rect 9786 10318 9791 10346
rect 11321 10318 11326 10346
rect 11354 10318 12558 10346
rect 12586 10318 12591 10346
rect 6225 10262 6230 10290
rect 6258 10262 6790 10290
rect 6818 10262 6823 10290
rect 7177 10262 7182 10290
rect 7210 10262 9254 10290
rect 9282 10262 9702 10290
rect 9730 10262 10206 10290
rect 10234 10262 10239 10290
rect 9913 10178 9918 10206
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 10050 10178 10055 10206
rect 13729 10150 13734 10178
rect 13762 10150 14210 10178
rect 14182 10122 14210 10150
rect 20600 10122 21000 10136
rect 11657 10094 11662 10122
rect 11690 10094 12782 10122
rect 12810 10094 12815 10122
rect 14177 10094 14182 10122
rect 14210 10094 14215 10122
rect 20001 10094 20006 10122
rect 20034 10094 21000 10122
rect 20600 10080 21000 10094
rect 8857 10038 8862 10066
rect 8890 10038 10206 10066
rect 10234 10038 10239 10066
rect 10318 10038 11046 10066
rect 11074 10038 11079 10066
rect 11433 10038 11438 10066
rect 11466 10038 12278 10066
rect 12306 10038 13062 10066
rect 13090 10038 13095 10066
rect 10318 10010 10346 10038
rect 2137 9982 2142 10010
rect 2170 9982 4942 10010
rect 4970 9982 4975 10010
rect 8409 9982 8414 10010
rect 8442 9982 10346 10010
rect 10593 9982 10598 10010
rect 10626 9982 11214 10010
rect 11242 9982 11247 10010
rect 11713 9982 11718 10010
rect 11746 9982 12838 10010
rect 12866 9982 12871 10010
rect 9193 9926 9198 9954
rect 9226 9926 9926 9954
rect 9954 9926 11774 9954
rect 11802 9926 11807 9954
rect 12217 9926 12222 9954
rect 12250 9926 12670 9954
rect 12698 9926 13454 9954
rect 13482 9926 13487 9954
rect 14009 9926 14014 9954
rect 14042 9926 14462 9954
rect 14490 9926 14495 9954
rect 961 9870 966 9898
rect 994 9870 999 9898
rect 8913 9870 8918 9898
rect 8946 9870 9534 9898
rect 9562 9870 11718 9898
rect 11746 9870 11751 9898
rect 12273 9870 12278 9898
rect 12306 9870 13510 9898
rect 13538 9870 13543 9898
rect 0 9786 400 9800
rect 966 9786 994 9870
rect 10089 9814 10094 9842
rect 10122 9814 10262 9842
rect 10290 9814 10654 9842
rect 10682 9814 12110 9842
rect 12138 9814 12143 9842
rect 2233 9786 2238 9814
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2370 9786 2375 9814
rect 17593 9786 17598 9814
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17730 9786 17735 9814
rect 0 9758 994 9786
rect 12889 9758 12894 9786
rect 12922 9758 13902 9786
rect 13930 9758 13935 9786
rect 0 9744 400 9758
rect 9697 9702 9702 9730
rect 9730 9702 10150 9730
rect 10178 9702 10822 9730
rect 10850 9702 12726 9730
rect 12754 9702 13174 9730
rect 13202 9702 13207 9730
rect 13426 9702 13622 9730
rect 13650 9702 13655 9730
rect 13426 9674 13454 9702
rect 9753 9646 9758 9674
rect 9786 9646 12782 9674
rect 12810 9646 13454 9674
rect 4937 9590 4942 9618
rect 4970 9590 6734 9618
rect 6762 9590 6767 9618
rect 8857 9590 8862 9618
rect 8890 9590 9366 9618
rect 9394 9590 9399 9618
rect 10201 9590 10206 9618
rect 10234 9590 10654 9618
rect 10682 9590 10687 9618
rect 8241 9534 8246 9562
rect 8274 9534 9702 9562
rect 9730 9534 9735 9562
rect 10761 9534 10766 9562
rect 10794 9534 10990 9562
rect 11018 9534 11023 9562
rect 14177 9534 14182 9562
rect 14210 9534 14574 9562
rect 14602 9534 14607 9562
rect 6393 9478 6398 9506
rect 6426 9478 6678 9506
rect 6706 9478 8358 9506
rect 8386 9478 9422 9506
rect 9450 9478 9455 9506
rect 12161 9478 12166 9506
rect 12194 9478 12894 9506
rect 12922 9478 12927 9506
rect 13729 9478 13734 9506
rect 13762 9478 15470 9506
rect 15498 9478 18830 9506
rect 18858 9478 18863 9506
rect 8857 9422 8862 9450
rect 8890 9422 9366 9450
rect 9394 9422 9399 9450
rect 9913 9394 9918 9422
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 10050 9394 10055 9422
rect 13057 9366 13062 9394
rect 13090 9366 14686 9394
rect 14714 9366 15246 9394
rect 15274 9366 15279 9394
rect 6225 9310 6230 9338
rect 6258 9310 8750 9338
rect 8778 9310 8783 9338
rect 11769 9310 11774 9338
rect 11802 9310 12894 9338
rect 12922 9310 12927 9338
rect 13426 9310 13846 9338
rect 13874 9310 14238 9338
rect 14266 9310 14271 9338
rect 13426 9282 13454 9310
rect 6337 9254 6342 9282
rect 6370 9254 6846 9282
rect 6874 9254 6879 9282
rect 9473 9254 9478 9282
rect 9506 9254 10290 9282
rect 11433 9254 11438 9282
rect 11466 9254 13454 9282
rect 14009 9254 14014 9282
rect 14042 9254 14462 9282
rect 14490 9254 15526 9282
rect 15554 9254 15559 9282
rect 10262 9226 10290 9254
rect 6449 9198 6454 9226
rect 6482 9198 7126 9226
rect 7154 9198 7159 9226
rect 7737 9198 7742 9226
rect 7770 9198 8638 9226
rect 8666 9198 8671 9226
rect 9585 9198 9590 9226
rect 9618 9198 10150 9226
rect 10178 9198 10183 9226
rect 10262 9198 11634 9226
rect 12105 9198 12110 9226
rect 12138 9198 12950 9226
rect 12978 9198 13174 9226
rect 13202 9198 13207 9226
rect 13286 9198 13566 9226
rect 13594 9198 13734 9226
rect 13762 9198 13767 9226
rect 11606 9170 11634 9198
rect 13286 9170 13314 9198
rect 9249 9142 9254 9170
rect 9282 9142 9870 9170
rect 9898 9142 10374 9170
rect 10402 9142 10766 9170
rect 10794 9142 10799 9170
rect 11601 9142 11606 9170
rect 11634 9142 13314 9170
rect 13393 9142 13398 9170
rect 13426 9142 14238 9170
rect 14266 9142 14271 9170
rect 8409 9086 8414 9114
rect 8442 9086 8918 9114
rect 8946 9086 8951 9114
rect 13426 9058 13454 9142
rect 8017 9030 8022 9058
rect 8050 9030 11158 9058
rect 11186 9030 13454 9058
rect 2233 9002 2238 9030
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2370 9002 2375 9030
rect 17593 9002 17598 9030
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17730 9002 17735 9030
rect 7793 8974 7798 9002
rect 7826 8974 8470 9002
rect 8498 8974 8974 9002
rect 9002 8974 9007 9002
rect 10313 8918 10318 8946
rect 10346 8918 10710 8946
rect 10738 8918 11158 8946
rect 11186 8918 11270 8946
rect 11298 8918 11303 8946
rect 6393 8862 6398 8890
rect 6426 8862 6958 8890
rect 6986 8862 6991 8890
rect 7121 8862 7126 8890
rect 7154 8862 7742 8890
rect 7770 8862 7775 8890
rect 8409 8862 8414 8890
rect 8442 8862 12054 8890
rect 12082 8862 12087 8890
rect 14121 8862 14126 8890
rect 14154 8862 15470 8890
rect 15498 8862 15974 8890
rect 15946 8834 15974 8862
rect 2137 8806 2142 8834
rect 2170 8806 5558 8834
rect 5586 8806 5591 8834
rect 6897 8806 6902 8834
rect 6930 8806 7462 8834
rect 7490 8806 8722 8834
rect 10705 8806 10710 8834
rect 10738 8806 11046 8834
rect 11074 8806 11079 8834
rect 13393 8806 13398 8834
rect 13426 8806 14014 8834
rect 14042 8806 14574 8834
rect 14602 8806 14607 8834
rect 15946 8806 18830 8834
rect 18858 8806 18863 8834
rect 5558 8778 5586 8806
rect 5558 8750 7014 8778
rect 7042 8750 7047 8778
rect 7233 8750 7238 8778
rect 7266 8750 7271 8778
rect 7737 8750 7742 8778
rect 7770 8750 8134 8778
rect 8162 8750 8167 8778
rect 7238 8722 7266 8750
rect 8694 8722 8722 8806
rect 20600 8778 21000 8792
rect 14681 8750 14686 8778
rect 14714 8750 15246 8778
rect 15274 8750 15279 8778
rect 20001 8750 20006 8778
rect 20034 8750 21000 8778
rect 20600 8736 21000 8750
rect 7238 8694 7574 8722
rect 7625 8694 7630 8722
rect 7658 8694 8414 8722
rect 8442 8694 8447 8722
rect 8689 8694 8694 8722
rect 8722 8694 8727 8722
rect 9814 8694 10206 8722
rect 10234 8694 10710 8722
rect 10738 8694 10934 8722
rect 10962 8694 11326 8722
rect 11354 8694 11359 8722
rect 11433 8694 11438 8722
rect 11466 8694 11886 8722
rect 11914 8694 11919 8722
rect 14233 8694 14238 8722
rect 14266 8694 14854 8722
rect 14882 8694 14887 8722
rect 7546 8666 7574 8694
rect 9814 8666 9842 8694
rect 7546 8638 9842 8666
rect 11265 8638 11270 8666
rect 11298 8638 14070 8666
rect 14098 8638 15134 8666
rect 15162 8638 15167 8666
rect 9913 8610 9918 8638
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 10050 8610 10055 8638
rect 7457 8470 7462 8498
rect 7490 8470 8190 8498
rect 8218 8470 8223 8498
rect 14233 8470 14238 8498
rect 14266 8470 15078 8498
rect 15106 8470 15111 8498
rect 0 8442 400 8456
rect 20600 8442 21000 8456
rect 0 8414 966 8442
rect 994 8414 999 8442
rect 7513 8414 7518 8442
rect 7546 8414 8302 8442
rect 8330 8414 8335 8442
rect 9193 8414 9198 8442
rect 9226 8414 9478 8442
rect 9506 8414 9814 8442
rect 9842 8414 9847 8442
rect 11321 8414 11326 8442
rect 11354 8414 11774 8442
rect 11802 8414 11998 8442
rect 12026 8414 12031 8442
rect 15241 8414 15246 8442
rect 15274 8414 18830 8442
rect 18858 8414 18863 8442
rect 20001 8414 20006 8442
rect 20034 8414 21000 8442
rect 0 8400 400 8414
rect 20600 8400 21000 8414
rect 8241 8358 8246 8386
rect 8274 8358 13006 8386
rect 13034 8358 13039 8386
rect 13113 8358 13118 8386
rect 13146 8358 13510 8386
rect 13538 8358 13543 8386
rect 2233 8218 2238 8246
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2370 8218 2375 8246
rect 17593 8218 17598 8246
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17730 8218 17735 8246
rect 9585 8022 9590 8050
rect 9618 8022 10094 8050
rect 10122 8022 10127 8050
rect 10257 8022 10262 8050
rect 10290 8022 10878 8050
rect 10906 8022 11662 8050
rect 11690 8022 11695 8050
rect 9697 7910 9702 7938
rect 9730 7910 10822 7938
rect 10850 7910 10855 7938
rect 9913 7826 9918 7854
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 10050 7826 10055 7854
rect 10985 7742 10990 7770
rect 11018 7742 11438 7770
rect 11466 7742 12110 7770
rect 12138 7742 12143 7770
rect 11545 7686 11550 7714
rect 11578 7686 11830 7714
rect 11858 7686 11863 7714
rect 11657 7630 11662 7658
rect 11690 7630 11886 7658
rect 11914 7630 12726 7658
rect 12754 7630 13230 7658
rect 13258 7630 13263 7658
rect 13393 7630 13398 7658
rect 13426 7630 14518 7658
rect 14546 7630 18830 7658
rect 18858 7630 18863 7658
rect 6841 7574 6846 7602
rect 6874 7574 7014 7602
rect 7042 7574 8414 7602
rect 8442 7574 9366 7602
rect 9394 7574 10878 7602
rect 10906 7574 10911 7602
rect 10990 7574 11102 7602
rect 11130 7574 11135 7602
rect 10990 7546 11018 7574
rect 10201 7518 10206 7546
rect 10234 7518 11018 7546
rect 11769 7518 11774 7546
rect 11802 7518 11998 7546
rect 12026 7518 12166 7546
rect 12194 7518 12199 7546
rect 2233 7434 2238 7462
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2370 7434 2375 7462
rect 17593 7434 17598 7462
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17730 7434 17735 7462
rect 20600 7434 21000 7448
rect 20001 7406 20006 7434
rect 20034 7406 21000 7434
rect 20600 7392 21000 7406
rect 9305 7126 9310 7154
rect 9338 7126 11550 7154
rect 11578 7126 11583 7154
rect 11769 7126 11774 7154
rect 11802 7126 12110 7154
rect 12138 7126 12143 7154
rect 13057 7126 13062 7154
rect 13090 7126 13454 7154
rect 13482 7126 13487 7154
rect 13561 7126 13566 7154
rect 13594 7126 14014 7154
rect 14042 7126 14742 7154
rect 14770 7126 14775 7154
rect 9913 7042 9918 7070
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 10050 7042 10055 7070
rect 12217 6958 12222 6986
rect 12250 6958 12726 6986
rect 12754 6958 12759 6986
rect 11993 6902 11998 6930
rect 12026 6902 12558 6930
rect 12586 6902 12591 6930
rect 12329 6790 12334 6818
rect 12362 6790 12670 6818
rect 12698 6790 12703 6818
rect 10369 6734 10374 6762
rect 10402 6734 11074 6762
rect 11046 6706 11074 6734
rect 12782 6734 13062 6762
rect 13090 6734 13566 6762
rect 13594 6734 13599 6762
rect 12782 6706 12810 6734
rect 11046 6678 11102 6706
rect 11130 6678 11942 6706
rect 11970 6678 12782 6706
rect 12810 6678 12815 6706
rect 2233 6650 2238 6678
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2370 6650 2375 6678
rect 17593 6650 17598 6678
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17730 6650 17735 6678
rect 8129 6510 8134 6538
rect 8162 6510 9366 6538
rect 9394 6510 9814 6538
rect 9842 6510 9847 6538
rect 9913 6258 9918 6286
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 10050 6258 10055 6286
rect 2233 5866 2238 5894
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2370 5866 2375 5894
rect 17593 5866 17598 5894
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17730 5866 17735 5894
rect 9913 5474 9918 5502
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 10050 5474 10055 5502
rect 2233 5082 2238 5110
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2370 5082 2375 5110
rect 17593 5082 17598 5110
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17730 5082 17735 5110
rect 9913 4690 9918 4718
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 10050 4690 10055 4718
rect 2233 4298 2238 4326
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2370 4298 2375 4326
rect 17593 4298 17598 4326
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17730 4298 17735 4326
rect 9913 3906 9918 3934
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 10050 3906 10055 3934
rect 2233 3514 2238 3542
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2370 3514 2375 3542
rect 17593 3514 17598 3542
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17730 3514 17735 3542
rect 9913 3122 9918 3150
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 10050 3122 10055 3150
rect 2233 2730 2238 2758
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2370 2730 2375 2758
rect 17593 2730 17598 2758
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17730 2730 17735 2758
rect 12833 2590 12838 2618
rect 12866 2590 13398 2618
rect 13426 2590 13431 2618
rect 9913 2338 9918 2366
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 10050 2338 10055 2366
rect 12441 2030 12446 2058
rect 12474 2030 13118 2058
rect 13146 2030 13151 2058
rect 2233 1946 2238 1974
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2370 1946 2375 1974
rect 17593 1946 17598 1974
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17730 1946 17735 1974
rect 10761 1806 10766 1834
rect 10794 1806 11214 1834
rect 11242 1806 11247 1834
rect 11769 1806 11774 1834
rect 11802 1806 12782 1834
rect 12810 1806 12815 1834
rect 8409 1694 8414 1722
rect 8442 1694 9030 1722
rect 9058 1694 9063 1722
rect 9913 1554 9918 1582
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 10050 1554 10055 1582
<< via3 >>
rect 2238 19194 2266 19222
rect 2290 19194 2318 19222
rect 2342 19194 2370 19222
rect 17598 19194 17626 19222
rect 17650 19194 17678 19222
rect 17702 19194 17730 19222
rect 9918 18802 9946 18830
rect 9970 18802 9998 18830
rect 10022 18802 10050 18830
rect 2238 18410 2266 18438
rect 2290 18410 2318 18438
rect 2342 18410 2370 18438
rect 17598 18410 17626 18438
rect 17650 18410 17678 18438
rect 17702 18410 17730 18438
rect 9918 18018 9946 18046
rect 9970 18018 9998 18046
rect 10022 18018 10050 18046
rect 2238 17626 2266 17654
rect 2290 17626 2318 17654
rect 2342 17626 2370 17654
rect 17598 17626 17626 17654
rect 17650 17626 17678 17654
rect 17702 17626 17730 17654
rect 9918 17234 9946 17262
rect 9970 17234 9998 17262
rect 10022 17234 10050 17262
rect 2238 16842 2266 16870
rect 2290 16842 2318 16870
rect 2342 16842 2370 16870
rect 17598 16842 17626 16870
rect 17650 16842 17678 16870
rect 17702 16842 17730 16870
rect 9918 16450 9946 16478
rect 9970 16450 9998 16478
rect 10022 16450 10050 16478
rect 2238 16058 2266 16086
rect 2290 16058 2318 16086
rect 2342 16058 2370 16086
rect 17598 16058 17626 16086
rect 17650 16058 17678 16086
rect 17702 16058 17730 16086
rect 9918 15666 9946 15694
rect 9970 15666 9998 15694
rect 10022 15666 10050 15694
rect 2238 15274 2266 15302
rect 2290 15274 2318 15302
rect 2342 15274 2370 15302
rect 17598 15274 17626 15302
rect 17650 15274 17678 15302
rect 17702 15274 17730 15302
rect 9918 14882 9946 14910
rect 9970 14882 9998 14910
rect 10022 14882 10050 14910
rect 2238 14490 2266 14518
rect 2290 14490 2318 14518
rect 2342 14490 2370 14518
rect 17598 14490 17626 14518
rect 17650 14490 17678 14518
rect 17702 14490 17730 14518
rect 9918 14098 9946 14126
rect 9970 14098 9998 14126
rect 10022 14098 10050 14126
rect 2238 13706 2266 13734
rect 2290 13706 2318 13734
rect 2342 13706 2370 13734
rect 17598 13706 17626 13734
rect 17650 13706 17678 13734
rect 17702 13706 17730 13734
rect 9918 13314 9946 13342
rect 9970 13314 9998 13342
rect 10022 13314 10050 13342
rect 2238 12922 2266 12950
rect 2290 12922 2318 12950
rect 2342 12922 2370 12950
rect 17598 12922 17626 12950
rect 17650 12922 17678 12950
rect 17702 12922 17730 12950
rect 9918 12530 9946 12558
rect 9970 12530 9998 12558
rect 10022 12530 10050 12558
rect 2238 12138 2266 12166
rect 2290 12138 2318 12166
rect 2342 12138 2370 12166
rect 17598 12138 17626 12166
rect 17650 12138 17678 12166
rect 17702 12138 17730 12166
rect 9918 11746 9946 11774
rect 9970 11746 9998 11774
rect 10022 11746 10050 11774
rect 2238 11354 2266 11382
rect 2290 11354 2318 11382
rect 2342 11354 2370 11382
rect 17598 11354 17626 11382
rect 17650 11354 17678 11382
rect 17702 11354 17730 11382
rect 9918 10962 9946 10990
rect 9970 10962 9998 10990
rect 10022 10962 10050 10990
rect 2238 10570 2266 10598
rect 2290 10570 2318 10598
rect 2342 10570 2370 10598
rect 17598 10570 17626 10598
rect 17650 10570 17678 10598
rect 17702 10570 17730 10598
rect 9918 10178 9946 10206
rect 9970 10178 9998 10206
rect 10022 10178 10050 10206
rect 2238 9786 2266 9814
rect 2290 9786 2318 9814
rect 2342 9786 2370 9814
rect 17598 9786 17626 9814
rect 17650 9786 17678 9814
rect 17702 9786 17730 9814
rect 9918 9394 9946 9422
rect 9970 9394 9998 9422
rect 10022 9394 10050 9422
rect 2238 9002 2266 9030
rect 2290 9002 2318 9030
rect 2342 9002 2370 9030
rect 17598 9002 17626 9030
rect 17650 9002 17678 9030
rect 17702 9002 17730 9030
rect 9918 8610 9946 8638
rect 9970 8610 9998 8638
rect 10022 8610 10050 8638
rect 2238 8218 2266 8246
rect 2290 8218 2318 8246
rect 2342 8218 2370 8246
rect 17598 8218 17626 8246
rect 17650 8218 17678 8246
rect 17702 8218 17730 8246
rect 9918 7826 9946 7854
rect 9970 7826 9998 7854
rect 10022 7826 10050 7854
rect 2238 7434 2266 7462
rect 2290 7434 2318 7462
rect 2342 7434 2370 7462
rect 17598 7434 17626 7462
rect 17650 7434 17678 7462
rect 17702 7434 17730 7462
rect 9918 7042 9946 7070
rect 9970 7042 9998 7070
rect 10022 7042 10050 7070
rect 2238 6650 2266 6678
rect 2290 6650 2318 6678
rect 2342 6650 2370 6678
rect 17598 6650 17626 6678
rect 17650 6650 17678 6678
rect 17702 6650 17730 6678
rect 9918 6258 9946 6286
rect 9970 6258 9998 6286
rect 10022 6258 10050 6286
rect 2238 5866 2266 5894
rect 2290 5866 2318 5894
rect 2342 5866 2370 5894
rect 17598 5866 17626 5894
rect 17650 5866 17678 5894
rect 17702 5866 17730 5894
rect 9918 5474 9946 5502
rect 9970 5474 9998 5502
rect 10022 5474 10050 5502
rect 2238 5082 2266 5110
rect 2290 5082 2318 5110
rect 2342 5082 2370 5110
rect 17598 5082 17626 5110
rect 17650 5082 17678 5110
rect 17702 5082 17730 5110
rect 9918 4690 9946 4718
rect 9970 4690 9998 4718
rect 10022 4690 10050 4718
rect 2238 4298 2266 4326
rect 2290 4298 2318 4326
rect 2342 4298 2370 4326
rect 17598 4298 17626 4326
rect 17650 4298 17678 4326
rect 17702 4298 17730 4326
rect 9918 3906 9946 3934
rect 9970 3906 9998 3934
rect 10022 3906 10050 3934
rect 2238 3514 2266 3542
rect 2290 3514 2318 3542
rect 2342 3514 2370 3542
rect 17598 3514 17626 3542
rect 17650 3514 17678 3542
rect 17702 3514 17730 3542
rect 9918 3122 9946 3150
rect 9970 3122 9998 3150
rect 10022 3122 10050 3150
rect 2238 2730 2266 2758
rect 2290 2730 2318 2758
rect 2342 2730 2370 2758
rect 17598 2730 17626 2758
rect 17650 2730 17678 2758
rect 17702 2730 17730 2758
rect 9918 2338 9946 2366
rect 9970 2338 9998 2366
rect 10022 2338 10050 2366
rect 2238 1946 2266 1974
rect 2290 1946 2318 1974
rect 2342 1946 2370 1974
rect 17598 1946 17626 1974
rect 17650 1946 17678 1974
rect 17702 1946 17730 1974
rect 9918 1554 9946 1582
rect 9970 1554 9998 1582
rect 10022 1554 10050 1582
<< metal4 >>
rect 2224 19222 2384 19238
rect 2224 19194 2238 19222
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2370 19194 2384 19222
rect 2224 18438 2384 19194
rect 2224 18410 2238 18438
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2370 18410 2384 18438
rect 2224 17654 2384 18410
rect 2224 17626 2238 17654
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2370 17626 2384 17654
rect 2224 16870 2384 17626
rect 2224 16842 2238 16870
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2370 16842 2384 16870
rect 2224 16086 2384 16842
rect 2224 16058 2238 16086
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2370 16058 2384 16086
rect 2224 15302 2384 16058
rect 2224 15274 2238 15302
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2370 15274 2384 15302
rect 2224 14518 2384 15274
rect 2224 14490 2238 14518
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2370 14490 2384 14518
rect 2224 13734 2384 14490
rect 2224 13706 2238 13734
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2370 13706 2384 13734
rect 2224 12950 2384 13706
rect 2224 12922 2238 12950
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2370 12922 2384 12950
rect 2224 12166 2384 12922
rect 2224 12138 2238 12166
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2370 12138 2384 12166
rect 2224 11382 2384 12138
rect 2224 11354 2238 11382
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2370 11354 2384 11382
rect 2224 10598 2384 11354
rect 2224 10570 2238 10598
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2370 10570 2384 10598
rect 2224 9814 2384 10570
rect 2224 9786 2238 9814
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2370 9786 2384 9814
rect 2224 9030 2384 9786
rect 2224 9002 2238 9030
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2370 9002 2384 9030
rect 2224 8246 2384 9002
rect 2224 8218 2238 8246
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2370 8218 2384 8246
rect 2224 7462 2384 8218
rect 2224 7434 2238 7462
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2370 7434 2384 7462
rect 2224 6678 2384 7434
rect 2224 6650 2238 6678
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2370 6650 2384 6678
rect 2224 5894 2384 6650
rect 2224 5866 2238 5894
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2370 5866 2384 5894
rect 2224 5110 2384 5866
rect 2224 5082 2238 5110
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2370 5082 2384 5110
rect 2224 4326 2384 5082
rect 2224 4298 2238 4326
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2370 4298 2384 4326
rect 2224 3542 2384 4298
rect 2224 3514 2238 3542
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2370 3514 2384 3542
rect 2224 2758 2384 3514
rect 2224 2730 2238 2758
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2370 2730 2384 2758
rect 2224 1974 2384 2730
rect 2224 1946 2238 1974
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2370 1946 2384 1974
rect 2224 1538 2384 1946
rect 9904 18830 10064 19238
rect 9904 18802 9918 18830
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 10050 18802 10064 18830
rect 9904 18046 10064 18802
rect 9904 18018 9918 18046
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 10050 18018 10064 18046
rect 9904 17262 10064 18018
rect 9904 17234 9918 17262
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 10050 17234 10064 17262
rect 9904 16478 10064 17234
rect 9904 16450 9918 16478
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 10050 16450 10064 16478
rect 9904 15694 10064 16450
rect 9904 15666 9918 15694
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 10050 15666 10064 15694
rect 9904 14910 10064 15666
rect 9904 14882 9918 14910
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 10050 14882 10064 14910
rect 9904 14126 10064 14882
rect 9904 14098 9918 14126
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 10050 14098 10064 14126
rect 9904 13342 10064 14098
rect 9904 13314 9918 13342
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 10050 13314 10064 13342
rect 9904 12558 10064 13314
rect 9904 12530 9918 12558
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 10050 12530 10064 12558
rect 9904 11774 10064 12530
rect 9904 11746 9918 11774
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 10050 11746 10064 11774
rect 9904 10990 10064 11746
rect 9904 10962 9918 10990
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 10050 10962 10064 10990
rect 9904 10206 10064 10962
rect 9904 10178 9918 10206
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 10050 10178 10064 10206
rect 9904 9422 10064 10178
rect 9904 9394 9918 9422
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 10050 9394 10064 9422
rect 9904 8638 10064 9394
rect 9904 8610 9918 8638
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 10050 8610 10064 8638
rect 9904 7854 10064 8610
rect 9904 7826 9918 7854
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 10050 7826 10064 7854
rect 9904 7070 10064 7826
rect 9904 7042 9918 7070
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 10050 7042 10064 7070
rect 9904 6286 10064 7042
rect 9904 6258 9918 6286
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 10050 6258 10064 6286
rect 9904 5502 10064 6258
rect 9904 5474 9918 5502
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 10050 5474 10064 5502
rect 9904 4718 10064 5474
rect 9904 4690 9918 4718
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 10050 4690 10064 4718
rect 9904 3934 10064 4690
rect 9904 3906 9918 3934
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 10050 3906 10064 3934
rect 9904 3150 10064 3906
rect 9904 3122 9918 3150
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 10050 3122 10064 3150
rect 9904 2366 10064 3122
rect 9904 2338 9918 2366
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 10050 2338 10064 2366
rect 9904 1582 10064 2338
rect 9904 1554 9918 1582
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 10050 1554 10064 1582
rect 9904 1538 10064 1554
rect 17584 19222 17744 19238
rect 17584 19194 17598 19222
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17730 19194 17744 19222
rect 17584 18438 17744 19194
rect 17584 18410 17598 18438
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17730 18410 17744 18438
rect 17584 17654 17744 18410
rect 17584 17626 17598 17654
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17730 17626 17744 17654
rect 17584 16870 17744 17626
rect 17584 16842 17598 16870
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17730 16842 17744 16870
rect 17584 16086 17744 16842
rect 17584 16058 17598 16086
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17730 16058 17744 16086
rect 17584 15302 17744 16058
rect 17584 15274 17598 15302
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17730 15274 17744 15302
rect 17584 14518 17744 15274
rect 17584 14490 17598 14518
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17730 14490 17744 14518
rect 17584 13734 17744 14490
rect 17584 13706 17598 13734
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17730 13706 17744 13734
rect 17584 12950 17744 13706
rect 17584 12922 17598 12950
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17730 12922 17744 12950
rect 17584 12166 17744 12922
rect 17584 12138 17598 12166
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17730 12138 17744 12166
rect 17584 11382 17744 12138
rect 17584 11354 17598 11382
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17730 11354 17744 11382
rect 17584 10598 17744 11354
rect 17584 10570 17598 10598
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17730 10570 17744 10598
rect 17584 9814 17744 10570
rect 17584 9786 17598 9814
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17730 9786 17744 9814
rect 17584 9030 17744 9786
rect 17584 9002 17598 9030
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17730 9002 17744 9030
rect 17584 8246 17744 9002
rect 17584 8218 17598 8246
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17730 8218 17744 8246
rect 17584 7462 17744 8218
rect 17584 7434 17598 7462
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17730 7434 17744 7462
rect 17584 6678 17744 7434
rect 17584 6650 17598 6678
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17730 6650 17744 6678
rect 17584 5894 17744 6650
rect 17584 5866 17598 5894
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17730 5866 17744 5894
rect 17584 5110 17744 5866
rect 17584 5082 17598 5110
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17730 5082 17744 5110
rect 17584 4326 17744 5082
rect 17584 4298 17598 4326
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17730 4298 17744 4326
rect 17584 3542 17744 4298
rect 17584 3514 17598 3542
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17730 3514 17744 3542
rect 17584 2758 17744 3514
rect 17584 2730 17598 2758
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17730 2730 17744 2758
rect 17584 1974 17744 2730
rect 17584 1946 17598 1974
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17730 1946 17744 1974
rect 17584 1538 17744 1946
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _118_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9632 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _119_
timestamp 1698175906
transform -1 0 10472 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _120_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9856 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _121_
timestamp 1698175906
transform -1 0 10752 0 -1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _122_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8792 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _123_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 12880 0 -1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _124_
timestamp 1698175906
transform -1 0 9800 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _125_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9016 0 1 9408
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _126_
timestamp 1698175906
transform -1 0 11704 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _127_
timestamp 1698175906
transform 1 0 11144 0 1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _128_
timestamp 1698175906
transform 1 0 11424 0 -1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _129_
timestamp 1698175906
transform 1 0 11592 0 1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _130_
timestamp 1698175906
transform -1 0 10360 0 -1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _131_
timestamp 1698175906
transform 1 0 11480 0 1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _132_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 11872 0 -1 7840
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _133_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 11480 0 -1 7840
box -43 -43 659 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _134_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9408 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _135_
timestamp 1698175906
transform 1 0 10080 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _136_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 10920 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _137_
timestamp 1698175906
transform -1 0 11312 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _138_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 11312 0 1 8624
box -43 -43 771 435
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _139_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 12992 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _140_
timestamp 1698175906
transform -1 0 10304 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _141_
timestamp 1698175906
transform 1 0 13216 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _142_
timestamp 1698175906
transform -1 0 13216 0 -1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _143_
timestamp 1698175906
transform -1 0 9296 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _144_
timestamp 1698175906
transform -1 0 8512 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _145_
timestamp 1698175906
transform 1 0 8120 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _146_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 12936 0 1 8624
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _147_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 14952 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _148_
timestamp 1698175906
transform -1 0 13720 0 1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _149_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 12152 0 -1 10192
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _150_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 13776 0 -1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _151_
timestamp 1698175906
transform 1 0 14952 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _152_
timestamp 1698175906
transform 1 0 10920 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _153_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 11088 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _154_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 14336 0 1 8624
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _155_
timestamp 1698175906
transform 1 0 14504 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _156_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 9464 0 1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _157_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8120 0 1 7840
box -43 -43 715 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _158_
timestamp 1698175906
transform 1 0 8624 0 -1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _159_
timestamp 1698175906
transform 1 0 9016 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _160_
timestamp 1698175906
transform 1 0 8288 0 1 12544
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _161_
timestamp 1698175906
transform -1 0 10920 0 1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _162_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 10304 0 1 9408
box -43 -43 771 435
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _163_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 10248 0 1 10192
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _164_
timestamp 1698175906
transform 1 0 9520 0 1 11760
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _165_
timestamp 1698175906
transform 1 0 9352 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _166_
timestamp 1698175906
transform 1 0 9688 0 -1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _167_
timestamp 1698175906
transform 1 0 10584 0 -1 10192
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _168_
timestamp 1698175906
transform 1 0 10752 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _169_
timestamp 1698175906
transform 1 0 11424 0 -1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _170_
timestamp 1698175906
transform -1 0 9632 0 -1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _171_
timestamp 1698175906
transform 1 0 11480 0 1 9408
box -43 -43 771 435
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _172_
timestamp 1698175906
transform -1 0 9688 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _173_
timestamp 1698175906
transform 1 0 8792 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _174_
timestamp 1698175906
transform 1 0 8568 0 1 8624
box -43 -43 771 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _175_
timestamp 1698175906
transform -1 0 7560 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _176_
timestamp 1698175906
transform 1 0 8624 0 -1 9408
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _177_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 7336 0 1 8624
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _178_
timestamp 1698175906
transform -1 0 9016 0 1 9408
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _179_
timestamp 1698175906
transform 1 0 6216 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _180_
timestamp 1698175906
transform 1 0 11536 0 -1 9408
box -43 -43 771 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _181_
timestamp 1698175906
transform -1 0 12376 0 -1 12544
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _182_
timestamp 1698175906
transform 1 0 11200 0 1 13328
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _183_
timestamp 1698175906
transform -1 0 11592 0 1 12544
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _184_
timestamp 1698175906
transform 1 0 13496 0 1 8624
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _185_
timestamp 1698175906
transform 1 0 14000 0 1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _186_
timestamp 1698175906
transform 1 0 13496 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _187_
timestamp 1698175906
transform -1 0 10472 0 1 10976
box -43 -43 771 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _188_
timestamp 1698175906
transform 1 0 12320 0 1 12544
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _189_
timestamp 1698175906
transform 1 0 12544 0 -1 14112
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _190_
timestamp 1698175906
transform 1 0 13720 0 1 12544
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _191_
timestamp 1698175906
transform -1 0 14168 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _192_
timestamp 1698175906
transform -1 0 7840 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _193_
timestamp 1698175906
transform -1 0 8120 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _194_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 7840 0 -1 8624
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _195_
timestamp 1698175906
transform -1 0 7616 0 1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _196_
timestamp 1698175906
transform -1 0 10528 0 -1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _197_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9688 0 1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _198_
timestamp 1698175906
transform 1 0 9632 0 -1 13328
box -43 -43 659 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _199_
timestamp 1698175906
transform 1 0 8344 0 1 10192
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _200_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 6664 0 1 10192
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _201_
timestamp 1698175906
transform -1 0 6328 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _202_
timestamp 1698175906
transform -1 0 7000 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _203_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 7112 0 -1 9408
box -43 -43 883 435
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _204_
timestamp 1698175906
transform -1 0 6552 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _205_
timestamp 1698175906
transform 1 0 13216 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _206_
timestamp 1698175906
transform -1 0 13216 0 -1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _207_
timestamp 1698175906
transform 1 0 10080 0 1 7840
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _208_
timestamp 1698175906
transform 1 0 10584 0 1 7840
box -43 -43 659 435
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _209_
timestamp 1698175906
transform 1 0 12544 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _210_
timestamp 1698175906
transform -1 0 12768 0 1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _211_
timestamp 1698175906
transform -1 0 8064 0 1 13328
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _212_
timestamp 1698175906
transform -1 0 7672 0 1 13328
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _213_
timestamp 1698175906
transform -1 0 13832 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _214_
timestamp 1698175906
transform 1 0 12768 0 1 12544
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _215_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10584 0 1 10976
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _216_
timestamp 1698175906
transform -1 0 13944 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _217_
timestamp 1698175906
transform 1 0 13944 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _218_
timestamp 1698175906
transform 1 0 8960 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _219_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 9072 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _220_
timestamp 1698175906
transform 1 0 8624 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _221_
timestamp 1698175906
transform -1 0 7504 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _222_
timestamp 1698175906
transform 1 0 6664 0 1 10976
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _223_
timestamp 1698175906
transform 1 0 7504 0 -1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _224_
timestamp 1698175906
transform -1 0 7840 0 -1 13328
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _225_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 7672 0 -1 12544
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _226_
timestamp 1698175906
transform 1 0 8960 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _227_
timestamp 1698175906
transform 1 0 11088 0 -1 8624
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _228_
timestamp 1698175906
transform 1 0 11704 0 1 8624
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _229_
timestamp 1698175906
transform 1 0 11984 0 -1 7056
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _230_
timestamp 1698175906
transform 1 0 11368 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _231_
timestamp 1698175906
transform 1 0 13776 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _232_
timestamp 1698175906
transform 1 0 12768 0 1 10976
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _233_
timestamp 1698175906
transform 1 0 13328 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _234_
timestamp 1698175906
transform 1 0 12544 0 -1 7056
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _235_
timestamp 1698175906
transform 1 0 11928 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _236_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10248 0 -1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _237_
timestamp 1698175906
transform 1 0 13776 0 -1 8624
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _238_
timestamp 1698175906
transform 1 0 13944 0 -1 7840
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _239_
timestamp 1698175906
transform 1 0 6720 0 -1 10192
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _240_
timestamp 1698175906
transform 1 0 8008 0 1 6272
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _241_
timestamp 1698175906
transform 1 0 9408 0 -1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _242_
timestamp 1698175906
transform 1 0 11144 0 1 10976
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _243_
timestamp 1698175906
transform 1 0 8064 0 1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _244_
timestamp 1698175906
transform -1 0 7112 0 -1 8624
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _245_
timestamp 1698175906
transform 1 0 10696 0 -1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _246_
timestamp 1698175906
transform 1 0 13944 0 -1 10976
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _247_
timestamp 1698175906
transform 1 0 11592 0 1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _248_
timestamp 1698175906
transform 1 0 13496 0 -1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _249_
timestamp 1698175906
transform 1 0 6664 0 -1 7840
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _250_
timestamp 1698175906
transform 1 0 8904 0 -1 14112
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _251_
timestamp 1698175906
transform -1 0 6552 0 1 10192
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _252_
timestamp 1698175906
transform -1 0 6496 0 1 9408
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _253_
timestamp 1698175906
transform 1 0 12992 0 -1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _254_
timestamp 1698175906
transform 1 0 9240 0 -1 7840
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _255_
timestamp 1698175906
transform 1 0 6552 0 -1 14112
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _256_
timestamp 1698175906
transform 1 0 12712 0 -1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _257_
timestamp 1698175906
transform 1 0 13944 0 -1 9408
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _258_
timestamp 1698175906
transform -1 0 9240 0 1 10976
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _259_
timestamp 1698175906
transform -1 0 7056 0 -1 11760
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _260_
timestamp 1698175906
transform -1 0 8288 0 1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _261_
timestamp 1698175906
transform 1 0 11032 0 1 6272
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _262_
timestamp 1698175906
transform 1 0 13272 0 -1 11760
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _263_
timestamp 1698175906
transform 1 0 11816 0 1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _264_
timestamp 1698175906
transform -1 0 7168 0 1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _265_
timestamp 1698175906
transform 1 0 8176 0 -1 14112
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__236__CLK dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 11984 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__237__CLK
timestamp 1698175906
transform 1 0 15512 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__238__CLK
timestamp 1698175906
transform 1 0 15680 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__239__CLK
timestamp 1698175906
transform 1 0 8344 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__240__CLK
timestamp 1698175906
transform -1 0 9856 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__241__CLK
timestamp 1698175906
transform 1 0 11144 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__242__CLK
timestamp 1698175906
transform 1 0 13160 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__243__CLK
timestamp 1698175906
transform 1 0 10248 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__244__CLK
timestamp 1698175906
transform 1 0 7224 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__245__CLK
timestamp 1698175906
transform 1 0 12208 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__246__CLK
timestamp 1698175906
transform 1 0 15680 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__247__CLK
timestamp 1698175906
transform 1 0 13328 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__248__CLK
timestamp 1698175906
transform 1 0 15232 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__249__CLK
timestamp 1698175906
transform 1 0 8400 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__250__CLK
timestamp 1698175906
transform 1 0 10640 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__251__CLK
timestamp 1698175906
transform 1 0 6552 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__252__CLK
timestamp 1698175906
transform 1 0 6664 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__253__CLK
timestamp 1698175906
transform 1 0 14728 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__254__CLK
timestamp 1698175906
transform 1 0 10864 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__255__CLK
timestamp 1698175906
transform -1 0 8288 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__256__CLK
timestamp 1698175906
transform 1 0 14448 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__257__CLK
timestamp 1698175906
transform 1 0 15680 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__258__CLK
timestamp 1698175906
transform 1 0 9520 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__259__CLK
timestamp 1698175906
transform 1 0 7280 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__260__CLK
timestamp 1698175906
transform 1 0 8736 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__261__CLK
timestamp 1698175906
transform 1 0 12768 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__262__CLK
timestamp 1698175906
transform 1 0 15008 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__263__CLK
timestamp 1698175906
transform 1 0 13552 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1698175906
transform -1 0 10472 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10584 0 1 10192
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1698175906
transform -1 0 11424 0 -1 10976
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1698175906
transform 1 0 12544 0 -1 10192
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 784 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698175906
transform 1 0 2688 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698175906
transform 1 0 4592 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698175906
transform 1 0 6496 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_138 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8400 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_165 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9912 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_169
timestamp 1698175906
transform 1 0 10136 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_172
timestamp 1698175906
transform 1 0 10304 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_176 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10528 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_232
timestamp 1698175906
transform 1 0 13664 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_236
timestamp 1698175906
transform 1 0 13888 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_240
timestamp 1698175906
transform 1 0 14112 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_274
timestamp 1698175906
transform 1 0 16016 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_308
timestamp 1698175906
transform 1 0 17920 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_342
timestamp 1698175906
transform 1 0 19824 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_346
timestamp 1698175906
transform 1 0 20048 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_348
timestamp 1698175906
transform 1 0 20160 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 784 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698175906
transform 1 0 4368 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698175906
transform 1 0 4704 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698175906
transform 1 0 8288 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_142
timestamp 1698175906
transform 1 0 8624 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_206
timestamp 1698175906
transform 1 0 12208 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_238
timestamp 1698175906
transform 1 0 14000 0 -1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_270 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 15792 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_278
timestamp 1698175906
transform 1 0 16240 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_282
timestamp 1698175906
transform 1 0 16464 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_346
timestamp 1698175906
transform 1 0 20048 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_348
timestamp 1698175906
transform 1 0 20160 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698175906
transform 1 0 784 0 1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698175906
transform 1 0 2576 0 1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698175906
transform 1 0 2744 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698175906
transform 1 0 6328 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_107
timestamp 1698175906
transform 1 0 6664 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_171
timestamp 1698175906
transform 1 0 10248 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_177
timestamp 1698175906
transform 1 0 10584 0 1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_209
timestamp 1698175906
transform 1 0 12376 0 1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_243
timestamp 1698175906
transform 1 0 14280 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698175906
transform 1 0 14504 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698175906
transform 1 0 18088 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_317
timestamp 1698175906
transform 1 0 18424 0 1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698175906
transform 1 0 784 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698175906
transform 1 0 4368 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698175906
transform 1 0 4704 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698175906
transform 1 0 8288 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_142
timestamp 1698175906
transform 1 0 8624 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_206
timestamp 1698175906
transform 1 0 12208 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_212
timestamp 1698175906
transform 1 0 12544 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_276
timestamp 1698175906
transform 1 0 16128 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_282
timestamp 1698175906
transform 1 0 16464 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_346
timestamp 1698175906
transform 1 0 20048 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_348
timestamp 1698175906
transform 1 0 20160 0 -1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698175906
transform 1 0 784 0 1 3136
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698175906
transform 1 0 2576 0 1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698175906
transform 1 0 2744 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698175906
transform 1 0 6328 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_107
timestamp 1698175906
transform 1 0 6664 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698175906
transform 1 0 10248 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_177
timestamp 1698175906
transform 1 0 10584 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_241
timestamp 1698175906
transform 1 0 14168 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698175906
transform 1 0 14504 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698175906
transform 1 0 18088 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_317
timestamp 1698175906
transform 1 0 18424 0 1 3136
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698175906
transform 1 0 784 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698175906
transform 1 0 4368 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698175906
transform 1 0 4704 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698175906
transform 1 0 8288 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_142
timestamp 1698175906
transform 1 0 8624 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_206
timestamp 1698175906
transform 1 0 12208 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_212
timestamp 1698175906
transform 1 0 12544 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698175906
transform 1 0 16128 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_282
timestamp 1698175906
transform 1 0 16464 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_346
timestamp 1698175906
transform 1 0 20048 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_348
timestamp 1698175906
transform 1 0 20160 0 -1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698175906
transform 1 0 784 0 1 3920
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698175906
transform 1 0 2576 0 1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698175906
transform 1 0 2744 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698175906
transform 1 0 6328 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_107
timestamp 1698175906
transform 1 0 6664 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_171
timestamp 1698175906
transform 1 0 10248 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_177
timestamp 1698175906
transform 1 0 10584 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_241
timestamp 1698175906
transform 1 0 14168 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_247
timestamp 1698175906
transform 1 0 14504 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_311
timestamp 1698175906
transform 1 0 18088 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_317
timestamp 1698175906
transform 1 0 18424 0 1 3920
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698175906
transform 1 0 784 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698175906
transform 1 0 4368 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_72
timestamp 1698175906
transform 1 0 4704 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698175906
transform 1 0 8288 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_142
timestamp 1698175906
transform 1 0 8624 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_206
timestamp 1698175906
transform 1 0 12208 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_212
timestamp 1698175906
transform 1 0 12544 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_276
timestamp 1698175906
transform 1 0 16128 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_282
timestamp 1698175906
transform 1 0 16464 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_346
timestamp 1698175906
transform 1 0 20048 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_348
timestamp 1698175906
transform 1 0 20160 0 -1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698175906
transform 1 0 784 0 1 4704
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698175906
transform 1 0 2576 0 1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_37
timestamp 1698175906
transform 1 0 2744 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_101
timestamp 1698175906
transform 1 0 6328 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_107
timestamp 1698175906
transform 1 0 6664 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_171
timestamp 1698175906
transform 1 0 10248 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_177
timestamp 1698175906
transform 1 0 10584 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_241
timestamp 1698175906
transform 1 0 14168 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_247
timestamp 1698175906
transform 1 0 14504 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_311
timestamp 1698175906
transform 1 0 18088 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_317
timestamp 1698175906
transform 1 0 18424 0 1 4704
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698175906
transform 1 0 784 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698175906
transform 1 0 4368 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_72
timestamp 1698175906
transform 1 0 4704 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_136
timestamp 1698175906
transform 1 0 8288 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_142
timestamp 1698175906
transform 1 0 8624 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_206
timestamp 1698175906
transform 1 0 12208 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_212
timestamp 1698175906
transform 1 0 12544 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_276
timestamp 1698175906
transform 1 0 16128 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_282
timestamp 1698175906
transform 1 0 16464 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_346
timestamp 1698175906
transform 1 0 20048 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_348
timestamp 1698175906
transform 1 0 20160 0 -1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698175906
transform 1 0 784 0 1 5488
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698175906
transform 1 0 2576 0 1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_37
timestamp 1698175906
transform 1 0 2744 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698175906
transform 1 0 6328 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_107
timestamp 1698175906
transform 1 0 6664 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_171
timestamp 1698175906
transform 1 0 10248 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_177
timestamp 1698175906
transform 1 0 10584 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_241
timestamp 1698175906
transform 1 0 14168 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_247
timestamp 1698175906
transform 1 0 14504 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_311
timestamp 1698175906
transform 1 0 18088 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_317
timestamp 1698175906
transform 1 0 18424 0 1 5488
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2
timestamp 1698175906
transform 1 0 784 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698175906
transform 1 0 4368 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_72
timestamp 1698175906
transform 1 0 4704 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698175906
transform 1 0 8288 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_11_142
timestamp 1698175906
transform 1 0 8624 0 -1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_174 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10416 0 -1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_190
timestamp 1698175906
transform 1 0 11312 0 -1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_198
timestamp 1698175906
transform 1 0 11760 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_202
timestamp 1698175906
transform 1 0 11984 0 -1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_212
timestamp 1698175906
transform 1 0 12544 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_276
timestamp 1698175906
transform 1 0 16128 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_282
timestamp 1698175906
transform 1 0 16464 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_346
timestamp 1698175906
transform 1 0 20048 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_348
timestamp 1698175906
transform 1 0 20160 0 -1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698175906
transform 1 0 784 0 1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698175906
transform 1 0 2576 0 1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_37
timestamp 1698175906
transform 1 0 2744 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698175906
transform 1 0 6328 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_107
timestamp 1698175906
transform 1 0 6664 0 1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_123
timestamp 1698175906
transform 1 0 7560 0 1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_160
timestamp 1698175906
transform 1 0 9632 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_164
timestamp 1698175906
transform 1 0 9856 0 1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_172
timestamp 1698175906
transform 1 0 10304 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_174
timestamp 1698175906
transform 1 0 10416 0 1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_177
timestamp 1698175906
transform 1 0 10584 0 1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_214
timestamp 1698175906
transform 1 0 12656 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_218
timestamp 1698175906
transform 1 0 12880 0 1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_234
timestamp 1698175906
transform 1 0 13776 0 1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_242
timestamp 1698175906
transform 1 0 14224 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_244
timestamp 1698175906
transform 1 0 14336 0 1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_247
timestamp 1698175906
transform 1 0 14504 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_311
timestamp 1698175906
transform 1 0 18088 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_317
timestamp 1698175906
transform 1 0 18424 0 1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_2
timestamp 1698175906
transform 1 0 784 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_66
timestamp 1698175906
transform 1 0 4368 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_72
timestamp 1698175906
transform 1 0 4704 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_136
timestamp 1698175906
transform 1 0 8288 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_142
timestamp 1698175906
transform 1 0 8624 0 -1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_158
timestamp 1698175906
transform 1 0 9520 0 -1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_166
timestamp 1698175906
transform 1 0 9968 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_170
timestamp 1698175906
transform 1 0 10192 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_200
timestamp 1698175906
transform 1 0 11872 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_209
timestamp 1698175906
transform 1 0 12376 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_219
timestamp 1698175906
transform 1 0 12936 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_249
timestamp 1698175906
transform 1 0 14616 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_253
timestamp 1698175906
transform 1 0 14840 0 -1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_269
timestamp 1698175906
transform 1 0 15736 0 -1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_277
timestamp 1698175906
transform 1 0 16184 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_279
timestamp 1698175906
transform 1 0 16296 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_282
timestamp 1698175906
transform 1 0 16464 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_346
timestamp 1698175906
transform 1 0 20048 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_348
timestamp 1698175906
transform 1 0 20160 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698175906
transform 1 0 784 0 1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698175906
transform 1 0 2576 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_37
timestamp 1698175906
transform 1 0 2744 0 1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_101
timestamp 1698175906
transform 1 0 6328 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_107
timestamp 1698175906
transform 1 0 6664 0 1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_139
timestamp 1698175906
transform 1 0 8456 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_147
timestamp 1698175906
transform 1 0 8904 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_156
timestamp 1698175906
transform 1 0 9408 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_172
timestamp 1698175906
transform 1 0 10304 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_174
timestamp 1698175906
transform 1 0 10416 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_177
timestamp 1698175906
transform 1 0 10584 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_181
timestamp 1698175906
transform 1 0 10808 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_184
timestamp 1698175906
transform 1 0 10976 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_188
timestamp 1698175906
transform 1 0 11200 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_190
timestamp 1698175906
transform 1 0 11312 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_228
timestamp 1698175906
transform 1 0 13440 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_232
timestamp 1698175906
transform 1 0 13664 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_240
timestamp 1698175906
transform 1 0 14112 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_244
timestamp 1698175906
transform 1 0 14336 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_247
timestamp 1698175906
transform 1 0 14504 0 1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_311
timestamp 1698175906
transform 1 0 18088 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_317
timestamp 1698175906
transform 1 0 18424 0 1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_2
timestamp 1698175906
transform 1 0 784 0 -1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_66
timestamp 1698175906
transform 1 0 4368 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_72
timestamp 1698175906
transform 1 0 4704 0 -1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_104
timestamp 1698175906
transform 1 0 6496 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_106
timestamp 1698175906
transform 1 0 6608 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_136
timestamp 1698175906
transform 1 0 8288 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_148
timestamp 1698175906
transform 1 0 8960 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_152
timestamp 1698175906
transform 1 0 9184 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_200
timestamp 1698175906
transform 1 0 11872 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_209
timestamp 1698175906
transform 1 0 12376 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_212
timestamp 1698175906
transform 1 0 12544 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_216
timestamp 1698175906
transform 1 0 12768 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_232
timestamp 1698175906
transform 1 0 13664 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_236
timestamp 1698175906
transform 1 0 13888 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_266
timestamp 1698175906
transform 1 0 15568 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_270
timestamp 1698175906
transform 1 0 15792 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_278
timestamp 1698175906
transform 1 0 16240 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_282
timestamp 1698175906
transform 1 0 16464 0 -1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_314
timestamp 1698175906
transform 1 0 18256 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_322
timestamp 1698175906
transform 1 0 18704 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_2
timestamp 1698175906
transform 1 0 784 0 1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698175906
transform 1 0 2576 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_37
timestamp 1698175906
transform 1 0 2744 0 1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_101
timestamp 1698175906
transform 1 0 6328 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_107
timestamp 1698175906
transform 1 0 6664 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_115
timestamp 1698175906
transform 1 0 7112 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_117
timestamp 1698175906
transform 1 0 7224 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_124
timestamp 1698175906
transform 1 0 7616 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_132
timestamp 1698175906
transform 1 0 8064 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_145
timestamp 1698175906
transform 1 0 8792 0 1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_161
timestamp 1698175906
transform 1 0 9688 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_165
timestamp 1698175906
transform 1 0 9912 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_167
timestamp 1698175906
transform 1 0 10024 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_188
timestamp 1698175906
transform 1 0 11200 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_192
timestamp 1698175906
transform 1 0 11424 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_194
timestamp 1698175906
transform 1 0 11536 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_201
timestamp 1698175906
transform 1 0 11928 0 1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_233
timestamp 1698175906
transform 1 0 13720 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_241
timestamp 1698175906
transform 1 0 14168 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_247
timestamp 1698175906
transform 1 0 14504 0 1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_311
timestamp 1698175906
transform 1 0 18088 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_317
timestamp 1698175906
transform 1 0 18424 0 1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_2
timestamp 1698175906
transform 1 0 784 0 -1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_66
timestamp 1698175906
transform 1 0 4368 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_72
timestamp 1698175906
transform 1 0 4704 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_80
timestamp 1698175906
transform 1 0 5152 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_84
timestamp 1698175906
transform 1 0 5376 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_115
timestamp 1698175906
transform 1 0 7112 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_119
timestamp 1698175906
transform 1 0 7336 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_138
timestamp 1698175906
transform 1 0 8400 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_142
timestamp 1698175906
transform 1 0 8624 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_154
timestamp 1698175906
transform 1 0 9296 0 -1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_191
timestamp 1698175906
transform 1 0 11368 0 -1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_207
timestamp 1698175906
transform 1 0 12264 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_209
timestamp 1698175906
transform 1 0 12376 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_212
timestamp 1698175906
transform 1 0 12544 0 -1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_228
timestamp 1698175906
transform 1 0 13440 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_232
timestamp 1698175906
transform 1 0 13664 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_263
timestamp 1698175906
transform 1 0 15400 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_267
timestamp 1698175906
transform 1 0 15624 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_275
timestamp 1698175906
transform 1 0 16072 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_279
timestamp 1698175906
transform 1 0 16296 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_282
timestamp 1698175906
transform 1 0 16464 0 -1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_314
timestamp 1698175906
transform 1 0 18256 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_322
timestamp 1698175906
transform 1 0 18704 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_28
timestamp 1698175906
transform 1 0 2240 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_32
timestamp 1698175906
transform 1 0 2464 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698175906
transform 1 0 2576 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_37
timestamp 1698175906
transform 1 0 2744 0 1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_69
timestamp 1698175906
transform 1 0 4536 0 1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_85
timestamp 1698175906
transform 1 0 5432 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_93
timestamp 1698175906
transform 1 0 5880 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_97
timestamp 1698175906
transform 1 0 6104 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_107
timestamp 1698175906
transform 1 0 6664 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_109
timestamp 1698175906
transform 1 0 6776 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_123
timestamp 1698175906
transform 1 0 7560 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_154
timestamp 1698175906
transform 1 0 9296 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_161
timestamp 1698175906
transform 1 0 9688 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_190
timestamp 1698175906
transform 1 0 11312 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_207
timestamp 1698175906
transform 1 0 12264 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_215
timestamp 1698175906
transform 1 0 12712 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_244
timestamp 1698175906
transform 1 0 14336 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_263
timestamp 1698175906
transform 1 0 15400 0 1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_295
timestamp 1698175906
transform 1 0 17192 0 1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_311
timestamp 1698175906
transform 1 0 18088 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_317
timestamp 1698175906
transform 1 0 18424 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_321
timestamp 1698175906
transform 1 0 18648 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_2
timestamp 1698175906
transform 1 0 784 0 -1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_66
timestamp 1698175906
transform 1 0 4368 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_72
timestamp 1698175906
transform 1 0 4704 0 -1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_88
timestamp 1698175906
transform 1 0 5600 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_96
timestamp 1698175906
transform 1 0 6048 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_105
timestamp 1698175906
transform 1 0 6552 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_109
timestamp 1698175906
transform 1 0 6776 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_113
timestamp 1698175906
transform 1 0 7000 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_130
timestamp 1698175906
transform 1 0 7952 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_166
timestamp 1698175906
transform 1 0 9968 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_174
timestamp 1698175906
transform 1 0 10416 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_182
timestamp 1698175906
transform 1 0 10864 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_207
timestamp 1698175906
transform 1 0 12264 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_209
timestamp 1698175906
transform 1 0 12376 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_212
timestamp 1698175906
transform 1 0 12544 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_216
timestamp 1698175906
transform 1 0 12768 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_234
timestamp 1698175906
transform 1 0 13776 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_236
timestamp 1698175906
transform 1 0 13888 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_266
timestamp 1698175906
transform 1 0 15568 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_270
timestamp 1698175906
transform 1 0 15792 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_278
timestamp 1698175906
transform 1 0 16240 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_282
timestamp 1698175906
transform 1 0 16464 0 -1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_346
timestamp 1698175906
transform 1 0 20048 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_348
timestamp 1698175906
transform 1 0 20160 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_2
timestamp 1698175906
transform 1 0 784 0 1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698175906
transform 1 0 2576 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_37
timestamp 1698175906
transform 1 0 2744 0 1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_69
timestamp 1698175906
transform 1 0 4536 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_73
timestamp 1698175906
transform 1 0 4760 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_104
timestamp 1698175906
transform 1 0 6496 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_113
timestamp 1698175906
transform 1 0 7000 0 1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_129
timestamp 1698175906
transform 1 0 7896 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_139
timestamp 1698175906
transform 1 0 8456 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_143
timestamp 1698175906
transform 1 0 8680 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_158
timestamp 1698175906
transform 1 0 9520 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_172
timestamp 1698175906
transform 1 0 10304 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_174
timestamp 1698175906
transform 1 0 10416 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_189
timestamp 1698175906
transform 1 0 11256 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_206
timestamp 1698175906
transform 1 0 12208 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_210
timestamp 1698175906
transform 1 0 12432 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_228
timestamp 1698175906
transform 1 0 13440 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_253
timestamp 1698175906
transform 1 0 14840 0 1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_285
timestamp 1698175906
transform 1 0 16632 0 1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_301
timestamp 1698175906
transform 1 0 17528 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_309
timestamp 1698175906
transform 1 0 17976 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_313
timestamp 1698175906
transform 1 0 18200 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_317
timestamp 1698175906
transform 1 0 18424 0 1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_28
timestamp 1698175906
transform 1 0 2240 0 -1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_60
timestamp 1698175906
transform 1 0 4032 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_68
timestamp 1698175906
transform 1 0 4480 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_72
timestamp 1698175906
transform 1 0 4704 0 -1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_88
timestamp 1698175906
transform 1 0 5600 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_92
timestamp 1698175906
transform 1 0 5824 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_94
timestamp 1698175906
transform 1 0 5936 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_101
timestamp 1698175906
transform 1 0 6328 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_107
timestamp 1698175906
transform 1 0 6664 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_137
timestamp 1698175906
transform 1 0 8344 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_139
timestamp 1698175906
transform 1 0 8456 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_142
timestamp 1698175906
transform 1 0 8624 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_144
timestamp 1698175906
transform 1 0 8736 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_163
timestamp 1698175906
transform 1 0 9800 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_172
timestamp 1698175906
transform 1 0 10304 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_176
timestamp 1698175906
transform 1 0 10528 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_190
timestamp 1698175906
transform 1 0 11312 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_198
timestamp 1698175906
transform 1 0 11760 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_202
timestamp 1698175906
transform 1 0 11984 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_204
timestamp 1698175906
transform 1 0 12096 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_262
timestamp 1698175906
transform 1 0 15344 0 -1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_278
timestamp 1698175906
transform 1 0 16240 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_282
timestamp 1698175906
transform 1 0 16464 0 -1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_346
timestamp 1698175906
transform 1 0 20048 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_348
timestamp 1698175906
transform 1 0 20160 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_2
timestamp 1698175906
transform 1 0 784 0 1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698175906
transform 1 0 2576 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_37
timestamp 1698175906
transform 1 0 2744 0 1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_69
timestamp 1698175906
transform 1 0 4536 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_73
timestamp 1698175906
transform 1 0 4760 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_75
timestamp 1698175906
transform 1 0 4872 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_117
timestamp 1698175906
transform 1 0 7224 0 1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_133
timestamp 1698175906
transform 1 0 8120 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_150
timestamp 1698175906
transform 1 0 9072 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_171
timestamp 1698175906
transform 1 0 10248 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_233
timestamp 1698175906
transform 1 0 13720 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_237
timestamp 1698175906
transform 1 0 13944 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_244
timestamp 1698175906
transform 1 0 14336 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_247
timestamp 1698175906
transform 1 0 14504 0 1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_311
timestamp 1698175906
transform 1 0 18088 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_317
timestamp 1698175906
transform 1 0 18424 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_321
timestamp 1698175906
transform 1 0 18648 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_28
timestamp 1698175906
transform 1 0 2240 0 -1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_60
timestamp 1698175906
transform 1 0 4032 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_68
timestamp 1698175906
transform 1 0 4480 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_72
timestamp 1698175906
transform 1 0 4704 0 -1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_136
timestamp 1698175906
transform 1 0 8288 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_198
timestamp 1698175906
transform 1 0 11760 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_206
timestamp 1698175906
transform 1 0 12208 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_228
timestamp 1698175906
transform 1 0 13440 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_266
timestamp 1698175906
transform 1 0 15568 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_270
timestamp 1698175906
transform 1 0 15792 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_278
timestamp 1698175906
transform 1 0 16240 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_282
timestamp 1698175906
transform 1 0 16464 0 -1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_346
timestamp 1698175906
transform 1 0 20048 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_348
timestamp 1698175906
transform 1 0 20160 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_2
timestamp 1698175906
transform 1 0 784 0 1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698175906
transform 1 0 2576 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_37
timestamp 1698175906
transform 1 0 2744 0 1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_101
timestamp 1698175906
transform 1 0 6328 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_117
timestamp 1698175906
transform 1 0 7224 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_121
timestamp 1698175906
transform 1 0 7448 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_123
timestamp 1698175906
transform 1 0 7560 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_161
timestamp 1698175906
transform 1 0 9688 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_221
timestamp 1698175906
transform 1 0 13048 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_225
timestamp 1698175906
transform 1 0 13272 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_240
timestamp 1698175906
transform 1 0 14112 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_244
timestamp 1698175906
transform 1 0 14336 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_247
timestamp 1698175906
transform 1 0 14504 0 1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_311
timestamp 1698175906
transform 1 0 18088 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_317
timestamp 1698175906
transform 1 0 18424 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_321
timestamp 1698175906
transform 1 0 18648 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_28
timestamp 1698175906
transform 1 0 2240 0 -1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_60
timestamp 1698175906
transform 1 0 4032 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_68
timestamp 1698175906
transform 1 0 4480 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_72
timestamp 1698175906
transform 1 0 4704 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_80
timestamp 1698175906
transform 1 0 5152 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_84
timestamp 1698175906
transform 1 0 5376 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_128
timestamp 1698175906
transform 1 0 7840 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_136
timestamp 1698175906
transform 1 0 8288 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_142
timestamp 1698175906
transform 1 0 8624 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_146
timestamp 1698175906
transform 1 0 8848 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_156
timestamp 1698175906
transform 1 0 9408 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_160
timestamp 1698175906
transform 1 0 9632 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_173
timestamp 1698175906
transform 1 0 10360 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_184
timestamp 1698175906
transform 1 0 10976 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_198
timestamp 1698175906
transform 1 0 11760 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_206
timestamp 1698175906
transform 1 0 12208 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_212
timestamp 1698175906
transform 1 0 12544 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_220
timestamp 1698175906
transform 1 0 12992 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_224
timestamp 1698175906
transform 1 0 13216 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_254
timestamp 1698175906
transform 1 0 14896 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_258
timestamp 1698175906
transform 1 0 15120 0 -1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_274
timestamp 1698175906
transform 1 0 16016 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_278
timestamp 1698175906
transform 1 0 16240 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_282
timestamp 1698175906
transform 1 0 16464 0 -1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_346
timestamp 1698175906
transform 1 0 20048 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_348
timestamp 1698175906
transform 1 0 20160 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_28
timestamp 1698175906
transform 1 0 2240 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_32
timestamp 1698175906
transform 1 0 2464 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698175906
transform 1 0 2576 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_37
timestamp 1698175906
transform 1 0 2744 0 1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_101
timestamp 1698175906
transform 1 0 6328 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_107
timestamp 1698175906
transform 1 0 6664 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_109
timestamp 1698175906
transform 1 0 6776 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_116
timestamp 1698175906
transform 1 0 7168 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_120
timestamp 1698175906
transform 1 0 7392 0 1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_136
timestamp 1698175906
transform 1 0 8288 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_140
timestamp 1698175906
transform 1 0 8512 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_150
timestamp 1698175906
transform 1 0 9072 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_168
timestamp 1698175906
transform 1 0 10080 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_172
timestamp 1698175906
transform 1 0 10304 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_174
timestamp 1698175906
transform 1 0 10416 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_183
timestamp 1698175906
transform 1 0 10920 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_199
timestamp 1698175906
transform 1 0 11816 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_207
timestamp 1698175906
transform 1 0 12264 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_209
timestamp 1698175906
transform 1 0 12376 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_216
timestamp 1698175906
transform 1 0 12768 0 1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_232
timestamp 1698175906
transform 1 0 13664 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_241
timestamp 1698175906
transform 1 0 14168 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_247
timestamp 1698175906
transform 1 0 14504 0 1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_311
timestamp 1698175906
transform 1 0 18088 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_317
timestamp 1698175906
transform 1 0 18424 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_321
timestamp 1698175906
transform 1 0 18648 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_28
timestamp 1698175906
transform 1 0 2240 0 -1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_60
timestamp 1698175906
transform 1 0 4032 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_68
timestamp 1698175906
transform 1 0 4480 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_72
timestamp 1698175906
transform 1 0 4704 0 -1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_104
timestamp 1698175906
transform 1 0 6496 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_112
timestamp 1698175906
transform 1 0 6944 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_114
timestamp 1698175906
transform 1 0 7056 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_125
timestamp 1698175906
transform 1 0 7672 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_133
timestamp 1698175906
transform 1 0 8120 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_137
timestamp 1698175906
transform 1 0 8344 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_139
timestamp 1698175906
transform 1 0 8456 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_142
timestamp 1698175906
transform 1 0 8624 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_150
timestamp 1698175906
transform 1 0 9072 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_154
timestamp 1698175906
transform 1 0 9296 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_185
timestamp 1698175906
transform 1 0 11032 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_189
timestamp 1698175906
transform 1 0 11256 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_197
timestamp 1698175906
transform 1 0 11704 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_201
timestamp 1698175906
transform 1 0 11928 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_209
timestamp 1698175906
transform 1 0 12376 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_212
timestamp 1698175906
transform 1 0 12544 0 -1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_228
timestamp 1698175906
transform 1 0 13440 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_258
timestamp 1698175906
transform 1 0 15120 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_262
timestamp 1698175906
transform 1 0 15344 0 -1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_278
timestamp 1698175906
transform 1 0 16240 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_282
timestamp 1698175906
transform 1 0 16464 0 -1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_346
timestamp 1698175906
transform 1 0 20048 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_348
timestamp 1698175906
transform 1 0 20160 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_28
timestamp 1698175906
transform 1 0 2240 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_32
timestamp 1698175906
transform 1 0 2464 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698175906
transform 1 0 2576 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_37
timestamp 1698175906
transform 1 0 2744 0 1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_101
timestamp 1698175906
transform 1 0 6328 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_142
timestamp 1698175906
transform 1 0 8624 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_146
timestamp 1698175906
transform 1 0 8848 0 1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_162
timestamp 1698175906
transform 1 0 9744 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_170
timestamp 1698175906
transform 1 0 10192 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_174
timestamp 1698175906
transform 1 0 10416 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_177
timestamp 1698175906
transform 1 0 10584 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_185
timestamp 1698175906
transform 1 0 11032 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_189
timestamp 1698175906
transform 1 0 11256 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_195
timestamp 1698175906
transform 1 0 11592 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_203
timestamp 1698175906
transform 1 0 12040 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_205
timestamp 1698175906
transform 1 0 12152 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_215
timestamp 1698175906
transform 1 0 12712 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_225
timestamp 1698175906
transform 1 0 13272 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_238
timestamp 1698175906
transform 1 0 14000 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_242
timestamp 1698175906
transform 1 0 14224 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_244
timestamp 1698175906
transform 1 0 14336 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_247
timestamp 1698175906
transform 1 0 14504 0 1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_311
timestamp 1698175906
transform 1 0 18088 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_317
timestamp 1698175906
transform 1 0 18424 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_321
timestamp 1698175906
transform 1 0 18648 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_2
timestamp 1698175906
transform 1 0 784 0 -1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_66
timestamp 1698175906
transform 1 0 4368 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_72
timestamp 1698175906
transform 1 0 4704 0 -1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_104
timestamp 1698175906
transform 1 0 6496 0 -1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_120
timestamp 1698175906
transform 1 0 7392 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_128
timestamp 1698175906
transform 1 0 7840 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_136
timestamp 1698175906
transform 1 0 8288 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_142
timestamp 1698175906
transform 1 0 8624 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_144
timestamp 1698175906
transform 1 0 8736 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_153
timestamp 1698175906
transform 1 0 9240 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_176
timestamp 1698175906
transform 1 0 10528 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_178
timestamp 1698175906
transform 1 0 10640 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_208
timestamp 1698175906
transform 1 0 12320 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_212
timestamp 1698175906
transform 1 0 12544 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_214
timestamp 1698175906
transform 1 0 12656 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_244
timestamp 1698175906
transform 1 0 14336 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_248
timestamp 1698175906
transform 1 0 14560 0 -1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_282
timestamp 1698175906
transform 1 0 16464 0 -1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_346
timestamp 1698175906
transform 1 0 20048 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_348
timestamp 1698175906
transform 1 0 20160 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_2
timestamp 1698175906
transform 1 0 784 0 1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698175906
transform 1 0 2576 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_37
timestamp 1698175906
transform 1 0 2744 0 1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_101
timestamp 1698175906
transform 1 0 6328 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_107
timestamp 1698175906
transform 1 0 6664 0 1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_115
timestamp 1698175906
transform 1 0 7112 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_125
timestamp 1698175906
transform 1 0 7672 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_169
timestamp 1698175906
transform 1 0 10136 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_173
timestamp 1698175906
transform 1 0 10360 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_177
timestamp 1698175906
transform 1 0 10584 0 1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_185
timestamp 1698175906
transform 1 0 11032 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_187
timestamp 1698175906
transform 1 0 11144 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_224
timestamp 1698175906
transform 1 0 13216 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_228
timestamp 1698175906
transform 1 0 13440 0 1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_244
timestamp 1698175906
transform 1 0 14336 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_247
timestamp 1698175906
transform 1 0 14504 0 1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_311
timestamp 1698175906
transform 1 0 18088 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_317
timestamp 1698175906
transform 1 0 18424 0 1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_2
timestamp 1698175906
transform 1 0 784 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_66
timestamp 1698175906
transform 1 0 4368 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_72
timestamp 1698175906
transform 1 0 4704 0 -1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_104
timestamp 1698175906
transform 1 0 6496 0 -1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_142
timestamp 1698175906
transform 1 0 8624 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_146
timestamp 1698175906
transform 1 0 8848 0 -1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_176
timestamp 1698175906
transform 1 0 10528 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_180
timestamp 1698175906
transform 1 0 10752 0 -1 14112
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_196
timestamp 1698175906
transform 1 0 11648 0 -1 14112
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_204
timestamp 1698175906
transform 1 0 12096 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_208
timestamp 1698175906
transform 1 0 12320 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_217
timestamp 1698175906
transform 1 0 12824 0 -1 14112
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_225
timestamp 1698175906
transform 1 0 13272 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_229
timestamp 1698175906
transform 1 0 13496 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_235
timestamp 1698175906
transform 1 0 13832 0 -1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_267
timestamp 1698175906
transform 1 0 15624 0 -1 14112
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_275
timestamp 1698175906
transform 1 0 16072 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_279
timestamp 1698175906
transform 1 0 16296 0 -1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_282
timestamp 1698175906
transform 1 0 16464 0 -1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_314
timestamp 1698175906
transform 1 0 18256 0 -1 14112
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_322
timestamp 1698175906
transform 1 0 18704 0 -1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_2
timestamp 1698175906
transform 1 0 784 0 1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698175906
transform 1 0 2576 0 1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_37
timestamp 1698175906
transform 1 0 2744 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_101
timestamp 1698175906
transform 1 0 6328 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_107
timestamp 1698175906
transform 1 0 6664 0 1 14112
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_123
timestamp 1698175906
transform 1 0 7560 0 1 14112
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_131
timestamp 1698175906
transform 1 0 8008 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_133
timestamp 1698175906
transform 1 0 8120 0 1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_136
timestamp 1698175906
transform 1 0 8288 0 1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_168
timestamp 1698175906
transform 1 0 10080 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_172
timestamp 1698175906
transform 1 0 10304 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_174
timestamp 1698175906
transform 1 0 10416 0 1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_177
timestamp 1698175906
transform 1 0 10584 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_241
timestamp 1698175906
transform 1 0 14168 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_247
timestamp 1698175906
transform 1 0 14504 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_311
timestamp 1698175906
transform 1 0 18088 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_317
timestamp 1698175906
transform 1 0 18424 0 1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_2
timestamp 1698175906
transform 1 0 784 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_66
timestamp 1698175906
transform 1 0 4368 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_72
timestamp 1698175906
transform 1 0 4704 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_136
timestamp 1698175906
transform 1 0 8288 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_142
timestamp 1698175906
transform 1 0 8624 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_206
timestamp 1698175906
transform 1 0 12208 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_212
timestamp 1698175906
transform 1 0 12544 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_276
timestamp 1698175906
transform 1 0 16128 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_282
timestamp 1698175906
transform 1 0 16464 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_346
timestamp 1698175906
transform 1 0 20048 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_348
timestamp 1698175906
transform 1 0 20160 0 -1 14896
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698175906
transform 1 0 784 0 1 14896
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698175906
transform 1 0 2576 0 1 14896
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_37
timestamp 1698175906
transform 1 0 2744 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_101
timestamp 1698175906
transform 1 0 6328 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_107
timestamp 1698175906
transform 1 0 6664 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_171
timestamp 1698175906
transform 1 0 10248 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_177
timestamp 1698175906
transform 1 0 10584 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_241
timestamp 1698175906
transform 1 0 14168 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_247
timestamp 1698175906
transform 1 0 14504 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_311
timestamp 1698175906
transform 1 0 18088 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_317
timestamp 1698175906
transform 1 0 18424 0 1 14896
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2
timestamp 1698175906
transform 1 0 784 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_66
timestamp 1698175906
transform 1 0 4368 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_72
timestamp 1698175906
transform 1 0 4704 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_136
timestamp 1698175906
transform 1 0 8288 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_142
timestamp 1698175906
transform 1 0 8624 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_206
timestamp 1698175906
transform 1 0 12208 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_212
timestamp 1698175906
transform 1 0 12544 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_276
timestamp 1698175906
transform 1 0 16128 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_282
timestamp 1698175906
transform 1 0 16464 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_346
timestamp 1698175906
transform 1 0 20048 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_348
timestamp 1698175906
transform 1 0 20160 0 -1 15680
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_2
timestamp 1698175906
transform 1 0 784 0 1 15680
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698175906
transform 1 0 2576 0 1 15680
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_37
timestamp 1698175906
transform 1 0 2744 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_101
timestamp 1698175906
transform 1 0 6328 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_107
timestamp 1698175906
transform 1 0 6664 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_171
timestamp 1698175906
transform 1 0 10248 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_177
timestamp 1698175906
transform 1 0 10584 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_241
timestamp 1698175906
transform 1 0 14168 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_247
timestamp 1698175906
transform 1 0 14504 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_311
timestamp 1698175906
transform 1 0 18088 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_317
timestamp 1698175906
transform 1 0 18424 0 1 15680
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2
timestamp 1698175906
transform 1 0 784 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_66
timestamp 1698175906
transform 1 0 4368 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_72
timestamp 1698175906
transform 1 0 4704 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_136
timestamp 1698175906
transform 1 0 8288 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_142
timestamp 1698175906
transform 1 0 8624 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_206
timestamp 1698175906
transform 1 0 12208 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_212
timestamp 1698175906
transform 1 0 12544 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_276
timestamp 1698175906
transform 1 0 16128 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_282
timestamp 1698175906
transform 1 0 16464 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_346
timestamp 1698175906
transform 1 0 20048 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_348
timestamp 1698175906
transform 1 0 20160 0 -1 16464
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698175906
transform 1 0 784 0 1 16464
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698175906
transform 1 0 2576 0 1 16464
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_37
timestamp 1698175906
transform 1 0 2744 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_101
timestamp 1698175906
transform 1 0 6328 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_107
timestamp 1698175906
transform 1 0 6664 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_171
timestamp 1698175906
transform 1 0 10248 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_177
timestamp 1698175906
transform 1 0 10584 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_241
timestamp 1698175906
transform 1 0 14168 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_247
timestamp 1698175906
transform 1 0 14504 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_311
timestamp 1698175906
transform 1 0 18088 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_317
timestamp 1698175906
transform 1 0 18424 0 1 16464
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_2
timestamp 1698175906
transform 1 0 784 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_66
timestamp 1698175906
transform 1 0 4368 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_72
timestamp 1698175906
transform 1 0 4704 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_136
timestamp 1698175906
transform 1 0 8288 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_142
timestamp 1698175906
transform 1 0 8624 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_206
timestamp 1698175906
transform 1 0 12208 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_212
timestamp 1698175906
transform 1 0 12544 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_276
timestamp 1698175906
transform 1 0 16128 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_282
timestamp 1698175906
transform 1 0 16464 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_346
timestamp 1698175906
transform 1 0 20048 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_348
timestamp 1698175906
transform 1 0 20160 0 -1 17248
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698175906
transform 1 0 784 0 1 17248
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698175906
transform 1 0 2576 0 1 17248
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_37
timestamp 1698175906
transform 1 0 2744 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_101
timestamp 1698175906
transform 1 0 6328 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_107
timestamp 1698175906
transform 1 0 6664 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_171
timestamp 1698175906
transform 1 0 10248 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_177
timestamp 1698175906
transform 1 0 10584 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_241
timestamp 1698175906
transform 1 0 14168 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_247
timestamp 1698175906
transform 1 0 14504 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_311
timestamp 1698175906
transform 1 0 18088 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_317
timestamp 1698175906
transform 1 0 18424 0 1 17248
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2
timestamp 1698175906
transform 1 0 784 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1698175906
transform 1 0 4368 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_72
timestamp 1698175906
transform 1 0 4704 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_136
timestamp 1698175906
transform 1 0 8288 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_142
timestamp 1698175906
transform 1 0 8624 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_206
timestamp 1698175906
transform 1 0 12208 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_212
timestamp 1698175906
transform 1 0 12544 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_276
timestamp 1698175906
transform 1 0 16128 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_282
timestamp 1698175906
transform 1 0 16464 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_346
timestamp 1698175906
transform 1 0 20048 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_348
timestamp 1698175906
transform 1 0 20160 0 -1 18032
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_2
timestamp 1698175906
transform 1 0 784 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698175906
transform 1 0 2576 0 1 18032
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_37
timestamp 1698175906
transform 1 0 2744 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_101
timestamp 1698175906
transform 1 0 6328 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_107
timestamp 1698175906
transform 1 0 6664 0 1 18032
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_123
timestamp 1698175906
transform 1 0 7560 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_153
timestamp 1698175906
transform 1 0 9240 0 1 18032
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_169
timestamp 1698175906
transform 1 0 10136 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_173
timestamp 1698175906
transform 1 0 10360 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_177
timestamp 1698175906
transform 1 0 10584 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_241
timestamp 1698175906
transform 1 0 14168 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_247
timestamp 1698175906
transform 1 0 14504 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_311
timestamp 1698175906
transform 1 0 18088 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_317
timestamp 1698175906
transform 1 0 18424 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_2
timestamp 1698175906
transform 1 0 784 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_66
timestamp 1698175906
transform 1 0 4368 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_72
timestamp 1698175906
transform 1 0 4704 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_136
timestamp 1698175906
transform 1 0 8288 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_142
timestamp 1698175906
transform 1 0 8624 0 -1 18816
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_150
timestamp 1698175906
transform 1 0 9072 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_154
timestamp 1698175906
transform 1 0 9296 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_156
timestamp 1698175906
transform 1 0 9408 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_183
timestamp 1698175906
transform 1 0 10920 0 -1 18816
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_199
timestamp 1698175906
transform 1 0 11816 0 -1 18816
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_207
timestamp 1698175906
transform 1 0 12264 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_209
timestamp 1698175906
transform 1 0 12376 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_212
timestamp 1698175906
transform 1 0 12544 0 -1 18816
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_220
timestamp 1698175906
transform 1 0 12992 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_222
timestamp 1698175906
transform 1 0 13104 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_249
timestamp 1698175906
transform 1 0 14616 0 -1 18816
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_265
timestamp 1698175906
transform 1 0 15512 0 -1 18816
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_273
timestamp 1698175906
transform 1 0 15960 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_277
timestamp 1698175906
transform 1 0 16184 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_279
timestamp 1698175906
transform 1 0 16296 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_282
timestamp 1698175906
transform 1 0 16464 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_346
timestamp 1698175906
transform 1 0 20048 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_348
timestamp 1698175906
transform 1 0 20160 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_2
timestamp 1698175906
transform 1 0 784 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_36
timestamp 1698175906
transform 1 0 2688 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_70
timestamp 1698175906
transform 1 0 4592 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_104
timestamp 1698175906
transform 1 0 6496 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_164
timestamp 1698175906
transform 1 0 9856 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_168
timestamp 1698175906
transform 1 0 10080 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_172
timestamp 1698175906
transform 1 0 10304 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_174
timestamp 1698175906
transform 1 0 10416 0 1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_201
timestamp 1698175906
transform 1 0 11928 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_203
timestamp 1698175906
transform 1 0 12040 0 1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_232
timestamp 1698175906
transform 1 0 13664 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_236
timestamp 1698175906
transform 1 0 13888 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_240
timestamp 1698175906
transform 1 0 14112 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_274
timestamp 1698175906
transform 1 0 16016 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_308
timestamp 1698175906
transform 1 0 17920 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_342
timestamp 1698175906
transform 1 0 19824 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_346
timestamp 1698175906
transform 1 0 20048 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_348
timestamp 1698175906
transform 1 0 20160 0 1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 7784 0 1 18032
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output2
timestamp 1698175906
transform -1 0 2240 0 1 12544
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output3
timestamp 1698175906
transform 1 0 12544 0 -1 2352
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output4
timestamp 1698175906
transform 1 0 18760 0 1 11760
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output5
timestamp 1698175906
transform 1 0 10472 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output6
timestamp 1698175906
transform -1 0 2240 0 -1 10976
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output7
timestamp 1698175906
transform 1 0 18760 0 -1 8624
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output8
timestamp 1698175906
transform 1 0 18760 0 -1 14112
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output9
timestamp 1698175906
transform -1 0 2240 0 -1 10192
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output10
timestamp 1698175906
transform 1 0 18760 0 1 8624
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output11
timestamp 1698175906
transform 1 0 18760 0 1 10192
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output12
timestamp 1698175906
transform -1 0 2240 0 -1 11760
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output13
timestamp 1698175906
transform -1 0 2240 0 -1 12544
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output14
timestamp 1698175906
transform -1 0 2240 0 1 11760
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output15
timestamp 1698175906
transform 1 0 8456 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output16
timestamp 1698175906
transform 1 0 10640 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output17
timestamp 1698175906
transform 1 0 8400 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output18
timestamp 1698175906
transform 1 0 18760 0 1 12544
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output19
timestamp 1698175906
transform 1 0 13160 0 -1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output20
timestamp 1698175906
transform 1 0 18760 0 1 10976
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output21
timestamp 1698175906
transform 1 0 12208 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output22
timestamp 1698175906
transform -1 0 2240 0 1 8624
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output23
timestamp 1698175906
transform 1 0 9464 0 -1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output24
timestamp 1698175906
transform 1 0 18760 0 -1 7840
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output25
timestamp 1698175906
transform 1 0 12208 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output26
timestamp 1698175906
transform 1 0 12824 0 1 2352
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_45 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 672 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698175906
transform -1 0 20328 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_46
timestamp 1698175906
transform 1 0 672 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698175906
transform -1 0 20328 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_47
timestamp 1698175906
transform 1 0 672 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698175906
transform -1 0 20328 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_48
timestamp 1698175906
transform 1 0 672 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698175906
transform -1 0 20328 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_49
timestamp 1698175906
transform 1 0 672 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698175906
transform -1 0 20328 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_50
timestamp 1698175906
transform 1 0 672 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698175906
transform -1 0 20328 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_51
timestamp 1698175906
transform 1 0 672 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698175906
transform -1 0 20328 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_52
timestamp 1698175906
transform 1 0 672 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698175906
transform -1 0 20328 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_53
timestamp 1698175906
transform 1 0 672 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698175906
transform -1 0 20328 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_54
timestamp 1698175906
transform 1 0 672 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698175906
transform -1 0 20328 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_55
timestamp 1698175906
transform 1 0 672 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698175906
transform -1 0 20328 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_56
timestamp 1698175906
transform 1 0 672 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698175906
transform -1 0 20328 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_57
timestamp 1698175906
transform 1 0 672 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698175906
transform -1 0 20328 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_58
timestamp 1698175906
transform 1 0 672 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698175906
transform -1 0 20328 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_59
timestamp 1698175906
transform 1 0 672 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698175906
transform -1 0 20328 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_60
timestamp 1698175906
transform 1 0 672 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698175906
transform -1 0 20328 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_61
timestamp 1698175906
transform 1 0 672 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698175906
transform -1 0 20328 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_62
timestamp 1698175906
transform 1 0 672 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698175906
transform -1 0 20328 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_63
timestamp 1698175906
transform 1 0 672 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698175906
transform -1 0 20328 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_64
timestamp 1698175906
transform 1 0 672 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698175906
transform -1 0 20328 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_65
timestamp 1698175906
transform 1 0 672 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698175906
transform -1 0 20328 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_66
timestamp 1698175906
transform 1 0 672 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698175906
transform -1 0 20328 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_67
timestamp 1698175906
transform 1 0 672 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698175906
transform -1 0 20328 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_68
timestamp 1698175906
transform 1 0 672 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698175906
transform -1 0 20328 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_69
timestamp 1698175906
transform 1 0 672 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698175906
transform -1 0 20328 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_70
timestamp 1698175906
transform 1 0 672 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698175906
transform -1 0 20328 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_71
timestamp 1698175906
transform 1 0 672 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698175906
transform -1 0 20328 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_72
timestamp 1698175906
transform 1 0 672 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698175906
transform -1 0 20328 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_73
timestamp 1698175906
transform 1 0 672 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698175906
transform -1 0 20328 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_74
timestamp 1698175906
transform 1 0 672 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698175906
transform -1 0 20328 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_75
timestamp 1698175906
transform 1 0 672 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698175906
transform -1 0 20328 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_76
timestamp 1698175906
transform 1 0 672 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698175906
transform -1 0 20328 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_77
timestamp 1698175906
transform 1 0 672 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698175906
transform -1 0 20328 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_78
timestamp 1698175906
transform 1 0 672 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698175906
transform -1 0 20328 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_79
timestamp 1698175906
transform 1 0 672 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698175906
transform -1 0 20328 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_80
timestamp 1698175906
transform 1 0 672 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698175906
transform -1 0 20328 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_81
timestamp 1698175906
transform 1 0 672 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698175906
transform -1 0 20328 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_82
timestamp 1698175906
transform 1 0 672 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698175906
transform -1 0 20328 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_83
timestamp 1698175906
transform 1 0 672 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698175906
transform -1 0 20328 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_84
timestamp 1698175906
transform 1 0 672 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698175906
transform -1 0 20328 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_85
timestamp 1698175906
transform 1 0 672 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698175906
transform -1 0 20328 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_86
timestamp 1698175906
transform 1 0 672 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698175906
transform -1 0 20328 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_87
timestamp 1698175906
transform 1 0 672 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698175906
transform -1 0 20328 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_88
timestamp 1698175906
transform 1 0 672 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698175906
transform -1 0 20328 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_89
timestamp 1698175906
transform 1 0 672 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698175906
transform -1 0 20328 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_90 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 2576 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_91
timestamp 1698175906
transform 1 0 4480 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_92
timestamp 1698175906
transform 1 0 6384 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_93
timestamp 1698175906
transform 1 0 8288 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_94
timestamp 1698175906
transform 1 0 10192 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_95
timestamp 1698175906
transform 1 0 12096 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_96
timestamp 1698175906
transform 1 0 14000 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_97
timestamp 1698175906
transform 1 0 15904 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_98
timestamp 1698175906
transform 1 0 17808 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_99
timestamp 1698175906
transform 1 0 19712 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_100
timestamp 1698175906
transform 1 0 4592 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_101
timestamp 1698175906
transform 1 0 8512 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_102
timestamp 1698175906
transform 1 0 12432 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_103
timestamp 1698175906
transform 1 0 16352 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_104
timestamp 1698175906
transform 1 0 2632 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_105
timestamp 1698175906
transform 1 0 6552 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_106
timestamp 1698175906
transform 1 0 10472 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_107
timestamp 1698175906
transform 1 0 14392 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_108
timestamp 1698175906
transform 1 0 18312 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_109
timestamp 1698175906
transform 1 0 4592 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_110
timestamp 1698175906
transform 1 0 8512 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_111
timestamp 1698175906
transform 1 0 12432 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_112
timestamp 1698175906
transform 1 0 16352 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_113
timestamp 1698175906
transform 1 0 2632 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_114
timestamp 1698175906
transform 1 0 6552 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_115
timestamp 1698175906
transform 1 0 10472 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_116
timestamp 1698175906
transform 1 0 14392 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_117
timestamp 1698175906
transform 1 0 18312 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_118
timestamp 1698175906
transform 1 0 4592 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_119
timestamp 1698175906
transform 1 0 8512 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_120
timestamp 1698175906
transform 1 0 12432 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_121
timestamp 1698175906
transform 1 0 16352 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_122
timestamp 1698175906
transform 1 0 2632 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_123
timestamp 1698175906
transform 1 0 6552 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_124
timestamp 1698175906
transform 1 0 10472 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_125
timestamp 1698175906
transform 1 0 14392 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_126
timestamp 1698175906
transform 1 0 18312 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_127
timestamp 1698175906
transform 1 0 4592 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_128
timestamp 1698175906
transform 1 0 8512 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_129
timestamp 1698175906
transform 1 0 12432 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_130
timestamp 1698175906
transform 1 0 16352 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_131
timestamp 1698175906
transform 1 0 2632 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_132
timestamp 1698175906
transform 1 0 6552 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_133
timestamp 1698175906
transform 1 0 10472 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_134
timestamp 1698175906
transform 1 0 14392 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_135
timestamp 1698175906
transform 1 0 18312 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_136
timestamp 1698175906
transform 1 0 4592 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_137
timestamp 1698175906
transform 1 0 8512 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_138
timestamp 1698175906
transform 1 0 12432 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_139
timestamp 1698175906
transform 1 0 16352 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_140
timestamp 1698175906
transform 1 0 2632 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_141
timestamp 1698175906
transform 1 0 6552 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_142
timestamp 1698175906
transform 1 0 10472 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_143
timestamp 1698175906
transform 1 0 14392 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_144
timestamp 1698175906
transform 1 0 18312 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_145
timestamp 1698175906
transform 1 0 4592 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_146
timestamp 1698175906
transform 1 0 8512 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_147
timestamp 1698175906
transform 1 0 12432 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_148
timestamp 1698175906
transform 1 0 16352 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_149
timestamp 1698175906
transform 1 0 2632 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_150
timestamp 1698175906
transform 1 0 6552 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_151
timestamp 1698175906
transform 1 0 10472 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_152
timestamp 1698175906
transform 1 0 14392 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_153
timestamp 1698175906
transform 1 0 18312 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_154
timestamp 1698175906
transform 1 0 4592 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_155
timestamp 1698175906
transform 1 0 8512 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_156
timestamp 1698175906
transform 1 0 12432 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_157
timestamp 1698175906
transform 1 0 16352 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_158
timestamp 1698175906
transform 1 0 2632 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_159
timestamp 1698175906
transform 1 0 6552 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_160
timestamp 1698175906
transform 1 0 10472 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_161
timestamp 1698175906
transform 1 0 14392 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_162
timestamp 1698175906
transform 1 0 18312 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_163
timestamp 1698175906
transform 1 0 4592 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_164
timestamp 1698175906
transform 1 0 8512 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_165
timestamp 1698175906
transform 1 0 12432 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_166
timestamp 1698175906
transform 1 0 16352 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_167
timestamp 1698175906
transform 1 0 2632 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_168
timestamp 1698175906
transform 1 0 6552 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_169
timestamp 1698175906
transform 1 0 10472 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_170
timestamp 1698175906
transform 1 0 14392 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_171
timestamp 1698175906
transform 1 0 18312 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_172
timestamp 1698175906
transform 1 0 4592 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_173
timestamp 1698175906
transform 1 0 8512 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_174
timestamp 1698175906
transform 1 0 12432 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_175
timestamp 1698175906
transform 1 0 16352 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_176
timestamp 1698175906
transform 1 0 2632 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_177
timestamp 1698175906
transform 1 0 6552 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_178
timestamp 1698175906
transform 1 0 10472 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_179
timestamp 1698175906
transform 1 0 14392 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_180
timestamp 1698175906
transform 1 0 18312 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_181
timestamp 1698175906
transform 1 0 4592 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_182
timestamp 1698175906
transform 1 0 8512 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_183
timestamp 1698175906
transform 1 0 12432 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_184
timestamp 1698175906
transform 1 0 16352 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_185
timestamp 1698175906
transform 1 0 2632 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_186
timestamp 1698175906
transform 1 0 6552 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_187
timestamp 1698175906
transform 1 0 10472 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_188
timestamp 1698175906
transform 1 0 14392 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_189
timestamp 1698175906
transform 1 0 18312 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_190
timestamp 1698175906
transform 1 0 4592 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_191
timestamp 1698175906
transform 1 0 8512 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_192
timestamp 1698175906
transform 1 0 12432 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_193
timestamp 1698175906
transform 1 0 16352 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_194
timestamp 1698175906
transform 1 0 2632 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_195
timestamp 1698175906
transform 1 0 6552 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_196
timestamp 1698175906
transform 1 0 10472 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_197
timestamp 1698175906
transform 1 0 14392 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_198
timestamp 1698175906
transform 1 0 18312 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_199
timestamp 1698175906
transform 1 0 4592 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_200
timestamp 1698175906
transform 1 0 8512 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_201
timestamp 1698175906
transform 1 0 12432 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_202
timestamp 1698175906
transform 1 0 16352 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_203
timestamp 1698175906
transform 1 0 2632 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_204
timestamp 1698175906
transform 1 0 6552 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_205
timestamp 1698175906
transform 1 0 10472 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_206
timestamp 1698175906
transform 1 0 14392 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_207
timestamp 1698175906
transform 1 0 18312 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_208
timestamp 1698175906
transform 1 0 4592 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_209
timestamp 1698175906
transform 1 0 8512 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_210
timestamp 1698175906
transform 1 0 12432 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_211
timestamp 1698175906
transform 1 0 16352 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_212
timestamp 1698175906
transform 1 0 2632 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_213
timestamp 1698175906
transform 1 0 6552 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_214
timestamp 1698175906
transform 1 0 10472 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_215
timestamp 1698175906
transform 1 0 14392 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_216
timestamp 1698175906
transform 1 0 18312 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_217
timestamp 1698175906
transform 1 0 4592 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_218
timestamp 1698175906
transform 1 0 8512 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_219
timestamp 1698175906
transform 1 0 12432 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_220
timestamp 1698175906
transform 1 0 16352 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_221
timestamp 1698175906
transform 1 0 2632 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_222
timestamp 1698175906
transform 1 0 6552 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_223
timestamp 1698175906
transform 1 0 10472 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_224
timestamp 1698175906
transform 1 0 14392 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_225
timestamp 1698175906
transform 1 0 18312 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_226
timestamp 1698175906
transform 1 0 4592 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_227
timestamp 1698175906
transform 1 0 8512 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_228
timestamp 1698175906
transform 1 0 12432 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_229
timestamp 1698175906
transform 1 0 16352 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_230
timestamp 1698175906
transform 1 0 2632 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_231
timestamp 1698175906
transform 1 0 6552 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_232
timestamp 1698175906
transform 1 0 10472 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_233
timestamp 1698175906
transform 1 0 14392 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_234
timestamp 1698175906
transform 1 0 18312 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_235
timestamp 1698175906
transform 1 0 4592 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_236
timestamp 1698175906
transform 1 0 8512 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_237
timestamp 1698175906
transform 1 0 12432 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_238
timestamp 1698175906
transform 1 0 16352 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_239
timestamp 1698175906
transform 1 0 2632 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_240
timestamp 1698175906
transform 1 0 6552 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_241
timestamp 1698175906
transform 1 0 10472 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_242
timestamp 1698175906
transform 1 0 14392 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_243
timestamp 1698175906
transform 1 0 18312 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_244
timestamp 1698175906
transform 1 0 4592 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_245
timestamp 1698175906
transform 1 0 8512 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_246
timestamp 1698175906
transform 1 0 12432 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_247
timestamp 1698175906
transform 1 0 16352 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_248
timestamp 1698175906
transform 1 0 2632 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_249
timestamp 1698175906
transform 1 0 6552 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_250
timestamp 1698175906
transform 1 0 10472 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_251
timestamp 1698175906
transform 1 0 14392 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_252
timestamp 1698175906
transform 1 0 18312 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_253
timestamp 1698175906
transform 1 0 4592 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_254
timestamp 1698175906
transform 1 0 8512 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_255
timestamp 1698175906
transform 1 0 12432 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_256
timestamp 1698175906
transform 1 0 16352 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_257
timestamp 1698175906
transform 1 0 2632 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_258
timestamp 1698175906
transform 1 0 6552 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_259
timestamp 1698175906
transform 1 0 10472 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_260
timestamp 1698175906
transform 1 0 14392 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_261
timestamp 1698175906
transform 1 0 18312 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_262
timestamp 1698175906
transform 1 0 4592 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_263
timestamp 1698175906
transform 1 0 8512 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_264
timestamp 1698175906
transform 1 0 12432 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_265
timestamp 1698175906
transform 1 0 16352 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_266
timestamp 1698175906
transform 1 0 2632 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_267
timestamp 1698175906
transform 1 0 6552 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_268
timestamp 1698175906
transform 1 0 10472 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_269
timestamp 1698175906
transform 1 0 14392 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_270
timestamp 1698175906
transform 1 0 18312 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_271
timestamp 1698175906
transform 1 0 4592 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_272
timestamp 1698175906
transform 1 0 8512 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_273
timestamp 1698175906
transform 1 0 12432 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_274
timestamp 1698175906
transform 1 0 16352 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_275
timestamp 1698175906
transform 1 0 2632 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_276
timestamp 1698175906
transform 1 0 6552 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_277
timestamp 1698175906
transform 1 0 10472 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_278
timestamp 1698175906
transform 1 0 14392 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_279
timestamp 1698175906
transform 1 0 18312 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_280
timestamp 1698175906
transform 1 0 4592 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_281
timestamp 1698175906
transform 1 0 8512 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_282
timestamp 1698175906
transform 1 0 12432 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_283
timestamp 1698175906
transform 1 0 16352 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_284
timestamp 1698175906
transform 1 0 2632 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_285
timestamp 1698175906
transform 1 0 6552 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_286
timestamp 1698175906
transform 1 0 10472 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_287
timestamp 1698175906
transform 1 0 14392 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_288
timestamp 1698175906
transform 1 0 18312 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_289
timestamp 1698175906
transform 1 0 4592 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_290
timestamp 1698175906
transform 1 0 8512 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_291
timestamp 1698175906
transform 1 0 12432 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_292
timestamp 1698175906
transform 1 0 16352 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_293
timestamp 1698175906
transform 1 0 2576 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_294
timestamp 1698175906
transform 1 0 4480 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_295
timestamp 1698175906
transform 1 0 6384 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_296
timestamp 1698175906
transform 1 0 8288 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_297
timestamp 1698175906
transform 1 0 10192 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_298
timestamp 1698175906
transform 1 0 12096 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_299
timestamp 1698175906
transform 1 0 14000 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_300
timestamp 1698175906
transform 1 0 15904 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_301
timestamp 1698175906
transform 1 0 17808 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_302
timestamp 1698175906
transform 1 0 19712 0 1 18816
box -43 -43 155 435
<< labels >>
flabel metal3 s 0 13440 400 13496 0 FreeSans 224 0 0 0 clk
port 0 nsew signal input
flabel metal2 s 7728 20600 7784 21000 0 FreeSans 224 90 0 0 segm[0]
port 1 nsew signal tristate
flabel metal3 s 0 12432 400 12488 0 FreeSans 224 0 0 0 segm[10]
port 2 nsew signal tristate
flabel metal2 s 12432 0 12488 400 0 FreeSans 224 90 0 0 segm[11]
port 3 nsew signal tristate
flabel metal3 s 20600 11760 21000 11816 0 FreeSans 224 0 0 0 segm[12]
port 4 nsew signal tristate
flabel metal2 s 10416 20600 10472 21000 0 FreeSans 224 90 0 0 segm[13]
port 5 nsew signal tristate
flabel metal3 s 0 10416 400 10472 0 FreeSans 224 0 0 0 segm[1]
port 6 nsew signal tristate
flabel metal3 s 20600 8400 21000 8456 0 FreeSans 224 0 0 0 segm[2]
port 7 nsew signal tristate
flabel metal3 s 20600 13776 21000 13832 0 FreeSans 224 0 0 0 segm[3]
port 8 nsew signal tristate
flabel metal3 s 0 9744 400 9800 0 FreeSans 224 0 0 0 segm[4]
port 9 nsew signal tristate
flabel metal3 s 20600 8736 21000 8792 0 FreeSans 224 0 0 0 segm[5]
port 10 nsew signal tristate
flabel metal3 s 20600 10080 21000 10136 0 FreeSans 224 0 0 0 segm[6]
port 11 nsew signal tristate
flabel metal3 s 0 11424 400 11480 0 FreeSans 224 0 0 0 segm[7]
port 12 nsew signal tristate
flabel metal3 s 0 12096 400 12152 0 FreeSans 224 0 0 0 segm[8]
port 13 nsew signal tristate
flabel metal3 s 0 11760 400 11816 0 FreeSans 224 0 0 0 segm[9]
port 14 nsew signal tristate
flabel metal2 s 8400 0 8456 400 0 FreeSans 224 90 0 0 sel[0]
port 15 nsew signal tristate
flabel metal2 s 10752 0 10808 400 0 FreeSans 224 90 0 0 sel[10]
port 16 nsew signal tristate
flabel metal2 s 8064 20600 8120 21000 0 FreeSans 224 90 0 0 sel[11]
port 17 nsew signal tristate
flabel metal3 s 20600 12432 21000 12488 0 FreeSans 224 0 0 0 sel[1]
port 18 nsew signal tristate
flabel metal2 s 13104 20600 13160 21000 0 FreeSans 224 90 0 0 sel[2]
port 19 nsew signal tristate
flabel metal3 s 20600 10752 21000 10808 0 FreeSans 224 0 0 0 sel[3]
port 20 nsew signal tristate
flabel metal2 s 12096 20600 12152 21000 0 FreeSans 224 90 0 0 sel[4]
port 21 nsew signal tristate
flabel metal3 s 0 8400 400 8456 0 FreeSans 224 0 0 0 sel[5]
port 22 nsew signal tristate
flabel metal2 s 9408 20600 9464 21000 0 FreeSans 224 90 0 0 sel[6]
port 23 nsew signal tristate
flabel metal3 s 20600 7392 21000 7448 0 FreeSans 224 0 0 0 sel[7]
port 24 nsew signal tristate
flabel metal2 s 11760 0 11816 400 0 FreeSans 224 90 0 0 sel[8]
port 25 nsew signal tristate
flabel metal2 s 12768 0 12824 400 0 FreeSans 224 90 0 0 sel[9]
port 26 nsew signal tristate
flabel metal4 s 2224 1538 2384 19238 0 FreeSans 640 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 17584 1538 17744 19238 0 FreeSans 640 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 9904 1538 10064 19238 0 FreeSans 640 90 0 0 vss
port 28 nsew ground bidirectional
rlabel metal1 10500 19208 10500 19208 0 vdd
rlabel metal1 10500 18816 10500 18816 0 vss
rlabel metal2 10780 6916 10780 6916 0 _000_
rlabel metal3 14672 8484 14672 8484 0 _001_
rlabel metal2 14420 8120 14420 8120 0 _002_
rlabel metal2 7308 9212 7308 9212 0 _003_
rlabel metal2 9156 6888 9156 6888 0 _004_
rlabel metal2 9660 12152 9660 12152 0 _005_
rlabel metal2 11564 11004 11564 11004 0 _006_
rlabel metal3 8764 13244 8764 13244 0 _007_
rlabel metal2 6636 8680 6636 8680 0 _008_
rlabel metal2 11340 12908 11340 12908 0 _009_
rlabel metal3 14140 10724 14140 10724 0 _010_
rlabel metal2 12068 13692 12068 13692 0 _011_
rlabel metal2 13972 12068 13972 12068 0 _012_
rlabel metal2 7140 7812 7140 7812 0 _013_
rlabel metal2 9380 13650 9380 13650 0 _014_
rlabel metal2 6076 10136 6076 10136 0 _015_
rlabel metal2 6188 9408 6188 9408 0 _016_
rlabel metal2 13468 7028 13468 7028 0 _017_
rlabel metal2 10836 7952 10836 7952 0 _018_
rlabel metal2 7420 13748 7420 13748 0 _019_
rlabel metal2 13160 12796 13160 12796 0 _020_
rlabel metal2 14420 9408 14420 9408 0 _021_
rlabel metal2 8764 11536 8764 11536 0 _022_
rlabel metal3 7112 11508 7112 11508 0 _023_
rlabel metal2 7308 12572 7308 12572 0 _024_
rlabel metal2 11508 6832 11508 6832 0 _025_
rlabel metal2 13468 11284 13468 11284 0 _026_
rlabel metal2 12292 7336 12292 7336 0 _027_
rlabel metal2 11172 13524 11172 13524 0 _028_
rlabel metal2 13664 10164 13664 10164 0 _029_
rlabel metal2 9772 10976 9772 10976 0 _030_
rlabel metal2 9604 8372 9604 8372 0 _031_
rlabel metal2 11676 10444 11676 10444 0 _032_
rlabel metal2 10836 10584 10836 10584 0 _033_
rlabel metal3 11200 10836 11200 10836 0 _034_
rlabel metal3 9212 13132 9212 13132 0 _035_
rlabel metal2 11732 9744 11732 9744 0 _036_
rlabel metal2 8876 12544 8876 12544 0 _037_
rlabel metal2 6748 10444 6748 10444 0 _038_
rlabel metal2 6972 8624 6972 8624 0 _039_
rlabel metal2 7140 8848 7140 8848 0 _040_
rlabel metal2 6412 8820 6412 8820 0 _041_
rlabel metal2 6244 9268 6244 9268 0 _042_
rlabel metal2 6916 10276 6916 10276 0 _043_
rlabel metal2 12124 12936 12124 12936 0 _044_
rlabel metal2 11564 13076 11564 13076 0 _045_
rlabel metal2 13804 11340 13804 11340 0 _046_
rlabel metal2 14140 10556 14140 10556 0 _047_
rlabel metal2 12740 13972 12740 13972 0 _048_
rlabel metal2 12600 13916 12600 13916 0 _049_
rlabel metal2 14084 12292 14084 12292 0 _050_
rlabel metal2 7868 8316 7868 8316 0 _051_
rlabel metal2 7868 9100 7868 9100 0 _052_
rlabel metal2 7532 8232 7532 8232 0 _053_
rlabel metal2 10136 13132 10136 13132 0 _054_
rlabel metal2 9828 13328 9828 13328 0 _055_
rlabel metal2 6972 10780 6972 10780 0 _056_
rlabel metal3 6524 10276 6524 10276 0 _057_
rlabel metal2 6356 9240 6356 9240 0 _058_
rlabel metal2 7140 11172 7140 11172 0 _059_
rlabel metal2 13132 7728 13132 7728 0 _060_
rlabel metal2 10556 7980 10556 7980 0 _061_
rlabel metal2 13860 11088 13860 11088 0 _062_
rlabel metal2 7476 12264 7476 12264 0 _063_
rlabel metal2 7700 13580 7700 13580 0 _064_
rlabel metal3 13384 13804 13384 13804 0 _065_
rlabel metal2 13692 11172 13692 11172 0 _066_
rlabel metal2 13916 9492 13916 9492 0 _067_
rlabel metal2 8876 10892 8876 10892 0 _068_
rlabel metal2 8708 11200 8708 11200 0 _069_
rlabel metal3 7532 11620 7532 11620 0 _070_
rlabel metal2 7140 11368 7140 11368 0 _071_
rlabel metal2 7588 12684 7588 12684 0 _072_
rlabel metal3 10444 7140 10444 7140 0 _073_
rlabel metal2 11788 8568 11788 8568 0 _074_
rlabel metal2 11452 7336 11452 7336 0 _075_
rlabel metal2 11788 7196 11788 7196 0 _076_
rlabel metal2 13524 11200 13524 11200 0 _077_
rlabel metal2 13412 11144 13412 11144 0 _078_
rlabel metal3 12516 6804 12516 6804 0 _079_
rlabel metal2 9884 9212 9884 9212 0 _080_
rlabel metal3 7252 8736 7252 8736 0 _081_
rlabel metal3 10612 7532 10612 7532 0 _082_
rlabel metal2 10276 10052 10276 10052 0 _083_
rlabel metal2 9016 9996 9016 9996 0 _084_
rlabel metal2 12628 10612 12628 10612 0 _085_
rlabel metal2 9380 9772 9380 9772 0 _086_
rlabel metal2 13580 9240 13580 9240 0 _087_
rlabel metal2 11004 7700 11004 7700 0 _088_
rlabel metal3 12684 10052 12684 10052 0 _089_
rlabel metal2 7476 11340 7476 11340 0 _090_
rlabel metal2 12180 6944 12180 6944 0 _091_
rlabel metal2 10864 11844 10864 11844 0 _092_
rlabel metal3 11984 7532 11984 7532 0 _093_
rlabel metal2 11452 7532 11452 7532 0 _094_
rlabel metal2 9576 9212 9576 9212 0 _095_
rlabel metal2 10780 8848 10780 8848 0 _096_
rlabel metal2 10640 9716 10640 9716 0 _097_
rlabel metal2 9016 7308 9016 7308 0 _098_
rlabel metal2 14140 10220 14140 10220 0 _099_
rlabel metal2 14252 8988 14252 8988 0 _100_
rlabel metal3 9576 9940 9576 9940 0 _101_
rlabel metal2 13244 10836 13244 10836 0 _102_
rlabel metal2 13524 8008 13524 8008 0 _103_
rlabel metal2 8792 8428 8792 8428 0 _104_
rlabel metal2 8260 8960 8260 8960 0 _105_
rlabel metal2 8428 8792 8428 8792 0 _106_
rlabel metal3 14308 8820 14308 8820 0 _107_
rlabel metal2 14980 8848 14980 8848 0 _108_
rlabel metal2 13468 10108 13468 10108 0 _109_
rlabel metal2 13524 9744 13524 9744 0 _110_
rlabel metal2 14700 9436 14700 9436 0 _111_
rlabel metal2 9604 10836 9604 10836 0 _112_
rlabel metal2 13860 9072 13860 9072 0 _113_
rlabel metal2 14196 9212 14196 9212 0 _114_
rlabel metal2 8708 7840 8708 7840 0 _115_
rlabel metal2 8372 12880 8372 12880 0 _116_
rlabel metal3 8232 13468 8232 13468 0 _117_
rlabel metal3 1239 13468 1239 13468 0 clk
rlabel metal2 12600 10332 12600 10332 0 clknet_0_clk
rlabel metal2 10276 13720 10276 13720 0 clknet_1_0__leaf_clk
rlabel metal2 14028 10976 14028 10976 0 clknet_1_1__leaf_clk
rlabel metal2 8344 9268 8344 9268 0 dut21.count\[0\]
rlabel metal2 9884 7252 9884 7252 0 dut21.count\[1\]
rlabel metal3 10976 11900 10976 11900 0 dut21.count\[2\]
rlabel metal2 12740 11004 12740 11004 0 dut21.count\[3\]
rlabel metal2 8260 14056 8260 14056 0 net1
rlabel metal2 14140 8848 14140 8848 0 net10
rlabel metal2 15484 9324 15484 9324 0 net11
rlabel metal2 2156 11648 2156 11648 0 net12
rlabel metal2 6916 12124 6916 12124 0 net13
rlabel metal2 2044 11732 2044 11732 0 net14
rlabel metal2 8540 2982 8540 2982 0 net15
rlabel metal2 10836 2982 10836 2982 0 net16
rlabel metal2 8428 14994 8428 14994 0 net17
rlabel metal2 14980 12292 14980 12292 0 net18
rlabel metal3 12908 13580 12908 13580 0 net19
rlabel metal2 6748 12768 6748 12768 0 net2
rlabel metal2 15484 10556 15484 10556 0 net20
rlabel metal3 11872 13468 11872 13468 0 net21
rlabel metal2 5572 8596 5572 8596 0 net22
rlabel metal2 9548 13580 9548 13580 0 net23
rlabel metal2 14532 7224 14532 7224 0 net24
rlabel metal2 12292 2982 12292 2982 0 net25
rlabel metal2 12908 3374 12908 3374 0 net26
rlabel metal2 12572 6188 12572 6188 0 net3
rlabel metal2 13972 11312 13972 11312 0 net4
rlabel metal2 10444 13832 10444 13832 0 net5
rlabel metal2 5012 10388 5012 10388 0 net6
rlabel metal2 15288 8372 15288 8372 0 net7
rlabel metal2 14252 13468 14252 13468 0 net8
rlabel metal2 4956 9632 4956 9632 0 net9
rlabel metal2 7756 19481 7756 19481 0 segm[0]
rlabel metal3 679 12460 679 12460 0 segm[10]
rlabel metal2 12460 1211 12460 1211 0 segm[11]
rlabel metal2 20020 11900 20020 11900 0 segm[12]
rlabel metal2 10444 19873 10444 19873 0 segm[13]
rlabel metal3 679 10444 679 10444 0 segm[1]
rlabel metal2 20020 8400 20020 8400 0 segm[2]
rlabel metal3 20321 13804 20321 13804 0 segm[3]
rlabel metal3 679 9772 679 9772 0 segm[4]
rlabel metal2 20020 8820 20020 8820 0 segm[5]
rlabel metal2 20020 10276 20020 10276 0 segm[6]
rlabel metal3 679 11452 679 11452 0 segm[7]
rlabel metal3 679 12124 679 12124 0 segm[8]
rlabel metal3 679 11788 679 11788 0 segm[9]
rlabel metal2 8428 1043 8428 1043 0 sel[0]
rlabel metal2 10780 1099 10780 1099 0 sel[10]
rlabel metal2 8092 19873 8092 19873 0 sel[11]
rlabel metal2 20020 12628 20020 12628 0 sel[1]
rlabel metal2 13132 19677 13132 19677 0 sel[2]
rlabel metal2 20020 11004 20020 11004 0 sel[3]
rlabel metal2 12124 19873 12124 19873 0 sel[4]
rlabel metal3 679 8428 679 8428 0 sel[5]
rlabel metal3 9744 18732 9744 18732 0 sel[6]
rlabel metal2 20020 7504 20020 7504 0 sel[7]
rlabel metal2 11788 1099 11788 1099 0 sel[8]
rlabel metal2 12796 791 12796 791 0 sel[9]
<< properties >>
string FIXED_BBOX 0 0 21000 21000
<< end >>
