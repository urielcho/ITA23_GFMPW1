magic
tech gf180mcuD
magscale 1 5
timestamp 1699641266
<< metal1 >>
rect 672 19221 20328 19238
rect 672 19195 2239 19221
rect 2265 19195 2291 19221
rect 2317 19195 2343 19221
rect 2369 19195 17599 19221
rect 17625 19195 17651 19221
rect 17677 19195 17703 19221
rect 17729 19195 20328 19221
rect 672 19178 20328 19195
rect 9311 19137 9337 19143
rect 9311 19105 9337 19111
rect 11215 19137 11241 19143
rect 11215 19105 11241 19111
rect 12783 19137 12809 19143
rect 12783 19105 12809 19111
rect 14687 19137 14713 19143
rect 14687 19105 14713 19111
rect 8913 18999 8919 19025
rect 8945 18999 8951 19025
rect 10873 18999 10879 19025
rect 10905 18999 10911 19025
rect 12273 18999 12279 19025
rect 12305 18999 12311 19025
rect 14289 18999 14295 19025
rect 14321 18999 14327 19025
rect 672 18829 20328 18846
rect 672 18803 9919 18829
rect 9945 18803 9971 18829
rect 9997 18803 10023 18829
rect 10049 18803 20328 18829
rect 672 18786 20328 18803
rect 10039 18745 10065 18751
rect 10039 18713 10065 18719
rect 13399 18745 13425 18751
rect 13399 18713 13425 18719
rect 9529 18607 9535 18633
rect 9561 18607 9567 18633
rect 12945 18607 12951 18633
rect 12977 18607 12983 18633
rect 672 18437 20328 18454
rect 672 18411 2239 18437
rect 2265 18411 2291 18437
rect 2317 18411 2343 18437
rect 2369 18411 17599 18437
rect 17625 18411 17651 18437
rect 17677 18411 17703 18437
rect 17729 18411 20328 18437
rect 672 18394 20328 18411
rect 8359 18353 8385 18359
rect 8359 18321 8385 18327
rect 7849 18215 7855 18241
rect 7881 18215 7887 18241
rect 672 18045 20328 18062
rect 672 18019 9919 18045
rect 9945 18019 9971 18045
rect 9997 18019 10023 18045
rect 10049 18019 20328 18045
rect 672 18002 20328 18019
rect 672 17653 20328 17670
rect 672 17627 2239 17653
rect 2265 17627 2291 17653
rect 2317 17627 2343 17653
rect 2369 17627 17599 17653
rect 17625 17627 17651 17653
rect 17677 17627 17703 17653
rect 17729 17627 20328 17653
rect 672 17610 20328 17627
rect 672 17261 20328 17278
rect 672 17235 9919 17261
rect 9945 17235 9971 17261
rect 9997 17235 10023 17261
rect 10049 17235 20328 17261
rect 672 17218 20328 17235
rect 672 16869 20328 16886
rect 672 16843 2239 16869
rect 2265 16843 2291 16869
rect 2317 16843 2343 16869
rect 2369 16843 17599 16869
rect 17625 16843 17651 16869
rect 17677 16843 17703 16869
rect 17729 16843 20328 16869
rect 672 16826 20328 16843
rect 672 16477 20328 16494
rect 672 16451 9919 16477
rect 9945 16451 9971 16477
rect 9997 16451 10023 16477
rect 10049 16451 20328 16477
rect 672 16434 20328 16451
rect 672 16085 20328 16102
rect 672 16059 2239 16085
rect 2265 16059 2291 16085
rect 2317 16059 2343 16085
rect 2369 16059 17599 16085
rect 17625 16059 17651 16085
rect 17677 16059 17703 16085
rect 17729 16059 20328 16085
rect 672 16042 20328 16059
rect 672 15693 20328 15710
rect 672 15667 9919 15693
rect 9945 15667 9971 15693
rect 9997 15667 10023 15693
rect 10049 15667 20328 15693
rect 672 15650 20328 15667
rect 672 15301 20328 15318
rect 672 15275 2239 15301
rect 2265 15275 2291 15301
rect 2317 15275 2343 15301
rect 2369 15275 17599 15301
rect 17625 15275 17651 15301
rect 17677 15275 17703 15301
rect 17729 15275 20328 15301
rect 672 15258 20328 15275
rect 672 14909 20328 14926
rect 672 14883 9919 14909
rect 9945 14883 9971 14909
rect 9997 14883 10023 14909
rect 10049 14883 20328 14909
rect 672 14866 20328 14883
rect 672 14517 20328 14534
rect 672 14491 2239 14517
rect 2265 14491 2291 14517
rect 2317 14491 2343 14517
rect 2369 14491 17599 14517
rect 17625 14491 17651 14517
rect 17677 14491 17703 14517
rect 17729 14491 20328 14517
rect 672 14474 20328 14491
rect 10935 14321 10961 14327
rect 10935 14289 10961 14295
rect 10879 14209 10905 14215
rect 10879 14177 10905 14183
rect 672 14125 20328 14142
rect 672 14099 9919 14125
rect 9945 14099 9971 14125
rect 9997 14099 10023 14125
rect 10049 14099 20328 14125
rect 672 14082 20328 14099
rect 12951 14041 12977 14047
rect 13113 14015 13119 14041
rect 13145 14015 13151 14041
rect 12951 14009 12977 14015
rect 12671 13985 12697 13991
rect 10593 13959 10599 13985
rect 10625 13959 10631 13985
rect 12671 13953 12697 13959
rect 11943 13929 11969 13935
rect 6225 13903 6231 13929
rect 6257 13903 6263 13929
rect 10257 13903 10263 13929
rect 10289 13903 10295 13929
rect 11943 13897 11969 13903
rect 7911 13873 7937 13879
rect 6561 13847 6567 13873
rect 6593 13847 6599 13873
rect 7625 13847 7631 13873
rect 7657 13847 7663 13873
rect 11657 13847 11663 13873
rect 11689 13847 11695 13873
rect 7911 13841 7937 13847
rect 12615 13817 12641 13823
rect 12615 13785 12641 13791
rect 672 13733 20328 13750
rect 672 13707 2239 13733
rect 2265 13707 2291 13733
rect 2317 13707 2343 13733
rect 2369 13707 17599 13733
rect 17625 13707 17651 13733
rect 17677 13707 17703 13733
rect 17729 13707 20328 13733
rect 672 13690 20328 13707
rect 7127 13649 7153 13655
rect 7127 13617 7153 13623
rect 10711 13593 10737 13599
rect 20007 13593 20033 13599
rect 8913 13567 8919 13593
rect 8945 13567 8951 13593
rect 13169 13567 13175 13593
rect 13201 13567 13207 13593
rect 10711 13561 10737 13567
rect 20007 13561 20033 13567
rect 9031 13537 9057 13543
rect 10375 13537 10401 13543
rect 7457 13511 7463 13537
rect 7489 13511 7495 13537
rect 9193 13511 9199 13537
rect 9225 13511 9231 13537
rect 9031 13505 9057 13511
rect 10375 13505 10401 13511
rect 10823 13537 10849 13543
rect 10823 13505 10849 13511
rect 11327 13537 11353 13543
rect 11327 13505 11353 13511
rect 11439 13537 11465 13543
rect 11439 13505 11465 13511
rect 11551 13537 11577 13543
rect 13399 13537 13425 13543
rect 11769 13511 11775 13537
rect 11801 13511 11807 13537
rect 18825 13511 18831 13537
rect 18857 13511 18863 13537
rect 11551 13505 11577 13511
rect 13399 13505 13425 13511
rect 7183 13481 7209 13487
rect 9311 13481 9337 13487
rect 7849 13455 7855 13481
rect 7881 13455 7887 13481
rect 7183 13449 7209 13455
rect 9311 13449 9337 13455
rect 10207 13481 10233 13487
rect 10207 13449 10233 13455
rect 10655 13481 10681 13487
rect 10655 13449 10681 13455
rect 10935 13481 10961 13487
rect 10935 13449 10961 13455
rect 11103 13481 11129 13487
rect 11209 13455 11215 13481
rect 11241 13455 11247 13481
rect 12105 13455 12111 13481
rect 12137 13455 12143 13481
rect 11103 13449 11129 13455
rect 9367 13425 9393 13431
rect 9367 13393 9393 13399
rect 9535 13425 9561 13431
rect 9535 13393 9561 13399
rect 10319 13425 10345 13431
rect 10319 13393 10345 13399
rect 11607 13425 11633 13431
rect 11607 13393 11633 13399
rect 672 13341 20328 13358
rect 672 13315 9919 13341
rect 9945 13315 9971 13341
rect 9997 13315 10023 13341
rect 10049 13315 20328 13341
rect 672 13298 20328 13315
rect 8919 13257 8945 13263
rect 14295 13257 14321 13263
rect 11825 13231 11831 13257
rect 11857 13231 11863 13257
rect 8919 13225 8945 13231
rect 14295 13225 14321 13231
rect 7911 13201 7937 13207
rect 7911 13169 7937 13175
rect 8079 13201 8105 13207
rect 9977 13175 9983 13201
rect 10009 13175 10015 13201
rect 11769 13175 11775 13201
rect 11801 13175 11807 13201
rect 12105 13175 12111 13201
rect 12137 13175 12143 13201
rect 8079 13169 8105 13175
rect 7687 13145 7713 13151
rect 8415 13145 8441 13151
rect 2137 13119 2143 13145
rect 2169 13119 2175 13145
rect 5609 13119 5615 13145
rect 5641 13119 5647 13145
rect 8017 13119 8023 13145
rect 8049 13119 8055 13145
rect 8185 13119 8191 13145
rect 8217 13119 8223 13145
rect 7687 13113 7713 13119
rect 8415 13113 8441 13119
rect 8695 13145 8721 13151
rect 9087 13145 9113 13151
rect 9025 13119 9031 13145
rect 9057 13119 9063 13145
rect 9193 13119 9199 13145
rect 9225 13119 9231 13145
rect 9585 13119 9591 13145
rect 9617 13119 9623 13145
rect 11265 13119 11271 13145
rect 11297 13119 11303 13145
rect 11713 13119 11719 13145
rect 11745 13119 11751 13145
rect 12217 13119 12223 13145
rect 12249 13119 12255 13145
rect 12609 13119 12615 13145
rect 12641 13119 12647 13145
rect 8695 13113 8721 13119
rect 9087 13113 9113 13119
rect 7239 13089 7265 13095
rect 5945 13063 5951 13089
rect 5977 13063 5983 13089
rect 7009 13063 7015 13089
rect 7041 13063 7047 13089
rect 7239 13057 7265 13063
rect 9423 13089 9449 13095
rect 11041 13063 11047 13089
rect 11073 13063 11079 13089
rect 13001 13063 13007 13089
rect 13033 13063 13039 13089
rect 14065 13063 14071 13089
rect 14097 13063 14103 13089
rect 9423 13057 9449 13063
rect 967 13033 993 13039
rect 967 13001 993 13007
rect 7743 13033 7769 13039
rect 7743 13001 7769 13007
rect 8359 13033 8385 13039
rect 8359 13001 8385 13007
rect 8751 13033 8777 13039
rect 8751 13001 8777 13007
rect 672 12949 20328 12966
rect 672 12923 2239 12949
rect 2265 12923 2291 12949
rect 2317 12923 2343 12949
rect 2369 12923 17599 12949
rect 17625 12923 17651 12949
rect 17677 12923 17703 12949
rect 17729 12923 20328 12949
rect 672 12906 20328 12923
rect 10319 12865 10345 12871
rect 10319 12833 10345 12839
rect 10655 12865 10681 12871
rect 10655 12833 10681 12839
rect 7575 12809 7601 12815
rect 7575 12777 7601 12783
rect 7799 12809 7825 12815
rect 12279 12809 12305 12815
rect 9697 12783 9703 12809
rect 9729 12783 9735 12809
rect 10817 12783 10823 12809
rect 10849 12783 10855 12809
rect 7799 12777 7825 12783
rect 12279 12777 12305 12783
rect 7463 12753 7489 12759
rect 7463 12721 7489 12727
rect 7743 12753 7769 12759
rect 11159 12753 11185 12759
rect 8241 12727 8247 12753
rect 8273 12727 8279 12753
rect 7743 12721 7769 12727
rect 11159 12721 11185 12727
rect 12055 12753 12081 12759
rect 12055 12721 12081 12727
rect 12335 12753 12361 12759
rect 12335 12721 12361 12727
rect 13175 12753 13201 12759
rect 13175 12721 13201 12727
rect 6231 12697 6257 12703
rect 6231 12665 6257 12671
rect 6399 12697 6425 12703
rect 10375 12697 10401 12703
rect 12167 12697 12193 12703
rect 7289 12671 7295 12697
rect 7321 12671 7327 12697
rect 8633 12671 8639 12697
rect 8665 12671 8671 12697
rect 10985 12671 10991 12697
rect 11017 12671 11023 12697
rect 6399 12665 6425 12671
rect 10375 12665 10401 12671
rect 12167 12665 12193 12671
rect 13287 12697 13313 12703
rect 13287 12665 13313 12671
rect 13343 12697 13369 12703
rect 13343 12665 13369 12671
rect 9927 12641 9953 12647
rect 9927 12609 9953 12615
rect 10319 12641 10345 12647
rect 10319 12609 10345 12615
rect 10767 12641 10793 12647
rect 10767 12609 10793 12615
rect 672 12557 20328 12574
rect 672 12531 9919 12557
rect 9945 12531 9971 12557
rect 9997 12531 10023 12557
rect 10049 12531 20328 12557
rect 672 12514 20328 12531
rect 7575 12473 7601 12479
rect 7575 12441 7601 12447
rect 7631 12473 7657 12479
rect 7631 12441 7657 12447
rect 9087 12473 9113 12479
rect 9087 12441 9113 12447
rect 9143 12473 9169 12479
rect 13679 12473 13705 12479
rect 10705 12447 10711 12473
rect 10737 12447 10743 12473
rect 9143 12441 9169 12447
rect 13679 12441 13705 12447
rect 7519 12361 7545 12367
rect 7519 12329 7545 12335
rect 7855 12361 7881 12367
rect 7855 12329 7881 12335
rect 9031 12361 9057 12367
rect 9031 12329 9057 12335
rect 9367 12361 9393 12367
rect 10817 12335 10823 12361
rect 10849 12335 10855 12361
rect 13841 12335 13847 12361
rect 13873 12335 13879 12361
rect 18825 12335 18831 12361
rect 18857 12335 18863 12361
rect 9367 12329 9393 12335
rect 14233 12279 14239 12305
rect 14265 12279 14271 12305
rect 15297 12279 15303 12305
rect 15329 12279 15335 12305
rect 20007 12249 20033 12255
rect 20007 12217 20033 12223
rect 672 12165 20328 12182
rect 672 12139 2239 12165
rect 2265 12139 2291 12165
rect 2317 12139 2343 12165
rect 2369 12139 17599 12165
rect 17625 12139 17651 12165
rect 17677 12139 17703 12165
rect 17729 12139 20328 12165
rect 672 12122 20328 12139
rect 7127 12081 7153 12087
rect 7127 12049 7153 12055
rect 967 12025 993 12031
rect 11831 12025 11857 12031
rect 6953 11999 6959 12025
rect 6985 11999 6991 12025
rect 967 11993 993 11999
rect 11831 11993 11857 11999
rect 13455 12025 13481 12031
rect 13455 11993 13481 11999
rect 20007 12025 20033 12031
rect 20007 11993 20033 11999
rect 11943 11969 11969 11975
rect 2137 11943 2143 11969
rect 2169 11943 2175 11969
rect 8689 11943 8695 11969
rect 8721 11943 8727 11969
rect 10761 11943 10767 11969
rect 10793 11943 10799 11969
rect 11943 11937 11969 11943
rect 13959 11969 13985 11975
rect 18825 11943 18831 11969
rect 18857 11943 18863 11969
rect 13959 11937 13985 11943
rect 7015 11913 7041 11919
rect 7015 11881 7041 11887
rect 8583 11913 8609 11919
rect 12279 11913 12305 11919
rect 10873 11887 10879 11913
rect 10905 11887 10911 11913
rect 11153 11887 11159 11913
rect 11185 11887 11191 11913
rect 12105 11887 12111 11913
rect 12137 11887 12143 11913
rect 8583 11881 8609 11887
rect 12279 11881 12305 11887
rect 7631 11857 7657 11863
rect 12447 11857 12473 11863
rect 11209 11831 11215 11857
rect 11241 11831 11247 11857
rect 7631 11825 7657 11831
rect 12447 11825 12473 11831
rect 13847 11857 13873 11863
rect 13847 11825 13873 11831
rect 13903 11857 13929 11863
rect 13903 11825 13929 11831
rect 14071 11857 14097 11863
rect 14071 11825 14097 11831
rect 672 11773 20328 11790
rect 672 11747 9919 11773
rect 9945 11747 9971 11773
rect 9997 11747 10023 11773
rect 10049 11747 20328 11773
rect 672 11730 20328 11747
rect 9759 11689 9785 11695
rect 9305 11663 9311 11689
rect 9337 11663 9343 11689
rect 9759 11657 9785 11663
rect 11831 11689 11857 11695
rect 11831 11657 11857 11663
rect 13287 11689 13313 11695
rect 13287 11657 13313 11663
rect 9647 11633 9673 11639
rect 9647 11601 9673 11607
rect 9871 11633 9897 11639
rect 9871 11601 9897 11607
rect 10543 11633 10569 11639
rect 11943 11633 11969 11639
rect 11041 11607 11047 11633
rect 11073 11607 11079 11633
rect 10543 11601 10569 11607
rect 11943 11601 11969 11607
rect 11999 11633 12025 11639
rect 11999 11601 12025 11607
rect 13399 11633 13425 11639
rect 13399 11601 13425 11607
rect 13455 11633 13481 11639
rect 15409 11607 15415 11633
rect 15441 11607 15447 11633
rect 13455 11601 13481 11607
rect 2137 11551 2143 11577
rect 2169 11551 2175 11577
rect 7513 11557 7519 11583
rect 7545 11557 7551 11583
rect 7687 11577 7713 11583
rect 7687 11545 7713 11551
rect 7799 11577 7825 11583
rect 7799 11545 7825 11551
rect 7967 11577 7993 11583
rect 7967 11545 7993 11551
rect 9479 11577 9505 11583
rect 11439 11577 11465 11583
rect 10313 11551 10319 11577
rect 10345 11551 10351 11577
rect 10705 11551 10711 11577
rect 10737 11551 10743 11577
rect 10985 11551 10991 11577
rect 11017 11551 11023 11577
rect 9479 11545 9505 11551
rect 11439 11545 11465 11551
rect 12895 11577 12921 11583
rect 15247 11577 15273 11583
rect 13113 11551 13119 11577
rect 13145 11551 13151 11577
rect 13617 11551 13623 11577
rect 13649 11551 13655 11577
rect 18825 11551 18831 11577
rect 18857 11551 18863 11577
rect 12895 11545 12921 11551
rect 15247 11545 15273 11551
rect 7743 11521 7769 11527
rect 6057 11495 6063 11521
rect 6089 11495 6095 11521
rect 7121 11495 7127 11521
rect 7153 11495 7159 11521
rect 10089 11495 10095 11521
rect 10121 11495 10127 11521
rect 11209 11495 11215 11521
rect 11241 11495 11247 11521
rect 11657 11495 11663 11521
rect 11689 11495 11695 11521
rect 14009 11495 14015 11521
rect 14041 11495 14047 11521
rect 15073 11495 15079 11521
rect 15105 11495 15111 11521
rect 7743 11489 7769 11495
rect 967 11465 993 11471
rect 967 11433 993 11439
rect 9591 11465 9617 11471
rect 9591 11433 9617 11439
rect 20007 11465 20033 11471
rect 20007 11433 20033 11439
rect 672 11381 20328 11398
rect 672 11355 2239 11381
rect 2265 11355 2291 11381
rect 2317 11355 2343 11381
rect 2369 11355 17599 11381
rect 17625 11355 17651 11381
rect 17677 11355 17703 11381
rect 17729 11355 20328 11381
rect 672 11338 20328 11355
rect 7631 11297 7657 11303
rect 7631 11265 7657 11271
rect 14183 11297 14209 11303
rect 14183 11265 14209 11271
rect 10375 11241 10401 11247
rect 7513 11215 7519 11241
rect 7545 11215 7551 11241
rect 9193 11215 9199 11241
rect 9225 11215 9231 11241
rect 10375 11209 10401 11215
rect 11719 11241 11745 11247
rect 13903 11241 13929 11247
rect 12441 11215 12447 11241
rect 12473 11215 12479 11241
rect 13505 11215 13511 11241
rect 13537 11215 13543 11241
rect 11719 11209 11745 11215
rect 13903 11209 13929 11215
rect 6847 11185 6873 11191
rect 6847 11153 6873 11159
rect 6959 11185 6985 11191
rect 8751 11185 8777 11191
rect 10095 11185 10121 11191
rect 8353 11159 8359 11185
rect 8385 11159 8391 11185
rect 9081 11159 9087 11185
rect 9113 11159 9119 11185
rect 9473 11159 9479 11185
rect 9505 11159 9511 11185
rect 6959 11153 6985 11159
rect 8751 11153 8777 11159
rect 10095 11153 10121 11159
rect 10935 11185 10961 11191
rect 10935 11153 10961 11159
rect 11103 11185 11129 11191
rect 13791 11185 13817 11191
rect 11769 11159 11775 11185
rect 11801 11159 11807 11185
rect 12105 11159 12111 11185
rect 12137 11159 12143 11185
rect 11103 11153 11129 11159
rect 13791 11153 13817 11159
rect 14015 11185 14041 11191
rect 14015 11153 14041 11159
rect 7519 11129 7545 11135
rect 13679 11129 13705 11135
rect 8577 11103 8583 11129
rect 8609 11103 8615 11129
rect 8913 11103 8919 11129
rect 8945 11103 8951 11129
rect 7519 11097 7545 11103
rect 13679 11097 13705 11103
rect 14127 11129 14153 11135
rect 14127 11097 14153 11103
rect 14183 11129 14209 11135
rect 14183 11097 14209 11103
rect 6903 11073 6929 11079
rect 6903 11041 6929 11047
rect 7071 11073 7097 11079
rect 10655 11073 10681 11079
rect 8241 11047 8247 11073
rect 8273 11047 8279 11073
rect 7071 11041 7097 11047
rect 10655 11041 10681 11047
rect 11383 11073 11409 11079
rect 11383 11041 11409 11047
rect 11551 11073 11577 11079
rect 11551 11041 11577 11047
rect 11663 11073 11689 11079
rect 11663 11041 11689 11047
rect 672 10989 20328 11006
rect 672 10963 9919 10989
rect 9945 10963 9971 10989
rect 9997 10963 10023 10989
rect 10049 10963 20328 10989
rect 672 10946 20328 10963
rect 8751 10905 8777 10911
rect 8751 10873 8777 10879
rect 8807 10905 8833 10911
rect 13063 10905 13089 10911
rect 9697 10879 9703 10905
rect 9729 10879 9735 10905
rect 10145 10879 10151 10905
rect 10177 10879 10183 10905
rect 10593 10879 10599 10905
rect 10625 10879 10631 10905
rect 8807 10873 8833 10879
rect 13063 10873 13089 10879
rect 13791 10905 13817 10911
rect 13791 10873 13817 10879
rect 14015 10905 14041 10911
rect 14015 10873 14041 10879
rect 13287 10849 13313 10855
rect 6617 10823 6623 10849
rect 6649 10823 6655 10849
rect 8409 10823 8415 10849
rect 8441 10823 8447 10849
rect 9361 10823 9367 10849
rect 9393 10823 9399 10849
rect 9641 10823 9647 10849
rect 9673 10823 9679 10849
rect 10649 10823 10655 10849
rect 10681 10823 10687 10849
rect 13287 10817 13313 10823
rect 13511 10849 13537 10855
rect 13511 10817 13537 10823
rect 13567 10849 13593 10855
rect 13567 10817 13593 10823
rect 9087 10793 9113 10799
rect 7009 10767 7015 10793
rect 7041 10767 7047 10793
rect 8297 10767 8303 10793
rect 8329 10767 8335 10793
rect 8913 10767 8919 10793
rect 8945 10767 8951 10793
rect 9087 10761 9113 10767
rect 9759 10793 9785 10799
rect 9759 10761 9785 10767
rect 10319 10793 10345 10799
rect 13231 10793 13257 10799
rect 10593 10767 10599 10793
rect 10625 10767 10631 10793
rect 12049 10767 12055 10793
rect 12081 10767 12087 10793
rect 12329 10767 12335 10793
rect 12361 10767 12367 10793
rect 10319 10761 10345 10767
rect 13231 10761 13257 10767
rect 7239 10737 7265 10743
rect 5553 10711 5559 10737
rect 5585 10711 5591 10737
rect 7239 10705 7265 10711
rect 12783 10737 12809 10743
rect 12783 10705 12809 10711
rect 13287 10681 13313 10687
rect 13287 10649 13313 10655
rect 672 10597 20328 10614
rect 672 10571 2239 10597
rect 2265 10571 2291 10597
rect 2317 10571 2343 10597
rect 2369 10571 17599 10597
rect 17625 10571 17651 10597
rect 17677 10571 17703 10597
rect 17729 10571 20328 10597
rect 672 10554 20328 10571
rect 11439 10513 11465 10519
rect 11439 10481 11465 10487
rect 7351 10457 7377 10463
rect 11495 10457 11521 10463
rect 7065 10431 7071 10457
rect 7097 10431 7103 10457
rect 7849 10431 7855 10457
rect 7881 10431 7887 10457
rect 13729 10431 13735 10457
rect 13761 10431 13767 10457
rect 7351 10425 7377 10431
rect 11495 10425 11521 10431
rect 11215 10401 11241 10407
rect 10033 10375 10039 10401
rect 10065 10375 10071 10401
rect 11215 10369 11241 10375
rect 11271 10401 11297 10407
rect 11657 10375 11663 10401
rect 11689 10375 11695 10401
rect 11271 10369 11297 10375
rect 10817 10319 10823 10345
rect 10849 10319 10855 10345
rect 11097 10319 11103 10345
rect 11129 10319 11135 10345
rect 6847 10289 6873 10295
rect 6847 10257 6873 10263
rect 672 10205 20328 10222
rect 672 10179 9919 10205
rect 9945 10179 9971 10205
rect 9997 10179 10023 10205
rect 10049 10179 20328 10205
rect 672 10162 20328 10179
rect 13791 10065 13817 10071
rect 6001 10039 6007 10065
rect 6033 10039 6039 10065
rect 7401 10039 7407 10065
rect 7433 10039 7439 10065
rect 7737 10039 7743 10065
rect 7769 10039 7775 10065
rect 8185 10039 8191 10065
rect 8217 10039 8223 10065
rect 11041 10039 11047 10065
rect 11073 10039 11079 10065
rect 13393 10039 13399 10065
rect 13425 10039 13431 10065
rect 13791 10033 13817 10039
rect 7239 10009 7265 10015
rect 5609 9983 5615 10009
rect 5641 9983 5647 10009
rect 7239 9977 7265 9983
rect 7575 10009 7601 10015
rect 7575 9977 7601 9983
rect 8023 10009 8049 10015
rect 8023 9977 8049 9983
rect 9143 10009 9169 10015
rect 13847 10009 13873 10015
rect 9249 9983 9255 10009
rect 9281 9983 9287 10009
rect 9697 9983 9703 10009
rect 9729 9983 9735 10009
rect 12721 9983 12727 10009
rect 12753 9983 12759 10009
rect 13113 9983 13119 10009
rect 13145 9983 13151 10009
rect 14009 9983 14015 10009
rect 14041 9983 14047 10009
rect 18825 9983 18831 10009
rect 18857 9983 18863 10009
rect 9143 9977 9169 9983
rect 13847 9977 13873 9983
rect 7911 9953 7937 9959
rect 7065 9927 7071 9953
rect 7097 9927 7103 9953
rect 7911 9921 7937 9927
rect 8751 9953 8777 9959
rect 9081 9927 9087 9953
rect 9113 9927 9119 9953
rect 13057 9927 13063 9953
rect 13089 9927 13095 9953
rect 14401 9927 14407 9953
rect 14433 9927 14439 9953
rect 15465 9927 15471 9953
rect 15497 9927 15503 9953
rect 8751 9921 8777 9927
rect 13791 9897 13817 9903
rect 9249 9871 9255 9897
rect 9281 9871 9287 9897
rect 13791 9865 13817 9871
rect 20007 9897 20033 9903
rect 20007 9865 20033 9871
rect 672 9813 20328 9830
rect 672 9787 2239 9813
rect 2265 9787 2291 9813
rect 2317 9787 2343 9813
rect 2369 9787 17599 9813
rect 17625 9787 17651 9813
rect 17677 9787 17703 9813
rect 17729 9787 20328 9813
rect 672 9770 20328 9787
rect 8639 9729 8665 9735
rect 8639 9697 8665 9703
rect 10711 9729 10737 9735
rect 13287 9729 13313 9735
rect 11601 9703 11607 9729
rect 11633 9703 11639 9729
rect 10711 9697 10737 9703
rect 13287 9697 13313 9703
rect 13679 9729 13705 9735
rect 13679 9697 13705 9703
rect 15079 9729 15105 9735
rect 15079 9697 15105 9703
rect 6735 9673 6761 9679
rect 14127 9673 14153 9679
rect 6897 9647 6903 9673
rect 6929 9647 6935 9673
rect 10985 9647 10991 9673
rect 11017 9647 11023 9673
rect 11881 9647 11887 9673
rect 11913 9647 11919 9673
rect 6735 9641 6761 9647
rect 14127 9641 14153 9647
rect 14799 9673 14825 9679
rect 14799 9641 14825 9647
rect 20007 9673 20033 9679
rect 20007 9641 20033 9647
rect 7967 9617 7993 9623
rect 8975 9617 9001 9623
rect 7065 9591 7071 9617
rect 7097 9591 7103 9617
rect 7737 9591 7743 9617
rect 7769 9591 7775 9617
rect 8409 9591 8415 9617
rect 8441 9591 8447 9617
rect 8801 9591 8807 9617
rect 8833 9591 8839 9617
rect 7967 9585 7993 9591
rect 8975 9585 9001 9591
rect 10039 9617 10065 9623
rect 10039 9585 10065 9591
rect 10375 9617 10401 9623
rect 11383 9617 11409 9623
rect 13175 9617 13201 9623
rect 13623 9617 13649 9623
rect 11153 9591 11159 9617
rect 11185 9591 11191 9617
rect 11825 9591 11831 9617
rect 11857 9591 11863 9617
rect 12217 9591 12223 9617
rect 12249 9591 12255 9617
rect 12945 9591 12951 9617
rect 12977 9591 12983 9617
rect 13449 9591 13455 9617
rect 13481 9591 13487 9617
rect 10375 9585 10401 9591
rect 11383 9585 11409 9591
rect 13175 9585 13201 9591
rect 13623 9585 13649 9591
rect 14575 9617 14601 9623
rect 14575 9585 14601 9591
rect 14911 9617 14937 9623
rect 18825 9591 18831 9617
rect 18857 9591 18863 9617
rect 14911 9585 14937 9591
rect 10655 9561 10681 9567
rect 8521 9535 8527 9561
rect 8553 9535 8559 9561
rect 10655 9529 10681 9535
rect 13959 9561 13985 9567
rect 13959 9529 13985 9535
rect 14071 9561 14097 9567
rect 14071 9529 14097 9535
rect 14183 9561 14209 9567
rect 14183 9529 14209 9535
rect 14687 9561 14713 9567
rect 14687 9529 14713 9535
rect 15023 9561 15049 9567
rect 15023 9529 15049 9535
rect 8695 9505 8721 9511
rect 9311 9505 9337 9511
rect 9647 9505 9673 9511
rect 13679 9505 13705 9511
rect 9137 9479 9143 9505
rect 9169 9479 9175 9505
rect 9473 9479 9479 9505
rect 9505 9479 9511 9505
rect 9865 9479 9871 9505
rect 9897 9479 9903 9505
rect 10201 9479 10207 9505
rect 10233 9479 10239 9505
rect 12105 9479 12111 9505
rect 12137 9479 12143 9505
rect 12833 9479 12839 9505
rect 12865 9479 12871 9505
rect 8695 9473 8721 9479
rect 9311 9473 9337 9479
rect 9647 9473 9673 9479
rect 13679 9473 13705 9479
rect 14239 9505 14265 9511
rect 14239 9473 14265 9479
rect 15079 9505 15105 9511
rect 15079 9473 15105 9479
rect 672 9421 20328 9438
rect 672 9395 9919 9421
rect 9945 9395 9971 9421
rect 9997 9395 10023 9421
rect 10049 9395 20328 9421
rect 672 9378 20328 9395
rect 8023 9337 8049 9343
rect 8023 9305 8049 9311
rect 8639 9337 8665 9343
rect 8639 9305 8665 9311
rect 10431 9337 10457 9343
rect 11825 9311 11831 9337
rect 11857 9311 11863 9337
rect 10431 9305 10457 9311
rect 8185 9255 8191 9281
rect 8217 9255 8223 9281
rect 10873 9255 10879 9281
rect 10905 9255 10911 9281
rect 14233 9255 14239 9281
rect 14265 9255 14271 9281
rect 7183 9225 7209 9231
rect 9759 9225 9785 9231
rect 5553 9199 5559 9225
rect 5585 9199 5591 9225
rect 8857 9199 8863 9225
rect 8889 9199 8895 9225
rect 8969 9199 8975 9225
rect 9001 9199 9007 9225
rect 7183 9193 7209 9199
rect 9759 9193 9785 9199
rect 9871 9225 9897 9231
rect 11439 9225 11465 9231
rect 10985 9199 10991 9225
rect 11017 9199 11023 9225
rect 9871 9193 9897 9199
rect 11439 9193 11465 9199
rect 11495 9225 11521 9231
rect 11495 9193 11521 9199
rect 11719 9225 11745 9231
rect 11937 9199 11943 9225
rect 11969 9199 11975 9225
rect 13841 9199 13847 9225
rect 13873 9199 13879 9225
rect 11719 9193 11745 9199
rect 9647 9169 9673 9175
rect 11607 9169 11633 9175
rect 5889 9143 5895 9169
rect 5921 9143 5927 9169
rect 6953 9143 6959 9169
rect 6985 9143 6991 9169
rect 9025 9143 9031 9169
rect 9057 9143 9063 9169
rect 10649 9143 10655 9169
rect 10681 9143 10687 9169
rect 9647 9137 9673 9143
rect 11607 9137 11633 9143
rect 13679 9169 13705 9175
rect 15297 9143 15303 9169
rect 15329 9143 15335 9169
rect 13679 9137 13705 9143
rect 10095 9113 10121 9119
rect 10095 9081 10121 9087
rect 672 9029 20328 9046
rect 672 9003 2239 9029
rect 2265 9003 2291 9029
rect 2317 9003 2343 9029
rect 2369 9003 17599 9029
rect 17625 9003 17651 9029
rect 17677 9003 17703 9029
rect 17729 9003 20328 9029
rect 672 8986 20328 9003
rect 9087 8945 9113 8951
rect 9087 8913 9113 8919
rect 9927 8945 9953 8951
rect 9927 8913 9953 8919
rect 11159 8945 11185 8951
rect 11159 8913 11185 8919
rect 7183 8889 7209 8895
rect 11433 8863 11439 8889
rect 11465 8863 11471 8889
rect 12497 8863 12503 8889
rect 12529 8863 12535 8889
rect 7183 8857 7209 8863
rect 9311 8833 9337 8839
rect 9025 8807 9031 8833
rect 9057 8807 9063 8833
rect 9311 8801 9337 8807
rect 9871 8833 9897 8839
rect 12889 8807 12895 8833
rect 12921 8807 12927 8833
rect 9871 8801 9897 8807
rect 9927 8777 9953 8783
rect 9193 8751 9199 8777
rect 9225 8751 9231 8777
rect 9927 8745 9953 8751
rect 11103 8777 11129 8783
rect 11103 8745 11129 8751
rect 11159 8777 11185 8783
rect 11159 8745 11185 8751
rect 8919 8721 8945 8727
rect 8919 8689 8945 8695
rect 13119 8721 13145 8727
rect 13119 8689 13145 8695
rect 672 8637 20328 8654
rect 672 8611 9919 8637
rect 9945 8611 9971 8637
rect 9997 8611 10023 8637
rect 10049 8611 20328 8637
rect 672 8594 20328 8611
rect 7519 8553 7545 8559
rect 7519 8521 7545 8527
rect 8191 8553 8217 8559
rect 8191 8521 8217 8527
rect 8303 8553 8329 8559
rect 8303 8521 8329 8527
rect 10487 8553 10513 8559
rect 10487 8521 10513 8527
rect 9535 8497 9561 8503
rect 9535 8465 9561 8471
rect 9591 8497 9617 8503
rect 14183 8497 14209 8503
rect 10313 8471 10319 8497
rect 10345 8471 10351 8497
rect 11265 8471 11271 8497
rect 11297 8471 11303 8497
rect 9591 8465 9617 8471
rect 14183 8465 14209 8471
rect 7407 8441 7433 8447
rect 2137 8415 2143 8441
rect 2169 8415 2175 8441
rect 7065 8415 7071 8441
rect 7097 8415 7103 8441
rect 7233 8415 7239 8441
rect 7265 8415 7271 8441
rect 7407 8409 7433 8415
rect 8415 8441 8441 8447
rect 9423 8441 9449 8447
rect 13847 8441 13873 8447
rect 8969 8415 8975 8441
rect 9001 8415 9007 8441
rect 9137 8415 9143 8441
rect 9169 8415 9175 8441
rect 10705 8415 10711 8441
rect 10737 8415 10743 8441
rect 11041 8415 11047 8441
rect 11073 8415 11079 8441
rect 11321 8415 11327 8441
rect 11353 8415 11359 8441
rect 8415 8409 8441 8415
rect 9423 8409 9449 8415
rect 13847 8409 13873 8415
rect 14071 8441 14097 8447
rect 18937 8415 18943 8441
rect 18969 8415 18975 8441
rect 14071 8409 14097 8415
rect 7463 8385 7489 8391
rect 5609 8359 5615 8385
rect 5641 8359 5647 8385
rect 6673 8359 6679 8385
rect 6705 8359 6711 8385
rect 7463 8353 7489 8359
rect 8359 8385 8385 8391
rect 11439 8385 11465 8391
rect 9193 8359 9199 8385
rect 9225 8359 9231 8385
rect 8359 8353 8385 8359
rect 11439 8353 11465 8359
rect 13959 8385 13985 8391
rect 19945 8359 19951 8385
rect 19977 8359 19983 8385
rect 13959 8353 13985 8359
rect 967 8329 993 8335
rect 9249 8303 9255 8329
rect 9281 8303 9287 8329
rect 967 8297 993 8303
rect 672 8245 20328 8262
rect 672 8219 2239 8245
rect 2265 8219 2291 8245
rect 2317 8219 2343 8245
rect 2369 8219 17599 8245
rect 17625 8219 17651 8245
rect 17677 8219 17703 8245
rect 17729 8219 20328 8245
rect 672 8202 20328 8219
rect 6959 8105 6985 8111
rect 9423 8105 9449 8111
rect 1017 8079 1023 8105
rect 1049 8079 1055 8105
rect 7905 8079 7911 8105
rect 7937 8079 7943 8105
rect 8969 8079 8975 8105
rect 9001 8079 9007 8105
rect 6959 8073 6985 8079
rect 9423 8073 9449 8079
rect 20007 8105 20033 8111
rect 20007 8073 20033 8079
rect 6903 8049 6929 8055
rect 2137 8023 2143 8049
rect 2169 8023 2175 8049
rect 6903 8017 6929 8023
rect 7015 8049 7041 8055
rect 9143 8049 9169 8055
rect 9367 8049 9393 8055
rect 7513 8023 7519 8049
rect 7545 8023 7551 8049
rect 9305 8023 9311 8049
rect 9337 8023 9343 8049
rect 7015 8017 7041 8023
rect 9143 8017 9169 8023
rect 9367 8017 9393 8023
rect 9479 8049 9505 8055
rect 9479 8017 9505 8023
rect 11887 8049 11913 8055
rect 11887 8017 11913 8023
rect 11999 8049 12025 8055
rect 11999 8017 12025 8023
rect 13679 8049 13705 8055
rect 13959 8049 13985 8055
rect 13841 8023 13847 8049
rect 13873 8023 13879 8049
rect 13679 8017 13705 8023
rect 13959 8017 13985 8023
rect 14071 8049 14097 8055
rect 14071 8017 14097 8023
rect 14519 8049 14545 8055
rect 14519 8017 14545 8023
rect 14687 8049 14713 8055
rect 14687 8017 14713 8023
rect 14911 8049 14937 8055
rect 18825 8023 18831 8049
rect 18857 8023 18863 8049
rect 14911 8017 14937 8023
rect 11775 7993 11801 7999
rect 11775 7961 11801 7967
rect 14183 7993 14209 7999
rect 14183 7961 14209 7967
rect 14855 7993 14881 7999
rect 14855 7961 14881 7967
rect 6791 7937 6817 7943
rect 6791 7905 6817 7911
rect 9759 7937 9785 7943
rect 9759 7905 9785 7911
rect 11887 7937 11913 7943
rect 11887 7905 11913 7911
rect 14127 7937 14153 7943
rect 14127 7905 14153 7911
rect 14631 7937 14657 7943
rect 14631 7905 14657 7911
rect 672 7853 20328 7870
rect 672 7827 9919 7853
rect 9945 7827 9971 7853
rect 9997 7827 10023 7853
rect 10049 7827 20328 7853
rect 672 7810 20328 7827
rect 7239 7769 7265 7775
rect 7239 7737 7265 7743
rect 7295 7769 7321 7775
rect 7295 7737 7321 7743
rect 7743 7769 7769 7775
rect 7743 7737 7769 7743
rect 9591 7769 9617 7775
rect 9591 7737 9617 7743
rect 9759 7769 9785 7775
rect 9759 7737 9785 7743
rect 11215 7769 11241 7775
rect 11215 7737 11241 7743
rect 11439 7769 11465 7775
rect 11439 7737 11465 7743
rect 11719 7769 11745 7775
rect 11719 7737 11745 7743
rect 11775 7769 11801 7775
rect 11775 7737 11801 7743
rect 15135 7769 15161 7775
rect 15135 7737 15161 7743
rect 7519 7713 7545 7719
rect 7519 7681 7545 7687
rect 9031 7713 9057 7719
rect 9031 7681 9057 7687
rect 9143 7713 9169 7719
rect 9143 7681 9169 7687
rect 9479 7713 9505 7719
rect 9479 7681 9505 7687
rect 10655 7713 10681 7719
rect 13841 7687 13847 7713
rect 13873 7687 13879 7713
rect 10655 7681 10681 7687
rect 8807 7657 8833 7663
rect 6729 7631 6735 7657
rect 6761 7631 6767 7657
rect 7065 7631 7071 7657
rect 7097 7631 7103 7657
rect 7401 7631 7407 7657
rect 7433 7631 7439 7657
rect 8807 7625 8833 7631
rect 8919 7657 8945 7663
rect 8919 7625 8945 7631
rect 9703 7657 9729 7663
rect 9703 7625 9729 7631
rect 10823 7657 10849 7663
rect 10823 7625 10849 7631
rect 10935 7657 10961 7663
rect 10935 7625 10961 7631
rect 11327 7657 11353 7663
rect 11327 7625 11353 7631
rect 11831 7657 11857 7663
rect 11831 7625 11857 7631
rect 12055 7657 12081 7663
rect 13449 7631 13455 7657
rect 13481 7631 13487 7657
rect 12055 7625 12081 7631
rect 9647 7601 9673 7607
rect 11383 7601 11409 7607
rect 5665 7575 5671 7601
rect 5697 7575 5703 7601
rect 10705 7575 10711 7601
rect 10737 7575 10743 7601
rect 14905 7575 14911 7601
rect 14937 7575 14943 7601
rect 9647 7569 9673 7575
rect 11383 7569 11409 7575
rect 10543 7545 10569 7551
rect 10543 7513 10569 7519
rect 672 7461 20328 7478
rect 672 7435 2239 7461
rect 2265 7435 2291 7461
rect 2317 7435 2343 7461
rect 2369 7435 17599 7461
rect 17625 7435 17651 7461
rect 17677 7435 17703 7461
rect 17729 7435 20328 7461
rect 672 7418 20328 7435
rect 6847 7377 6873 7383
rect 6847 7345 6873 7351
rect 9535 7377 9561 7383
rect 9535 7345 9561 7351
rect 10767 7377 10793 7383
rect 10767 7345 10793 7351
rect 11327 7377 11353 7383
rect 11327 7345 11353 7351
rect 12049 7295 12055 7321
rect 12081 7295 12087 7321
rect 13113 7295 13119 7321
rect 13145 7295 13151 7321
rect 7183 7265 7209 7271
rect 7009 7239 7015 7265
rect 7041 7239 7047 7265
rect 7183 7233 7209 7239
rect 8583 7265 8609 7271
rect 11103 7265 11129 7271
rect 9697 7239 9703 7265
rect 9729 7239 9735 7265
rect 10929 7239 10935 7265
rect 10961 7239 10967 7265
rect 11489 7239 11495 7265
rect 11521 7239 11527 7265
rect 11657 7239 11663 7265
rect 11689 7239 11695 7265
rect 8583 7233 8609 7239
rect 11103 7233 11129 7239
rect 6903 7209 6929 7215
rect 6903 7177 6929 7183
rect 8751 7209 8777 7215
rect 8751 7177 8777 7183
rect 8639 7153 8665 7159
rect 8639 7121 8665 7127
rect 8919 7153 8945 7159
rect 8919 7121 8945 7127
rect 9591 7153 9617 7159
rect 9591 7121 9617 7127
rect 10823 7153 10849 7159
rect 10823 7121 10849 7127
rect 11383 7153 11409 7159
rect 11383 7121 11409 7127
rect 13343 7153 13369 7159
rect 13343 7121 13369 7127
rect 672 7069 20328 7086
rect 672 7043 9919 7069
rect 9945 7043 9971 7069
rect 9997 7043 10023 7069
rect 10049 7043 20328 7069
rect 672 7026 20328 7043
rect 8751 6985 8777 6991
rect 8751 6953 8777 6959
rect 8975 6985 9001 6991
rect 8975 6953 9001 6959
rect 13511 6985 13537 6991
rect 13511 6953 13537 6959
rect 9087 6929 9113 6935
rect 7345 6903 7351 6929
rect 7377 6903 7383 6929
rect 9641 6903 9647 6929
rect 9673 6903 9679 6929
rect 11265 6903 11271 6929
rect 11297 6903 11303 6929
rect 14065 6903 14071 6929
rect 14097 6903 14103 6929
rect 9087 6897 9113 6903
rect 12671 6873 12697 6879
rect 7009 6847 7015 6873
rect 7041 6847 7047 6873
rect 9249 6847 9255 6873
rect 9281 6847 9287 6873
rect 10929 6847 10935 6873
rect 10961 6847 10967 6873
rect 13673 6847 13679 6873
rect 13705 6847 13711 6873
rect 12671 6841 12697 6847
rect 8409 6791 8415 6817
rect 8441 6791 8447 6817
rect 10705 6791 10711 6817
rect 10737 6791 10743 6817
rect 12329 6791 12335 6817
rect 12361 6791 12367 6817
rect 15129 6791 15135 6817
rect 15161 6791 15167 6817
rect 8919 6761 8945 6767
rect 8919 6729 8945 6735
rect 672 6677 20328 6694
rect 672 6651 2239 6677
rect 2265 6651 2291 6677
rect 2317 6651 2343 6677
rect 2369 6651 17599 6677
rect 17625 6651 17651 6677
rect 17677 6651 17703 6677
rect 17729 6651 20328 6677
rect 672 6634 20328 6651
rect 10207 6537 10233 6543
rect 8913 6511 8919 6537
rect 8945 6511 8951 6537
rect 9977 6511 9983 6537
rect 10009 6511 10015 6537
rect 10207 6505 10233 6511
rect 8577 6455 8583 6481
rect 8609 6455 8615 6481
rect 672 6285 20328 6302
rect 672 6259 9919 6285
rect 9945 6259 9971 6285
rect 9997 6259 10023 6285
rect 10049 6259 20328 6285
rect 672 6242 20328 6259
rect 672 5893 20328 5910
rect 672 5867 2239 5893
rect 2265 5867 2291 5893
rect 2317 5867 2343 5893
rect 2369 5867 17599 5893
rect 17625 5867 17651 5893
rect 17677 5867 17703 5893
rect 17729 5867 20328 5893
rect 672 5850 20328 5867
rect 672 5501 20328 5518
rect 672 5475 9919 5501
rect 9945 5475 9971 5501
rect 9997 5475 10023 5501
rect 10049 5475 20328 5501
rect 672 5458 20328 5475
rect 672 5109 20328 5126
rect 672 5083 2239 5109
rect 2265 5083 2291 5109
rect 2317 5083 2343 5109
rect 2369 5083 17599 5109
rect 17625 5083 17651 5109
rect 17677 5083 17703 5109
rect 17729 5083 20328 5109
rect 672 5066 20328 5083
rect 672 4717 20328 4734
rect 672 4691 9919 4717
rect 9945 4691 9971 4717
rect 9997 4691 10023 4717
rect 10049 4691 20328 4717
rect 672 4674 20328 4691
rect 672 4325 20328 4342
rect 672 4299 2239 4325
rect 2265 4299 2291 4325
rect 2317 4299 2343 4325
rect 2369 4299 17599 4325
rect 17625 4299 17651 4325
rect 17677 4299 17703 4325
rect 17729 4299 20328 4325
rect 672 4282 20328 4299
rect 672 3933 20328 3950
rect 672 3907 9919 3933
rect 9945 3907 9971 3933
rect 9997 3907 10023 3933
rect 10049 3907 20328 3933
rect 672 3890 20328 3907
rect 672 3541 20328 3558
rect 672 3515 2239 3541
rect 2265 3515 2291 3541
rect 2317 3515 2343 3541
rect 2369 3515 17599 3541
rect 17625 3515 17651 3541
rect 17677 3515 17703 3541
rect 17729 3515 20328 3541
rect 672 3498 20328 3515
rect 672 3149 20328 3166
rect 672 3123 9919 3149
rect 9945 3123 9971 3149
rect 9997 3123 10023 3149
rect 10049 3123 20328 3149
rect 672 3106 20328 3123
rect 672 2757 20328 2774
rect 672 2731 2239 2757
rect 2265 2731 2291 2757
rect 2317 2731 2343 2757
rect 2369 2731 17599 2757
rect 17625 2731 17651 2757
rect 17677 2731 17703 2757
rect 17729 2731 20328 2757
rect 672 2714 20328 2731
rect 9367 2617 9393 2623
rect 9367 2585 9393 2591
rect 8857 2535 8863 2561
rect 8889 2535 8895 2561
rect 672 2365 20328 2382
rect 672 2339 9919 2365
rect 9945 2339 9971 2365
rect 9997 2339 10023 2365
rect 10049 2339 20328 2365
rect 672 2322 20328 2339
rect 9865 2143 9871 2169
rect 9897 2143 9903 2169
rect 12609 2143 12615 2169
rect 12641 2143 12647 2169
rect 10375 2057 10401 2063
rect 10375 2025 10401 2031
rect 13119 2057 13145 2063
rect 13119 2025 13145 2031
rect 672 1973 20328 1990
rect 672 1947 2239 1973
rect 2265 1947 2291 1973
rect 2317 1947 2343 1973
rect 2369 1947 17599 1973
rect 17625 1947 17651 1973
rect 17677 1947 17703 1973
rect 17729 1947 20328 1973
rect 672 1930 20328 1947
rect 9311 1833 9337 1839
rect 9311 1801 9337 1807
rect 12783 1833 12809 1839
rect 12783 1801 12809 1807
rect 8801 1751 8807 1777
rect 8833 1751 8839 1777
rect 10705 1751 10711 1777
rect 10737 1751 10743 1777
rect 12273 1751 12279 1777
rect 12305 1751 12311 1777
rect 11215 1665 11241 1671
rect 11215 1633 11241 1639
rect 672 1581 20328 1598
rect 672 1555 9919 1581
rect 9945 1555 9971 1581
rect 9997 1555 10023 1581
rect 10049 1555 20328 1581
rect 672 1538 20328 1555
<< via1 >>
rect 2239 19195 2265 19221
rect 2291 19195 2317 19221
rect 2343 19195 2369 19221
rect 17599 19195 17625 19221
rect 17651 19195 17677 19221
rect 17703 19195 17729 19221
rect 9311 19111 9337 19137
rect 11215 19111 11241 19137
rect 12783 19111 12809 19137
rect 14687 19111 14713 19137
rect 8919 18999 8945 19025
rect 10879 18999 10905 19025
rect 12279 18999 12305 19025
rect 14295 18999 14321 19025
rect 9919 18803 9945 18829
rect 9971 18803 9997 18829
rect 10023 18803 10049 18829
rect 10039 18719 10065 18745
rect 13399 18719 13425 18745
rect 9535 18607 9561 18633
rect 12951 18607 12977 18633
rect 2239 18411 2265 18437
rect 2291 18411 2317 18437
rect 2343 18411 2369 18437
rect 17599 18411 17625 18437
rect 17651 18411 17677 18437
rect 17703 18411 17729 18437
rect 8359 18327 8385 18353
rect 7855 18215 7881 18241
rect 9919 18019 9945 18045
rect 9971 18019 9997 18045
rect 10023 18019 10049 18045
rect 2239 17627 2265 17653
rect 2291 17627 2317 17653
rect 2343 17627 2369 17653
rect 17599 17627 17625 17653
rect 17651 17627 17677 17653
rect 17703 17627 17729 17653
rect 9919 17235 9945 17261
rect 9971 17235 9997 17261
rect 10023 17235 10049 17261
rect 2239 16843 2265 16869
rect 2291 16843 2317 16869
rect 2343 16843 2369 16869
rect 17599 16843 17625 16869
rect 17651 16843 17677 16869
rect 17703 16843 17729 16869
rect 9919 16451 9945 16477
rect 9971 16451 9997 16477
rect 10023 16451 10049 16477
rect 2239 16059 2265 16085
rect 2291 16059 2317 16085
rect 2343 16059 2369 16085
rect 17599 16059 17625 16085
rect 17651 16059 17677 16085
rect 17703 16059 17729 16085
rect 9919 15667 9945 15693
rect 9971 15667 9997 15693
rect 10023 15667 10049 15693
rect 2239 15275 2265 15301
rect 2291 15275 2317 15301
rect 2343 15275 2369 15301
rect 17599 15275 17625 15301
rect 17651 15275 17677 15301
rect 17703 15275 17729 15301
rect 9919 14883 9945 14909
rect 9971 14883 9997 14909
rect 10023 14883 10049 14909
rect 2239 14491 2265 14517
rect 2291 14491 2317 14517
rect 2343 14491 2369 14517
rect 17599 14491 17625 14517
rect 17651 14491 17677 14517
rect 17703 14491 17729 14517
rect 10935 14295 10961 14321
rect 10879 14183 10905 14209
rect 9919 14099 9945 14125
rect 9971 14099 9997 14125
rect 10023 14099 10049 14125
rect 12951 14015 12977 14041
rect 13119 14015 13145 14041
rect 10599 13959 10625 13985
rect 12671 13959 12697 13985
rect 6231 13903 6257 13929
rect 10263 13903 10289 13929
rect 11943 13903 11969 13929
rect 6567 13847 6593 13873
rect 7631 13847 7657 13873
rect 7911 13847 7937 13873
rect 11663 13847 11689 13873
rect 12615 13791 12641 13817
rect 2239 13707 2265 13733
rect 2291 13707 2317 13733
rect 2343 13707 2369 13733
rect 17599 13707 17625 13733
rect 17651 13707 17677 13733
rect 17703 13707 17729 13733
rect 7127 13623 7153 13649
rect 8919 13567 8945 13593
rect 10711 13567 10737 13593
rect 13175 13567 13201 13593
rect 20007 13567 20033 13593
rect 7463 13511 7489 13537
rect 9031 13511 9057 13537
rect 9199 13511 9225 13537
rect 10375 13511 10401 13537
rect 10823 13511 10849 13537
rect 11327 13511 11353 13537
rect 11439 13511 11465 13537
rect 11551 13511 11577 13537
rect 11775 13511 11801 13537
rect 13399 13511 13425 13537
rect 18831 13511 18857 13537
rect 7183 13455 7209 13481
rect 7855 13455 7881 13481
rect 9311 13455 9337 13481
rect 10207 13455 10233 13481
rect 10655 13455 10681 13481
rect 10935 13455 10961 13481
rect 11103 13455 11129 13481
rect 11215 13455 11241 13481
rect 12111 13455 12137 13481
rect 9367 13399 9393 13425
rect 9535 13399 9561 13425
rect 10319 13399 10345 13425
rect 11607 13399 11633 13425
rect 9919 13315 9945 13341
rect 9971 13315 9997 13341
rect 10023 13315 10049 13341
rect 8919 13231 8945 13257
rect 11831 13231 11857 13257
rect 14295 13231 14321 13257
rect 7911 13175 7937 13201
rect 8079 13175 8105 13201
rect 9983 13175 10009 13201
rect 11775 13175 11801 13201
rect 12111 13175 12137 13201
rect 2143 13119 2169 13145
rect 5615 13119 5641 13145
rect 7687 13119 7713 13145
rect 8023 13119 8049 13145
rect 8191 13119 8217 13145
rect 8415 13119 8441 13145
rect 8695 13119 8721 13145
rect 9031 13119 9057 13145
rect 9087 13119 9113 13145
rect 9199 13119 9225 13145
rect 9591 13119 9617 13145
rect 11271 13119 11297 13145
rect 11719 13119 11745 13145
rect 12223 13119 12249 13145
rect 12615 13119 12641 13145
rect 5951 13063 5977 13089
rect 7015 13063 7041 13089
rect 7239 13063 7265 13089
rect 9423 13063 9449 13089
rect 11047 13063 11073 13089
rect 13007 13063 13033 13089
rect 14071 13063 14097 13089
rect 967 13007 993 13033
rect 7743 13007 7769 13033
rect 8359 13007 8385 13033
rect 8751 13007 8777 13033
rect 2239 12923 2265 12949
rect 2291 12923 2317 12949
rect 2343 12923 2369 12949
rect 17599 12923 17625 12949
rect 17651 12923 17677 12949
rect 17703 12923 17729 12949
rect 10319 12839 10345 12865
rect 10655 12839 10681 12865
rect 7575 12783 7601 12809
rect 7799 12783 7825 12809
rect 9703 12783 9729 12809
rect 10823 12783 10849 12809
rect 12279 12783 12305 12809
rect 7463 12727 7489 12753
rect 7743 12727 7769 12753
rect 8247 12727 8273 12753
rect 11159 12727 11185 12753
rect 12055 12727 12081 12753
rect 12335 12727 12361 12753
rect 13175 12727 13201 12753
rect 6231 12671 6257 12697
rect 6399 12671 6425 12697
rect 7295 12671 7321 12697
rect 8639 12671 8665 12697
rect 10375 12671 10401 12697
rect 10991 12671 11017 12697
rect 12167 12671 12193 12697
rect 13287 12671 13313 12697
rect 13343 12671 13369 12697
rect 9927 12615 9953 12641
rect 10319 12615 10345 12641
rect 10767 12615 10793 12641
rect 9919 12531 9945 12557
rect 9971 12531 9997 12557
rect 10023 12531 10049 12557
rect 7575 12447 7601 12473
rect 7631 12447 7657 12473
rect 9087 12447 9113 12473
rect 9143 12447 9169 12473
rect 10711 12447 10737 12473
rect 13679 12447 13705 12473
rect 7519 12335 7545 12361
rect 7855 12335 7881 12361
rect 9031 12335 9057 12361
rect 9367 12335 9393 12361
rect 10823 12335 10849 12361
rect 13847 12335 13873 12361
rect 18831 12335 18857 12361
rect 14239 12279 14265 12305
rect 15303 12279 15329 12305
rect 20007 12223 20033 12249
rect 2239 12139 2265 12165
rect 2291 12139 2317 12165
rect 2343 12139 2369 12165
rect 17599 12139 17625 12165
rect 17651 12139 17677 12165
rect 17703 12139 17729 12165
rect 7127 12055 7153 12081
rect 967 11999 993 12025
rect 6959 11999 6985 12025
rect 11831 11999 11857 12025
rect 13455 11999 13481 12025
rect 20007 11999 20033 12025
rect 2143 11943 2169 11969
rect 8695 11943 8721 11969
rect 10767 11943 10793 11969
rect 11943 11943 11969 11969
rect 13959 11943 13985 11969
rect 18831 11943 18857 11969
rect 7015 11887 7041 11913
rect 8583 11887 8609 11913
rect 10879 11887 10905 11913
rect 11159 11887 11185 11913
rect 12111 11887 12137 11913
rect 12279 11887 12305 11913
rect 7631 11831 7657 11857
rect 11215 11831 11241 11857
rect 12447 11831 12473 11857
rect 13847 11831 13873 11857
rect 13903 11831 13929 11857
rect 14071 11831 14097 11857
rect 9919 11747 9945 11773
rect 9971 11747 9997 11773
rect 10023 11747 10049 11773
rect 9311 11663 9337 11689
rect 9759 11663 9785 11689
rect 11831 11663 11857 11689
rect 13287 11663 13313 11689
rect 9647 11607 9673 11633
rect 9871 11607 9897 11633
rect 10543 11607 10569 11633
rect 11047 11607 11073 11633
rect 11943 11607 11969 11633
rect 11999 11607 12025 11633
rect 13399 11607 13425 11633
rect 13455 11607 13481 11633
rect 15415 11607 15441 11633
rect 2143 11551 2169 11577
rect 7519 11557 7545 11583
rect 7687 11551 7713 11577
rect 7799 11551 7825 11577
rect 7967 11551 7993 11577
rect 9479 11551 9505 11577
rect 10319 11551 10345 11577
rect 10711 11551 10737 11577
rect 10991 11551 11017 11577
rect 11439 11551 11465 11577
rect 12895 11551 12921 11577
rect 13119 11551 13145 11577
rect 13623 11551 13649 11577
rect 15247 11551 15273 11577
rect 18831 11551 18857 11577
rect 6063 11495 6089 11521
rect 7127 11495 7153 11521
rect 7743 11495 7769 11521
rect 10095 11495 10121 11521
rect 11215 11495 11241 11521
rect 11663 11495 11689 11521
rect 14015 11495 14041 11521
rect 15079 11495 15105 11521
rect 967 11439 993 11465
rect 9591 11439 9617 11465
rect 20007 11439 20033 11465
rect 2239 11355 2265 11381
rect 2291 11355 2317 11381
rect 2343 11355 2369 11381
rect 17599 11355 17625 11381
rect 17651 11355 17677 11381
rect 17703 11355 17729 11381
rect 7631 11271 7657 11297
rect 14183 11271 14209 11297
rect 7519 11215 7545 11241
rect 9199 11215 9225 11241
rect 10375 11215 10401 11241
rect 11719 11215 11745 11241
rect 12447 11215 12473 11241
rect 13511 11215 13537 11241
rect 13903 11215 13929 11241
rect 6847 11159 6873 11185
rect 6959 11159 6985 11185
rect 8359 11159 8385 11185
rect 8751 11159 8777 11185
rect 9087 11159 9113 11185
rect 9479 11159 9505 11185
rect 10095 11159 10121 11185
rect 10935 11159 10961 11185
rect 11103 11159 11129 11185
rect 11775 11159 11801 11185
rect 12111 11159 12137 11185
rect 13791 11159 13817 11185
rect 14015 11159 14041 11185
rect 7519 11103 7545 11129
rect 8583 11103 8609 11129
rect 8919 11103 8945 11129
rect 13679 11103 13705 11129
rect 14127 11103 14153 11129
rect 14183 11103 14209 11129
rect 6903 11047 6929 11073
rect 7071 11047 7097 11073
rect 8247 11047 8273 11073
rect 10655 11047 10681 11073
rect 11383 11047 11409 11073
rect 11551 11047 11577 11073
rect 11663 11047 11689 11073
rect 9919 10963 9945 10989
rect 9971 10963 9997 10989
rect 10023 10963 10049 10989
rect 8751 10879 8777 10905
rect 8807 10879 8833 10905
rect 9703 10879 9729 10905
rect 10151 10879 10177 10905
rect 10599 10879 10625 10905
rect 13063 10879 13089 10905
rect 13791 10879 13817 10905
rect 14015 10879 14041 10905
rect 6623 10823 6649 10849
rect 8415 10823 8441 10849
rect 9367 10823 9393 10849
rect 9647 10823 9673 10849
rect 10655 10823 10681 10849
rect 13287 10823 13313 10849
rect 13511 10823 13537 10849
rect 13567 10823 13593 10849
rect 7015 10767 7041 10793
rect 8303 10767 8329 10793
rect 8919 10767 8945 10793
rect 9087 10767 9113 10793
rect 9759 10767 9785 10793
rect 10319 10767 10345 10793
rect 10599 10767 10625 10793
rect 12055 10767 12081 10793
rect 12335 10767 12361 10793
rect 13231 10767 13257 10793
rect 5559 10711 5585 10737
rect 7239 10711 7265 10737
rect 12783 10711 12809 10737
rect 13287 10655 13313 10681
rect 2239 10571 2265 10597
rect 2291 10571 2317 10597
rect 2343 10571 2369 10597
rect 17599 10571 17625 10597
rect 17651 10571 17677 10597
rect 17703 10571 17729 10597
rect 11439 10487 11465 10513
rect 7071 10431 7097 10457
rect 7351 10431 7377 10457
rect 7855 10431 7881 10457
rect 11495 10431 11521 10457
rect 13735 10431 13761 10457
rect 10039 10375 10065 10401
rect 11215 10375 11241 10401
rect 11271 10375 11297 10401
rect 11663 10375 11689 10401
rect 10823 10319 10849 10345
rect 11103 10319 11129 10345
rect 6847 10263 6873 10289
rect 9919 10179 9945 10205
rect 9971 10179 9997 10205
rect 10023 10179 10049 10205
rect 6007 10039 6033 10065
rect 7407 10039 7433 10065
rect 7743 10039 7769 10065
rect 8191 10039 8217 10065
rect 11047 10039 11073 10065
rect 13399 10039 13425 10065
rect 13791 10039 13817 10065
rect 5615 9983 5641 10009
rect 7239 9983 7265 10009
rect 7575 9983 7601 10009
rect 8023 9983 8049 10009
rect 9143 9983 9169 10009
rect 9255 9983 9281 10009
rect 9703 9983 9729 10009
rect 12727 9983 12753 10009
rect 13119 9983 13145 10009
rect 13847 9983 13873 10009
rect 14015 9983 14041 10009
rect 18831 9983 18857 10009
rect 7071 9927 7097 9953
rect 7911 9927 7937 9953
rect 8751 9927 8777 9953
rect 9087 9927 9113 9953
rect 13063 9927 13089 9953
rect 14407 9927 14433 9953
rect 15471 9927 15497 9953
rect 9255 9871 9281 9897
rect 13791 9871 13817 9897
rect 20007 9871 20033 9897
rect 2239 9787 2265 9813
rect 2291 9787 2317 9813
rect 2343 9787 2369 9813
rect 17599 9787 17625 9813
rect 17651 9787 17677 9813
rect 17703 9787 17729 9813
rect 8639 9703 8665 9729
rect 10711 9703 10737 9729
rect 11607 9703 11633 9729
rect 13287 9703 13313 9729
rect 13679 9703 13705 9729
rect 15079 9703 15105 9729
rect 6735 9647 6761 9673
rect 6903 9647 6929 9673
rect 10991 9647 11017 9673
rect 11887 9647 11913 9673
rect 14127 9647 14153 9673
rect 14799 9647 14825 9673
rect 20007 9647 20033 9673
rect 7071 9591 7097 9617
rect 7743 9591 7769 9617
rect 7967 9591 7993 9617
rect 8415 9591 8441 9617
rect 8807 9591 8833 9617
rect 8975 9591 9001 9617
rect 10039 9591 10065 9617
rect 10375 9591 10401 9617
rect 11159 9591 11185 9617
rect 11383 9591 11409 9617
rect 11831 9591 11857 9617
rect 12223 9591 12249 9617
rect 12951 9591 12977 9617
rect 13175 9591 13201 9617
rect 13455 9591 13481 9617
rect 13623 9591 13649 9617
rect 14575 9591 14601 9617
rect 14911 9591 14937 9617
rect 18831 9591 18857 9617
rect 8527 9535 8553 9561
rect 10655 9535 10681 9561
rect 13959 9535 13985 9561
rect 14071 9535 14097 9561
rect 14183 9535 14209 9561
rect 14687 9535 14713 9561
rect 15023 9535 15049 9561
rect 8695 9479 8721 9505
rect 9143 9479 9169 9505
rect 9311 9479 9337 9505
rect 9479 9479 9505 9505
rect 9647 9479 9673 9505
rect 9871 9479 9897 9505
rect 10207 9479 10233 9505
rect 12111 9479 12137 9505
rect 12839 9479 12865 9505
rect 13679 9479 13705 9505
rect 14239 9479 14265 9505
rect 15079 9479 15105 9505
rect 9919 9395 9945 9421
rect 9971 9395 9997 9421
rect 10023 9395 10049 9421
rect 8023 9311 8049 9337
rect 8639 9311 8665 9337
rect 10431 9311 10457 9337
rect 11831 9311 11857 9337
rect 8191 9255 8217 9281
rect 10879 9255 10905 9281
rect 14239 9255 14265 9281
rect 5559 9199 5585 9225
rect 7183 9199 7209 9225
rect 8863 9199 8889 9225
rect 8975 9199 9001 9225
rect 9759 9199 9785 9225
rect 9871 9199 9897 9225
rect 10991 9199 11017 9225
rect 11439 9199 11465 9225
rect 11495 9199 11521 9225
rect 11719 9199 11745 9225
rect 11943 9199 11969 9225
rect 13847 9199 13873 9225
rect 5895 9143 5921 9169
rect 6959 9143 6985 9169
rect 9031 9143 9057 9169
rect 9647 9143 9673 9169
rect 10655 9143 10681 9169
rect 11607 9143 11633 9169
rect 13679 9143 13705 9169
rect 15303 9143 15329 9169
rect 10095 9087 10121 9113
rect 2239 9003 2265 9029
rect 2291 9003 2317 9029
rect 2343 9003 2369 9029
rect 17599 9003 17625 9029
rect 17651 9003 17677 9029
rect 17703 9003 17729 9029
rect 9087 8919 9113 8945
rect 9927 8919 9953 8945
rect 11159 8919 11185 8945
rect 7183 8863 7209 8889
rect 11439 8863 11465 8889
rect 12503 8863 12529 8889
rect 9031 8807 9057 8833
rect 9311 8807 9337 8833
rect 9871 8807 9897 8833
rect 12895 8807 12921 8833
rect 9199 8751 9225 8777
rect 9927 8751 9953 8777
rect 11103 8751 11129 8777
rect 11159 8751 11185 8777
rect 8919 8695 8945 8721
rect 13119 8695 13145 8721
rect 9919 8611 9945 8637
rect 9971 8611 9997 8637
rect 10023 8611 10049 8637
rect 7519 8527 7545 8553
rect 8191 8527 8217 8553
rect 8303 8527 8329 8553
rect 10487 8527 10513 8553
rect 9535 8471 9561 8497
rect 9591 8471 9617 8497
rect 10319 8471 10345 8497
rect 11271 8471 11297 8497
rect 14183 8471 14209 8497
rect 2143 8415 2169 8441
rect 7071 8415 7097 8441
rect 7239 8415 7265 8441
rect 7407 8415 7433 8441
rect 8415 8415 8441 8441
rect 8975 8415 9001 8441
rect 9143 8415 9169 8441
rect 9423 8415 9449 8441
rect 10711 8415 10737 8441
rect 11047 8415 11073 8441
rect 11327 8415 11353 8441
rect 13847 8415 13873 8441
rect 14071 8415 14097 8441
rect 18943 8415 18969 8441
rect 5615 8359 5641 8385
rect 6679 8359 6705 8385
rect 7463 8359 7489 8385
rect 8359 8359 8385 8385
rect 9199 8359 9225 8385
rect 11439 8359 11465 8385
rect 13959 8359 13985 8385
rect 19951 8359 19977 8385
rect 967 8303 993 8329
rect 9255 8303 9281 8329
rect 2239 8219 2265 8245
rect 2291 8219 2317 8245
rect 2343 8219 2369 8245
rect 17599 8219 17625 8245
rect 17651 8219 17677 8245
rect 17703 8219 17729 8245
rect 1023 8079 1049 8105
rect 6959 8079 6985 8105
rect 7911 8079 7937 8105
rect 8975 8079 9001 8105
rect 9423 8079 9449 8105
rect 20007 8079 20033 8105
rect 2143 8023 2169 8049
rect 6903 8023 6929 8049
rect 7015 8023 7041 8049
rect 7519 8023 7545 8049
rect 9143 8023 9169 8049
rect 9311 8023 9337 8049
rect 9367 8023 9393 8049
rect 9479 8023 9505 8049
rect 11887 8023 11913 8049
rect 11999 8023 12025 8049
rect 13679 8023 13705 8049
rect 13847 8023 13873 8049
rect 13959 8023 13985 8049
rect 14071 8023 14097 8049
rect 14519 8023 14545 8049
rect 14687 8023 14713 8049
rect 14911 8023 14937 8049
rect 18831 8023 18857 8049
rect 11775 7967 11801 7993
rect 14183 7967 14209 7993
rect 14855 7967 14881 7993
rect 6791 7911 6817 7937
rect 9759 7911 9785 7937
rect 11887 7911 11913 7937
rect 14127 7911 14153 7937
rect 14631 7911 14657 7937
rect 9919 7827 9945 7853
rect 9971 7827 9997 7853
rect 10023 7827 10049 7853
rect 7239 7743 7265 7769
rect 7295 7743 7321 7769
rect 7743 7743 7769 7769
rect 9591 7743 9617 7769
rect 9759 7743 9785 7769
rect 11215 7743 11241 7769
rect 11439 7743 11465 7769
rect 11719 7743 11745 7769
rect 11775 7743 11801 7769
rect 15135 7743 15161 7769
rect 7519 7687 7545 7713
rect 9031 7687 9057 7713
rect 9143 7687 9169 7713
rect 9479 7687 9505 7713
rect 10655 7687 10681 7713
rect 13847 7687 13873 7713
rect 6735 7631 6761 7657
rect 7071 7631 7097 7657
rect 7407 7631 7433 7657
rect 8807 7631 8833 7657
rect 8919 7631 8945 7657
rect 9703 7631 9729 7657
rect 10823 7631 10849 7657
rect 10935 7631 10961 7657
rect 11327 7631 11353 7657
rect 11831 7631 11857 7657
rect 12055 7631 12081 7657
rect 13455 7631 13481 7657
rect 5671 7575 5697 7601
rect 9647 7575 9673 7601
rect 10711 7575 10737 7601
rect 11383 7575 11409 7601
rect 14911 7575 14937 7601
rect 10543 7519 10569 7545
rect 2239 7435 2265 7461
rect 2291 7435 2317 7461
rect 2343 7435 2369 7461
rect 17599 7435 17625 7461
rect 17651 7435 17677 7461
rect 17703 7435 17729 7461
rect 6847 7351 6873 7377
rect 9535 7351 9561 7377
rect 10767 7351 10793 7377
rect 11327 7351 11353 7377
rect 12055 7295 12081 7321
rect 13119 7295 13145 7321
rect 7015 7239 7041 7265
rect 7183 7239 7209 7265
rect 8583 7239 8609 7265
rect 9703 7239 9729 7265
rect 10935 7239 10961 7265
rect 11103 7239 11129 7265
rect 11495 7239 11521 7265
rect 11663 7239 11689 7265
rect 6903 7183 6929 7209
rect 8751 7183 8777 7209
rect 8639 7127 8665 7153
rect 8919 7127 8945 7153
rect 9591 7127 9617 7153
rect 10823 7127 10849 7153
rect 11383 7127 11409 7153
rect 13343 7127 13369 7153
rect 9919 7043 9945 7069
rect 9971 7043 9997 7069
rect 10023 7043 10049 7069
rect 8751 6959 8777 6985
rect 8975 6959 9001 6985
rect 13511 6959 13537 6985
rect 7351 6903 7377 6929
rect 9087 6903 9113 6929
rect 9647 6903 9673 6929
rect 11271 6903 11297 6929
rect 14071 6903 14097 6929
rect 7015 6847 7041 6873
rect 9255 6847 9281 6873
rect 10935 6847 10961 6873
rect 12671 6847 12697 6873
rect 13679 6847 13705 6873
rect 8415 6791 8441 6817
rect 10711 6791 10737 6817
rect 12335 6791 12361 6817
rect 15135 6791 15161 6817
rect 8919 6735 8945 6761
rect 2239 6651 2265 6677
rect 2291 6651 2317 6677
rect 2343 6651 2369 6677
rect 17599 6651 17625 6677
rect 17651 6651 17677 6677
rect 17703 6651 17729 6677
rect 8919 6511 8945 6537
rect 9983 6511 10009 6537
rect 10207 6511 10233 6537
rect 8583 6455 8609 6481
rect 9919 6259 9945 6285
rect 9971 6259 9997 6285
rect 10023 6259 10049 6285
rect 2239 5867 2265 5893
rect 2291 5867 2317 5893
rect 2343 5867 2369 5893
rect 17599 5867 17625 5893
rect 17651 5867 17677 5893
rect 17703 5867 17729 5893
rect 9919 5475 9945 5501
rect 9971 5475 9997 5501
rect 10023 5475 10049 5501
rect 2239 5083 2265 5109
rect 2291 5083 2317 5109
rect 2343 5083 2369 5109
rect 17599 5083 17625 5109
rect 17651 5083 17677 5109
rect 17703 5083 17729 5109
rect 9919 4691 9945 4717
rect 9971 4691 9997 4717
rect 10023 4691 10049 4717
rect 2239 4299 2265 4325
rect 2291 4299 2317 4325
rect 2343 4299 2369 4325
rect 17599 4299 17625 4325
rect 17651 4299 17677 4325
rect 17703 4299 17729 4325
rect 9919 3907 9945 3933
rect 9971 3907 9997 3933
rect 10023 3907 10049 3933
rect 2239 3515 2265 3541
rect 2291 3515 2317 3541
rect 2343 3515 2369 3541
rect 17599 3515 17625 3541
rect 17651 3515 17677 3541
rect 17703 3515 17729 3541
rect 9919 3123 9945 3149
rect 9971 3123 9997 3149
rect 10023 3123 10049 3149
rect 2239 2731 2265 2757
rect 2291 2731 2317 2757
rect 2343 2731 2369 2757
rect 17599 2731 17625 2757
rect 17651 2731 17677 2757
rect 17703 2731 17729 2757
rect 9367 2591 9393 2617
rect 8863 2535 8889 2561
rect 9919 2339 9945 2365
rect 9971 2339 9997 2365
rect 10023 2339 10049 2365
rect 9871 2143 9897 2169
rect 12615 2143 12641 2169
rect 10375 2031 10401 2057
rect 13119 2031 13145 2057
rect 2239 1947 2265 1973
rect 2291 1947 2317 1973
rect 2343 1947 2369 1973
rect 17599 1947 17625 1973
rect 17651 1947 17677 1973
rect 17703 1947 17729 1973
rect 9311 1807 9337 1833
rect 12783 1807 12809 1833
rect 8807 1751 8833 1777
rect 10711 1751 10737 1777
rect 12279 1751 12305 1777
rect 11215 1639 11241 1665
rect 9919 1555 9945 1581
rect 9971 1555 9997 1581
rect 10023 1555 10049 1581
<< metal2 >>
rect 7728 20600 7784 21000
rect 8736 20600 8792 21000
rect 9408 20600 9464 21000
rect 11088 20600 11144 21000
rect 11424 20600 11480 21000
rect 12768 20600 12824 21000
rect 13104 20600 13160 21000
rect 2238 19222 2370 19227
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2238 19189 2370 19194
rect 2238 18438 2370 18443
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2238 18405 2370 18410
rect 7742 18354 7770 20600
rect 8750 19138 8778 20600
rect 8750 19105 8778 19110
rect 9310 19138 9338 19143
rect 9310 19091 9338 19110
rect 8918 19025 8946 19031
rect 8918 18999 8919 19025
rect 8945 18999 8946 19025
rect 7742 18321 7770 18326
rect 8358 18354 8386 18359
rect 8358 18307 8386 18326
rect 7854 18241 7882 18247
rect 7854 18215 7855 18241
rect 7881 18215 7882 18241
rect 2238 17654 2370 17659
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2238 17621 2370 17626
rect 2238 16870 2370 16875
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2238 16837 2370 16842
rect 2238 16086 2370 16091
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2238 16053 2370 16058
rect 7854 15974 7882 18215
rect 7630 15946 7882 15974
rect 2238 15302 2370 15307
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2238 15269 2370 15274
rect 2238 14518 2370 14523
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2238 14485 2370 14490
rect 6230 13929 6258 13935
rect 6230 13903 6231 13929
rect 6257 13903 6258 13929
rect 2086 13818 2114 13823
rect 966 13033 994 13039
rect 966 13007 967 13033
rect 993 13007 994 13033
rect 966 12810 994 13007
rect 966 12777 994 12782
rect 966 12025 994 12031
rect 966 11999 967 12025
rect 993 11999 994 12025
rect 966 11802 994 11999
rect 966 11769 994 11774
rect 966 11466 994 11471
rect 966 11419 994 11438
rect 2086 9954 2114 13790
rect 2238 13734 2370 13739
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2238 13701 2370 13706
rect 6230 13538 6258 13903
rect 6566 13874 6594 13879
rect 6566 13827 6594 13846
rect 7126 13874 7154 13879
rect 7126 13649 7154 13846
rect 7630 13874 7658 15946
rect 7630 13873 7714 13874
rect 7630 13847 7631 13873
rect 7657 13847 7714 13873
rect 7630 13846 7714 13847
rect 7630 13841 7658 13846
rect 7126 13623 7127 13649
rect 7153 13623 7154 13649
rect 7126 13617 7154 13623
rect 6230 13505 6258 13510
rect 7462 13538 7490 13543
rect 7182 13481 7210 13487
rect 7182 13455 7183 13481
rect 7209 13455 7210 13481
rect 5614 13426 5642 13431
rect 2142 13145 2170 13151
rect 2142 13119 2143 13145
rect 2169 13119 2170 13145
rect 2142 13090 2170 13119
rect 5614 13145 5642 13398
rect 7182 13202 7210 13455
rect 7182 13169 7210 13174
rect 5614 13119 5615 13145
rect 5641 13119 5642 13145
rect 5614 13113 5642 13119
rect 2142 13057 2170 13062
rect 5950 13090 5978 13095
rect 7014 13090 7042 13095
rect 5950 13089 6258 13090
rect 5950 13063 5951 13089
rect 5977 13063 6258 13089
rect 5950 13062 6258 13063
rect 5950 13057 5978 13062
rect 2238 12950 2370 12955
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2238 12917 2370 12922
rect 6230 12697 6258 13062
rect 7014 13043 7042 13062
rect 7238 13090 7266 13095
rect 7462 13090 7490 13510
rect 7686 13145 7714 13846
rect 7910 13873 7938 13879
rect 7910 13847 7911 13873
rect 7937 13847 7938 13873
rect 7910 13538 7938 13847
rect 7910 13505 7938 13510
rect 8190 13594 8218 13599
rect 8918 13594 8946 18999
rect 9422 18746 9450 20600
rect 11102 19138 11130 20600
rect 11214 19138 11242 19143
rect 11102 19137 11242 19138
rect 11102 19111 11215 19137
rect 11241 19111 11242 19137
rect 11102 19110 11242 19111
rect 11214 19105 11242 19110
rect 11438 19138 11466 20600
rect 12782 19306 12810 20600
rect 12782 19273 12810 19278
rect 11438 19105 11466 19110
rect 12782 19138 12810 19143
rect 12782 19091 12810 19110
rect 13118 19138 13146 20600
rect 13118 19105 13146 19110
rect 13398 19306 13426 19311
rect 10878 19025 10906 19031
rect 10878 18999 10879 19025
rect 10905 18999 10906 19025
rect 9918 18830 10050 18835
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 9918 18797 10050 18802
rect 9422 18713 9450 18718
rect 10038 18746 10066 18751
rect 10038 18699 10066 18718
rect 9534 18633 9562 18639
rect 9534 18607 9535 18633
rect 9561 18607 9562 18633
rect 9534 15974 9562 18607
rect 9918 18046 10050 18051
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 9918 18013 10050 18018
rect 9918 17262 10050 17267
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 9918 17229 10050 17234
rect 9918 16478 10050 16483
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 9918 16445 10050 16450
rect 9310 15946 9562 15974
rect 7854 13481 7882 13487
rect 7854 13455 7855 13481
rect 7881 13455 7882 13481
rect 7854 13314 7882 13455
rect 7854 13286 8162 13314
rect 7686 13119 7687 13145
rect 7713 13119 7714 13145
rect 7686 13113 7714 13119
rect 7910 13201 7938 13207
rect 7910 13175 7911 13201
rect 7937 13175 7938 13201
rect 7238 13089 7490 13090
rect 7238 13063 7239 13089
rect 7265 13063 7490 13089
rect 7238 13062 7490 13063
rect 7798 13090 7826 13095
rect 6230 12671 6231 12697
rect 6257 12671 6258 12697
rect 6230 12665 6258 12671
rect 6398 12698 6426 12703
rect 6398 12651 6426 12670
rect 7238 12642 7266 13062
rect 7574 13034 7602 13039
rect 7518 12978 7546 12983
rect 7462 12753 7490 12759
rect 7462 12727 7463 12753
rect 7489 12727 7490 12753
rect 7294 12698 7322 12703
rect 7294 12651 7322 12670
rect 7238 12609 7266 12614
rect 7462 12474 7490 12727
rect 7462 12441 7490 12446
rect 7518 12362 7546 12950
rect 7574 12809 7602 13006
rect 7742 13033 7770 13039
rect 7742 13007 7743 13033
rect 7769 13007 7770 13033
rect 7742 12978 7770 13007
rect 7742 12945 7770 12950
rect 7574 12783 7575 12809
rect 7601 12783 7602 12809
rect 7574 12777 7602 12783
rect 7798 12809 7826 13062
rect 7910 13090 7938 13175
rect 8078 13202 8106 13207
rect 8078 13155 8106 13174
rect 8022 13146 8050 13151
rect 7910 13057 7938 13062
rect 7966 13145 8050 13146
rect 7966 13119 8023 13145
rect 8049 13119 8050 13145
rect 7966 13118 8050 13119
rect 7798 12783 7799 12809
rect 7825 12783 7826 12809
rect 7798 12777 7826 12783
rect 7742 12754 7770 12759
rect 7630 12753 7770 12754
rect 7630 12727 7743 12753
rect 7769 12727 7770 12753
rect 7630 12726 7770 12727
rect 7574 12474 7602 12479
rect 7574 12427 7602 12446
rect 7630 12473 7658 12726
rect 7742 12721 7770 12726
rect 7630 12447 7631 12473
rect 7657 12447 7658 12473
rect 7630 12441 7658 12447
rect 7686 12642 7714 12647
rect 7126 12361 7546 12362
rect 7126 12335 7519 12361
rect 7545 12335 7546 12361
rect 7126 12334 7546 12335
rect 2238 12166 2370 12171
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2238 12133 2370 12138
rect 7126 12081 7154 12334
rect 7518 12329 7546 12334
rect 7126 12055 7127 12081
rect 7153 12055 7154 12081
rect 7126 12049 7154 12055
rect 6958 12026 6986 12031
rect 6846 12025 6986 12026
rect 6846 11999 6959 12025
rect 6985 11999 6986 12025
rect 6846 11998 6986 11999
rect 2142 11970 2170 11975
rect 2142 11923 2170 11942
rect 5558 11970 5586 11975
rect 2142 11578 2170 11583
rect 2142 11531 2170 11550
rect 2238 11382 2370 11387
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2238 11349 2370 11354
rect 5558 10737 5586 11942
rect 6062 11578 6090 11583
rect 6062 11521 6090 11550
rect 6062 11495 6063 11521
rect 6089 11495 6090 11521
rect 6062 11489 6090 11495
rect 6846 11185 6874 11998
rect 6958 11993 6986 11998
rect 7014 11970 7042 11975
rect 7014 11913 7042 11942
rect 7014 11887 7015 11913
rect 7041 11887 7042 11913
rect 7014 11881 7042 11887
rect 7630 11858 7658 11863
rect 7686 11858 7714 12614
rect 7518 11857 7714 11858
rect 7518 11831 7631 11857
rect 7657 11831 7714 11857
rect 7518 11830 7714 11831
rect 7854 12361 7882 12367
rect 7854 12335 7855 12361
rect 7881 12335 7882 12361
rect 7518 11583 7546 11830
rect 7630 11825 7658 11830
rect 7518 11557 7519 11583
rect 7545 11578 7546 11583
rect 7545 11557 7602 11578
rect 7518 11550 7602 11557
rect 7126 11522 7154 11527
rect 7126 11521 7546 11522
rect 7126 11495 7127 11521
rect 7153 11495 7546 11521
rect 7126 11494 7546 11495
rect 7126 11489 7154 11494
rect 6846 11159 6847 11185
rect 6873 11159 6874 11185
rect 6846 11153 6874 11159
rect 6958 11354 6986 11359
rect 6958 11185 6986 11326
rect 7518 11241 7546 11494
rect 7518 11215 7519 11241
rect 7545 11215 7546 11241
rect 7518 11209 7546 11215
rect 6958 11159 6959 11185
rect 6985 11159 6986 11185
rect 6958 11153 6986 11159
rect 7518 11130 7546 11135
rect 7518 11083 7546 11102
rect 6902 11073 6930 11079
rect 6902 11047 6903 11073
rect 6929 11047 6930 11073
rect 6902 10962 6930 11047
rect 7070 11074 7098 11079
rect 7070 11027 7098 11046
rect 7574 11018 7602 11550
rect 7686 11577 7714 11583
rect 7686 11551 7687 11577
rect 7713 11551 7714 11577
rect 7686 11466 7714 11551
rect 7798 11578 7826 11583
rect 7798 11531 7826 11550
rect 7686 11433 7714 11438
rect 7742 11521 7770 11527
rect 7742 11495 7743 11521
rect 7769 11495 7770 11521
rect 7742 11354 7770 11495
rect 7630 11326 7770 11354
rect 7630 11297 7658 11326
rect 7630 11271 7631 11297
rect 7657 11271 7658 11297
rect 7630 11265 7658 11271
rect 7854 11242 7882 12335
rect 7854 11209 7882 11214
rect 7966 11577 7994 13118
rect 8022 13113 8050 13118
rect 8134 13034 8162 13286
rect 8190 13145 8218 13566
rect 8694 13593 8946 13594
rect 8694 13567 8919 13593
rect 8945 13567 8946 13593
rect 8694 13566 8946 13567
rect 8190 13119 8191 13145
rect 8217 13119 8218 13145
rect 8190 13113 8218 13119
rect 8414 13146 8442 13151
rect 8414 13099 8442 13118
rect 8694 13145 8722 13566
rect 8918 13561 8946 13566
rect 9198 13594 9226 13599
rect 9030 13538 9058 13543
rect 8974 13537 9058 13538
rect 8974 13511 9031 13537
rect 9057 13511 9058 13537
rect 8974 13510 9058 13511
rect 8694 13119 8695 13145
rect 8721 13119 8722 13145
rect 8694 13113 8722 13119
rect 8918 13258 8946 13263
rect 8974 13258 9002 13510
rect 9030 13505 9058 13510
rect 9198 13537 9226 13566
rect 9198 13511 9199 13537
rect 9225 13511 9226 13537
rect 9198 13505 9226 13511
rect 9310 13538 9338 15946
rect 9918 15694 10050 15699
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 9918 15661 10050 15666
rect 9918 14910 10050 14915
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 9918 14877 10050 14882
rect 10878 14434 10906 18999
rect 12278 19025 12306 19031
rect 12278 18999 12279 19025
rect 12305 18999 12306 19025
rect 10878 14406 11018 14434
rect 10934 14321 10962 14327
rect 10934 14295 10935 14321
rect 10961 14295 10962 14321
rect 10934 14266 10962 14295
rect 10934 14233 10962 14238
rect 10878 14209 10906 14215
rect 10878 14183 10879 14209
rect 10905 14183 10906 14209
rect 9918 14126 10050 14131
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 9918 14093 10050 14098
rect 10878 14042 10906 14183
rect 10598 14014 10906 14042
rect 10598 13985 10626 14014
rect 10990 13986 11018 14406
rect 11830 14266 11858 14271
rect 10598 13959 10599 13985
rect 10625 13959 10626 13985
rect 10598 13953 10626 13959
rect 10822 13958 11074 13986
rect 10262 13930 10290 13935
rect 10262 13883 10290 13902
rect 10710 13594 10738 13599
rect 10374 13593 10738 13594
rect 10374 13567 10711 13593
rect 10737 13567 10738 13593
rect 10374 13566 10738 13567
rect 9310 13510 9730 13538
rect 9310 13481 9338 13510
rect 9310 13455 9311 13481
rect 9337 13455 9338 13481
rect 9310 13449 9338 13455
rect 8918 13257 9002 13258
rect 8918 13231 8919 13257
rect 8945 13231 9002 13257
rect 8918 13230 9002 13231
rect 9366 13425 9394 13431
rect 9366 13399 9367 13425
rect 9393 13399 9394 13425
rect 8582 13090 8610 13095
rect 8358 13034 8386 13039
rect 8134 13033 8386 13034
rect 8134 13007 8359 13033
rect 8385 13007 8386 13033
rect 8134 13006 8386 13007
rect 8358 13001 8386 13006
rect 8246 12753 8274 12759
rect 8246 12727 8247 12753
rect 8273 12727 8274 12753
rect 8246 12642 8274 12727
rect 8246 12609 8274 12614
rect 8582 11913 8610 13062
rect 8918 13090 8946 13230
rect 8918 13057 8946 13062
rect 9030 13145 9058 13151
rect 9030 13119 9031 13145
rect 9057 13119 9058 13145
rect 8750 13033 8778 13039
rect 8750 13007 8751 13033
rect 8777 13007 8778 13033
rect 8750 12978 8778 13007
rect 8638 12698 8666 12703
rect 8638 12651 8666 12670
rect 8750 12642 8778 12950
rect 9030 12866 9058 13119
rect 9086 13146 9114 13151
rect 9086 13099 9114 13118
rect 9198 13145 9226 13151
rect 9198 13119 9199 13145
rect 9225 13119 9226 13145
rect 9030 12833 9058 12838
rect 9030 12698 9058 12703
rect 9058 12670 9114 12698
rect 9030 12665 9058 12670
rect 8750 12614 8946 12642
rect 8582 11887 8583 11913
rect 8609 11887 8610 11913
rect 8582 11881 8610 11887
rect 8694 11969 8722 11975
rect 8694 11943 8695 11969
rect 8721 11943 8722 11969
rect 7966 11551 7967 11577
rect 7993 11551 7994 11577
rect 6622 10934 6930 10962
rect 7518 10990 7602 11018
rect 7630 11074 7658 11079
rect 6622 10849 6650 10934
rect 6622 10823 6623 10849
rect 6649 10823 6650 10849
rect 6622 10817 6650 10823
rect 5558 10711 5559 10737
rect 5585 10711 5586 10737
rect 5558 10705 5586 10711
rect 7014 10793 7042 10799
rect 7014 10767 7015 10793
rect 7041 10767 7042 10793
rect 7014 10738 7042 10767
rect 7238 10738 7266 10743
rect 7014 10737 7266 10738
rect 7014 10711 7239 10737
rect 7265 10711 7266 10737
rect 7014 10710 7266 10711
rect 2238 10598 2370 10603
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2238 10565 2370 10570
rect 7070 10457 7098 10463
rect 7070 10431 7071 10457
rect 7097 10431 7098 10457
rect 6006 10402 6034 10407
rect 6006 10065 6034 10374
rect 7070 10402 7098 10431
rect 7238 10458 7266 10710
rect 7350 10458 7378 10463
rect 7238 10430 7350 10458
rect 7070 10369 7098 10374
rect 6846 10289 6874 10295
rect 6846 10263 6847 10289
rect 6873 10263 6874 10289
rect 6846 10094 6874 10263
rect 6006 10039 6007 10065
rect 6033 10039 6034 10065
rect 6006 10033 6034 10039
rect 6734 10066 6874 10094
rect 5614 10010 5642 10015
rect 2086 9921 2114 9926
rect 5558 10009 5642 10010
rect 5558 9983 5615 10009
rect 5641 9983 5642 10009
rect 5558 9982 5642 9983
rect 2238 9814 2370 9819
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2238 9781 2370 9786
rect 5558 9226 5586 9982
rect 5614 9977 5642 9982
rect 6734 9673 6762 10066
rect 7070 10010 7098 10015
rect 7238 10010 7266 10015
rect 7070 9954 7098 9982
rect 7014 9953 7098 9954
rect 7014 9927 7071 9953
rect 7097 9927 7098 9953
rect 7014 9926 7098 9927
rect 6734 9647 6735 9673
rect 6761 9647 6762 9673
rect 6734 9641 6762 9647
rect 6902 9674 6930 9679
rect 7014 9674 7042 9926
rect 7070 9921 7098 9926
rect 7126 10009 7266 10010
rect 7126 9983 7239 10009
rect 7265 9983 7266 10009
rect 7126 9982 7266 9983
rect 6902 9673 7042 9674
rect 6902 9647 6903 9673
rect 6929 9647 7042 9673
rect 6902 9646 7042 9647
rect 6902 9641 6930 9646
rect 7070 9618 7098 9623
rect 7126 9618 7154 9982
rect 7238 9977 7266 9982
rect 5558 9179 5586 9198
rect 6958 9617 7154 9618
rect 6958 9591 7071 9617
rect 7097 9591 7154 9617
rect 6958 9590 7154 9591
rect 5894 9169 5922 9175
rect 5894 9143 5895 9169
rect 5921 9143 5922 9169
rect 2238 9030 2370 9035
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2238 8997 2370 9002
rect 2142 8441 2170 8447
rect 2142 8415 2143 8441
rect 2169 8415 2170 8441
rect 966 8329 994 8335
rect 966 8303 967 8329
rect 993 8303 994 8329
rect 966 8106 994 8303
rect 2142 8162 2170 8415
rect 5614 8385 5642 8391
rect 5614 8359 5615 8385
rect 5641 8359 5642 8385
rect 2238 8246 2370 8251
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2238 8213 2370 8218
rect 2142 8129 2170 8134
rect 966 8073 994 8078
rect 1022 8105 1050 8111
rect 1022 8079 1023 8105
rect 1049 8079 1050 8105
rect 1022 7770 1050 8079
rect 2142 8050 2170 8055
rect 2142 8003 2170 8022
rect 5614 8050 5642 8359
rect 5614 7826 5642 8022
rect 5614 7793 5642 7798
rect 5670 8162 5698 8167
rect 1022 7737 1050 7742
rect 5670 7770 5698 8134
rect 5894 8050 5922 9143
rect 6958 9169 6986 9590
rect 7070 9585 7098 9590
rect 6958 9143 6959 9169
rect 6985 9143 6986 9169
rect 6958 9137 6986 9143
rect 7182 9226 7210 9231
rect 7350 9226 7378 10430
rect 7518 10458 7546 10990
rect 7518 10425 7546 10430
rect 7406 10066 7434 10071
rect 7406 10019 7434 10038
rect 7574 10010 7602 10015
rect 7574 9963 7602 9982
rect 7210 9198 7378 9226
rect 7182 8890 7210 9198
rect 7070 8889 7210 8890
rect 7070 8863 7183 8889
rect 7209 8863 7210 8889
rect 7070 8862 7210 8863
rect 7014 8554 7042 8559
rect 6678 8386 6706 8391
rect 6678 8385 6986 8386
rect 6678 8359 6679 8385
rect 6705 8359 6986 8385
rect 6678 8358 6986 8359
rect 6678 8353 6706 8358
rect 6958 8105 6986 8358
rect 6958 8079 6959 8105
rect 6985 8079 6986 8105
rect 6958 8073 6986 8079
rect 5894 8017 5922 8022
rect 6902 8050 6930 8055
rect 6902 8003 6930 8022
rect 7014 8049 7042 8526
rect 7014 8023 7015 8049
rect 7041 8023 7042 8049
rect 7014 8017 7042 8023
rect 7070 8441 7098 8862
rect 7182 8857 7210 8862
rect 7518 8554 7546 8559
rect 7630 8554 7658 11046
rect 7966 10906 7994 11551
rect 8582 11466 8610 11471
rect 8358 11185 8386 11191
rect 8358 11159 8359 11185
rect 8385 11159 8386 11185
rect 8246 11074 8274 11079
rect 8246 11027 8274 11046
rect 8358 10962 8386 11159
rect 8582 11130 8610 11438
rect 8358 10929 8386 10934
rect 8470 11129 8610 11130
rect 8470 11103 8583 11129
rect 8609 11103 8610 11129
rect 8470 11102 8610 11103
rect 7966 10873 7994 10878
rect 8414 10850 8442 10855
rect 8414 10803 8442 10822
rect 8302 10793 8330 10799
rect 8302 10767 8303 10793
rect 8329 10767 8330 10793
rect 7854 10458 7882 10463
rect 7854 10411 7882 10430
rect 8302 10094 8330 10767
rect 7742 10065 7770 10071
rect 7742 10039 7743 10065
rect 7769 10039 7770 10065
rect 7742 9842 7770 10039
rect 7742 9617 7770 9814
rect 7742 9591 7743 9617
rect 7769 9591 7770 9617
rect 7742 9585 7770 9591
rect 7910 10066 7938 10071
rect 7910 9953 7938 10038
rect 8190 10066 8218 10071
rect 8302 10066 8442 10094
rect 8190 10019 8218 10038
rect 8022 10010 8050 10015
rect 8022 9963 8050 9982
rect 7910 9927 7911 9953
rect 7937 9927 7938 9953
rect 7910 9562 7938 9927
rect 8414 9842 8442 10066
rect 7910 9338 7938 9534
rect 7966 9617 7994 9623
rect 7966 9591 7967 9617
rect 7993 9591 7994 9617
rect 7966 9450 7994 9591
rect 8414 9617 8442 9814
rect 8414 9591 8415 9617
rect 8441 9591 8442 9617
rect 8414 9585 8442 9591
rect 7966 9417 7994 9422
rect 8022 9338 8050 9343
rect 7910 9337 8050 9338
rect 7910 9311 8023 9337
rect 8049 9311 8050 9337
rect 7910 9310 8050 9311
rect 8022 9305 8050 9310
rect 8190 9281 8218 9287
rect 8190 9255 8191 9281
rect 8217 9255 8218 9281
rect 8190 9170 8218 9255
rect 8190 9137 8218 9142
rect 8302 8722 8330 8727
rect 7518 8553 7630 8554
rect 7518 8527 7519 8553
rect 7545 8527 7630 8553
rect 7518 8526 7630 8527
rect 7518 8521 7546 8526
rect 7630 8507 7658 8526
rect 8190 8554 8218 8559
rect 8190 8507 8218 8526
rect 8302 8553 8330 8694
rect 8302 8527 8303 8553
rect 8329 8527 8330 8553
rect 8302 8521 8330 8527
rect 7070 8415 7071 8441
rect 7097 8415 7098 8441
rect 7070 8106 7098 8415
rect 6790 7938 6818 7943
rect 6790 7937 6874 7938
rect 6790 7911 6791 7937
rect 6817 7911 6874 7937
rect 6790 7910 6874 7911
rect 6790 7905 6818 7910
rect 5670 7601 5698 7742
rect 6790 7714 6818 7719
rect 6734 7686 6790 7714
rect 6734 7657 6762 7686
rect 6790 7681 6818 7686
rect 6734 7631 6735 7657
rect 6761 7631 6762 7657
rect 6734 7625 6762 7631
rect 5670 7575 5671 7601
rect 5697 7575 5698 7601
rect 5670 7569 5698 7575
rect 2238 7462 2370 7467
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2238 7429 2370 7434
rect 6846 7377 6874 7910
rect 6846 7351 6847 7377
rect 6873 7351 6874 7377
rect 6846 7345 6874 7351
rect 6902 7826 6930 7831
rect 6902 7209 6930 7798
rect 7070 7657 7098 8078
rect 7238 8441 7266 8447
rect 7238 8415 7239 8441
rect 7265 8415 7266 8441
rect 7238 7769 7266 8415
rect 7406 8442 7434 8447
rect 7406 8395 7434 8414
rect 8414 8441 8442 8447
rect 8414 8415 8415 8441
rect 8441 8415 8442 8441
rect 7462 8385 7490 8391
rect 7462 8359 7463 8385
rect 7489 8359 7490 8385
rect 7238 7743 7239 7769
rect 7265 7743 7266 7769
rect 7238 7737 7266 7743
rect 7294 7770 7322 7775
rect 7294 7723 7322 7742
rect 7462 7714 7490 8359
rect 8358 8385 8386 8391
rect 8358 8359 8359 8385
rect 8385 8359 8386 8385
rect 8358 8218 8386 8359
rect 7910 8190 8386 8218
rect 7518 8106 7546 8111
rect 7518 8050 7546 8078
rect 7910 8105 7938 8190
rect 7910 8079 7911 8105
rect 7937 8079 7938 8105
rect 7910 8073 7938 8079
rect 8414 8106 8442 8415
rect 8414 8073 8442 8078
rect 7518 8049 7770 8050
rect 7518 8023 7519 8049
rect 7545 8023 7770 8049
rect 7518 8022 7770 8023
rect 7518 8017 7546 8022
rect 7462 7681 7490 7686
rect 7518 7770 7546 7775
rect 7518 7713 7546 7742
rect 7518 7687 7519 7713
rect 7545 7687 7546 7713
rect 7070 7631 7071 7657
rect 7097 7631 7098 7657
rect 7014 7546 7042 7551
rect 7014 7265 7042 7518
rect 7014 7239 7015 7265
rect 7041 7239 7042 7265
rect 7014 7233 7042 7239
rect 6902 7183 6903 7209
rect 6929 7183 6930 7209
rect 6902 7177 6930 7183
rect 7014 6874 7042 6879
rect 7070 6874 7098 7631
rect 7350 7658 7378 7663
rect 7182 7602 7210 7607
rect 7182 7265 7210 7574
rect 7182 7239 7183 7265
rect 7209 7239 7210 7265
rect 7182 7233 7210 7239
rect 7350 6929 7378 7630
rect 7406 7657 7434 7663
rect 7406 7631 7407 7657
rect 7433 7631 7434 7657
rect 7406 7546 7434 7631
rect 7518 7602 7546 7687
rect 7518 7569 7546 7574
rect 7742 7769 7770 8022
rect 7742 7743 7743 7769
rect 7769 7743 7770 7769
rect 7742 7602 7770 7743
rect 7742 7569 7770 7574
rect 7406 7513 7434 7518
rect 8470 7546 8498 11102
rect 8582 11097 8610 11102
rect 8638 11242 8666 11247
rect 8582 10906 8610 10911
rect 8526 9618 8554 9623
rect 8526 9561 8554 9590
rect 8526 9535 8527 9561
rect 8553 9535 8554 9561
rect 8526 9529 8554 9535
rect 8582 9338 8610 10878
rect 8638 9729 8666 11214
rect 8694 10962 8722 11943
rect 8750 11186 8778 11191
rect 8750 11139 8778 11158
rect 8918 11129 8946 12614
rect 9086 12473 9114 12670
rect 9086 12447 9087 12473
rect 9113 12447 9114 12473
rect 9086 12441 9114 12447
rect 9142 12474 9170 12479
rect 9142 12427 9170 12446
rect 9030 12361 9058 12367
rect 9030 12335 9031 12361
rect 9057 12335 9058 12361
rect 9030 11746 9058 12335
rect 9030 11713 9058 11718
rect 9198 11690 9226 13119
rect 9366 12361 9394 13399
rect 9534 13425 9562 13431
rect 9534 13399 9535 13425
rect 9561 13399 9562 13425
rect 9422 13090 9450 13095
rect 9534 13090 9562 13399
rect 9590 13145 9618 13151
rect 9590 13119 9591 13145
rect 9617 13119 9618 13145
rect 9590 13090 9618 13119
rect 9422 13089 9618 13090
rect 9422 13063 9423 13089
rect 9449 13063 9618 13089
rect 9422 13062 9618 13063
rect 9422 12642 9450 13062
rect 9422 12609 9450 12614
rect 9534 12866 9562 12871
rect 9366 12335 9367 12361
rect 9393 12335 9394 12361
rect 9366 12329 9394 12335
rect 9310 11690 9338 11695
rect 9198 11662 9310 11690
rect 9310 11643 9338 11662
rect 9478 11578 9506 11583
rect 9198 11242 9226 11247
rect 9198 11195 9226 11214
rect 9086 11186 9114 11191
rect 8918 11103 8919 11129
rect 8945 11103 8946 11129
rect 8918 11097 8946 11103
rect 8974 11185 9114 11186
rect 8974 11159 9087 11185
rect 9113 11159 9114 11185
rect 8974 11158 9114 11159
rect 8750 10962 8778 10967
rect 8974 10962 9002 11158
rect 9086 11153 9114 11158
rect 9478 11186 9506 11550
rect 9478 11139 9506 11158
rect 8694 10934 8750 10962
rect 8750 10905 8778 10934
rect 8750 10879 8751 10905
rect 8777 10879 8778 10905
rect 8750 10873 8778 10879
rect 8806 10934 9002 10962
rect 9422 10962 9450 10967
rect 8806 10905 8834 10934
rect 8806 10879 8807 10905
rect 8833 10879 8834 10905
rect 8750 9954 8778 9959
rect 8750 9907 8778 9926
rect 8806 9730 8834 10879
rect 8638 9703 8639 9729
rect 8665 9703 8666 9729
rect 8638 9697 8666 9703
rect 8750 9702 8834 9730
rect 8862 10850 8890 10855
rect 8750 9618 8778 9702
rect 8694 9506 8722 9511
rect 8694 9459 8722 9478
rect 8638 9338 8666 9343
rect 8582 9337 8666 9338
rect 8582 9311 8639 9337
rect 8665 9311 8666 9337
rect 8582 9310 8666 9311
rect 8638 9305 8666 9310
rect 8750 9226 8778 9590
rect 8806 9618 8834 9623
rect 8862 9618 8890 10822
rect 9366 10850 9394 10855
rect 9366 10803 9394 10822
rect 8806 9617 8890 9618
rect 8806 9591 8807 9617
rect 8833 9591 8890 9617
rect 8806 9590 8890 9591
rect 8918 10793 8946 10799
rect 8918 10767 8919 10793
rect 8945 10767 8946 10793
rect 8806 9585 8834 9590
rect 8750 9193 8778 9198
rect 8862 9450 8890 9455
rect 8862 9225 8890 9422
rect 8918 9338 8946 10767
rect 9086 10794 9114 10799
rect 9086 10747 9114 10766
rect 9366 10402 9394 10407
rect 9366 10122 9394 10374
rect 9086 10010 9114 10015
rect 9086 9953 9114 9982
rect 9086 9927 9087 9953
rect 9113 9927 9114 9953
rect 9086 9921 9114 9927
rect 9142 10009 9170 10015
rect 9142 9983 9143 10009
rect 9169 9983 9170 10009
rect 9142 9842 9170 9983
rect 9254 10010 9282 10015
rect 9254 10009 9338 10010
rect 9254 9983 9255 10009
rect 9281 9983 9338 10009
rect 9254 9982 9338 9983
rect 9254 9977 9282 9982
rect 9254 9898 9282 9903
rect 9142 9809 9170 9814
rect 9198 9870 9254 9898
rect 8974 9618 9002 9623
rect 8974 9571 9002 9590
rect 8918 9305 8946 9310
rect 8974 9506 9002 9511
rect 8862 9199 8863 9225
rect 8889 9199 8890 9225
rect 8862 7826 8890 9199
rect 8974 9225 9002 9478
rect 8974 9199 8975 9225
rect 9001 9199 9002 9225
rect 8918 8722 8946 8727
rect 8918 8675 8946 8694
rect 8974 8442 9002 9199
rect 9142 9505 9170 9511
rect 9142 9479 9143 9505
rect 9169 9479 9170 9505
rect 9030 9170 9058 9175
rect 9142 9170 9170 9479
rect 9030 9169 9170 9170
rect 9030 9143 9031 9169
rect 9057 9143 9170 9169
rect 9030 9142 9170 9143
rect 9030 8833 9058 9142
rect 9086 8946 9114 8951
rect 9198 8946 9226 9870
rect 9254 9851 9282 9870
rect 9310 9786 9338 9982
rect 9254 9758 9338 9786
rect 9254 9562 9282 9758
rect 9254 9529 9282 9534
rect 9310 9505 9338 9511
rect 9310 9479 9311 9505
rect 9337 9479 9338 9505
rect 9310 9338 9338 9479
rect 9310 9305 9338 9310
rect 9086 8945 9226 8946
rect 9086 8919 9087 8945
rect 9113 8919 9226 8945
rect 9086 8918 9226 8919
rect 9086 8913 9114 8918
rect 9030 8807 9031 8833
rect 9057 8807 9058 8833
rect 9030 8498 9058 8807
rect 9310 8834 9338 8839
rect 9366 8834 9394 10094
rect 9310 8833 9394 8834
rect 9310 8807 9311 8833
rect 9337 8807 9394 8833
rect 9310 8806 9394 8807
rect 9310 8801 9338 8806
rect 9198 8778 9226 8783
rect 9198 8731 9226 8750
rect 9310 8554 9338 8559
rect 9254 8526 9310 8554
rect 9422 8554 9450 10934
rect 9534 9898 9562 12838
rect 9702 12809 9730 13510
rect 10374 13537 10402 13566
rect 10710 13561 10738 13566
rect 10766 13594 10794 13599
rect 10374 13511 10375 13537
rect 10401 13511 10402 13537
rect 10374 13505 10402 13511
rect 10206 13482 10234 13487
rect 10094 13481 10234 13482
rect 10094 13455 10207 13481
rect 10233 13455 10234 13481
rect 10094 13454 10234 13455
rect 9918 13342 10050 13347
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 9918 13309 10050 13314
rect 10094 13258 10122 13454
rect 10206 13449 10234 13454
rect 10654 13482 10682 13487
rect 10766 13482 10794 13566
rect 10822 13537 10850 13958
rect 10822 13511 10823 13537
rect 10849 13511 10850 13537
rect 10822 13505 10850 13511
rect 10654 13481 10794 13482
rect 10654 13455 10655 13481
rect 10681 13455 10794 13481
rect 10654 13454 10794 13455
rect 10934 13481 10962 13487
rect 10934 13455 10935 13481
rect 10961 13455 10962 13481
rect 10654 13449 10682 13454
rect 9982 13230 10122 13258
rect 10318 13425 10346 13431
rect 10318 13399 10319 13425
rect 10345 13399 10346 13425
rect 9982 13201 10010 13230
rect 9982 13175 9983 13201
rect 10009 13175 10010 13201
rect 9982 13169 10010 13175
rect 10318 12865 10346 13399
rect 10934 13426 10962 13455
rect 10318 12839 10319 12865
rect 10345 12839 10346 12865
rect 10318 12833 10346 12839
rect 10654 12866 10682 12871
rect 10654 12819 10682 12838
rect 9702 12783 9703 12809
rect 9729 12783 9730 12809
rect 9702 12777 9730 12783
rect 10822 12810 10850 12815
rect 10822 12763 10850 12782
rect 10598 12754 10626 12759
rect 10374 12698 10402 12703
rect 10374 12697 10570 12698
rect 10374 12671 10375 12697
rect 10401 12671 10570 12697
rect 10374 12670 10570 12671
rect 10374 12665 10402 12670
rect 9926 12642 9954 12661
rect 10318 12642 10346 12647
rect 9926 12609 9954 12614
rect 10262 12641 10346 12642
rect 10262 12615 10319 12641
rect 10345 12615 10346 12641
rect 10262 12614 10346 12615
rect 9918 12558 10050 12563
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 9918 12525 10050 12530
rect 10262 12474 10290 12614
rect 10318 12609 10346 12614
rect 9918 11774 10050 11779
rect 9758 11746 9786 11751
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 9918 11741 10050 11746
rect 9758 11689 9786 11718
rect 9758 11663 9759 11689
rect 9785 11663 9786 11689
rect 9646 11633 9674 11639
rect 9646 11607 9647 11633
rect 9673 11607 9674 11633
rect 9590 11465 9618 11471
rect 9590 11439 9591 11465
rect 9617 11439 9618 11465
rect 9590 11354 9618 11439
rect 9590 11321 9618 11326
rect 9646 11298 9674 11607
rect 9646 11265 9674 11270
rect 9758 10962 9786 11663
rect 9870 11634 9898 11639
rect 9702 10906 9730 10911
rect 9758 10906 9786 10934
rect 9702 10905 9786 10906
rect 9702 10879 9703 10905
rect 9729 10879 9786 10905
rect 9702 10878 9786 10879
rect 9814 11633 9898 11634
rect 9814 11607 9871 11633
rect 9897 11607 9898 11633
rect 9814 11606 9898 11607
rect 9702 10873 9730 10878
rect 9534 9865 9562 9870
rect 9646 10849 9674 10855
rect 9646 10823 9647 10849
rect 9673 10823 9674 10849
rect 9478 9506 9506 9511
rect 9478 9459 9506 9478
rect 9646 9505 9674 10823
rect 9814 10850 9842 11606
rect 9870 11601 9898 11606
rect 10150 11578 10178 11583
rect 10094 11521 10122 11527
rect 10094 11495 10095 11521
rect 10121 11495 10122 11521
rect 10094 11185 10122 11495
rect 10094 11159 10095 11185
rect 10121 11159 10122 11185
rect 9918 10990 10050 10995
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 9918 10957 10050 10962
rect 9814 10822 9898 10850
rect 9758 10794 9786 10799
rect 9758 10747 9786 10766
rect 9870 10682 9898 10822
rect 9870 10649 9898 10654
rect 10038 10401 10066 10407
rect 10038 10375 10039 10401
rect 10065 10375 10066 10401
rect 10038 10346 10066 10375
rect 10038 10313 10066 10318
rect 9918 10206 10050 10211
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 9918 10173 10050 10178
rect 10094 10066 10122 11159
rect 10150 10905 10178 11550
rect 10150 10879 10151 10905
rect 10177 10879 10178 10905
rect 10150 10873 10178 10879
rect 10094 10033 10122 10038
rect 9702 10009 9730 10015
rect 9702 9983 9703 10009
rect 9729 9983 9730 10009
rect 9702 9954 9730 9983
rect 9702 9921 9730 9926
rect 9870 9786 9898 9791
rect 9646 9479 9647 9505
rect 9673 9479 9674 9505
rect 9646 9170 9674 9479
rect 9814 9758 9870 9786
rect 9814 9338 9842 9758
rect 9870 9753 9898 9758
rect 10038 9730 10066 9735
rect 10038 9617 10066 9702
rect 10038 9591 10039 9617
rect 10065 9591 10066 9617
rect 10038 9585 10066 9591
rect 9870 9506 9898 9511
rect 9870 9505 10122 9506
rect 9870 9479 9871 9505
rect 9897 9479 10122 9505
rect 9870 9478 10122 9479
rect 9870 9473 9898 9478
rect 9918 9422 10050 9427
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 9918 9389 10050 9394
rect 10094 9338 10122 9478
rect 9814 9310 9954 9338
rect 9758 9226 9786 9231
rect 9870 9226 9898 9231
rect 9786 9198 9842 9226
rect 9758 9179 9786 9198
rect 9646 9123 9674 9142
rect 9590 9114 9618 9119
rect 9422 8526 9506 8554
rect 9142 8498 9170 8503
rect 9030 8470 9142 8498
rect 8974 8395 9002 8414
rect 9142 8441 9170 8470
rect 9254 8442 9282 8526
rect 9310 8521 9338 8526
rect 9422 8442 9450 8447
rect 9142 8415 9143 8441
rect 9169 8415 9170 8441
rect 9142 8409 9170 8415
rect 9198 8414 9282 8442
rect 9310 8441 9450 8442
rect 9310 8415 9423 8441
rect 9449 8415 9450 8441
rect 9310 8414 9450 8415
rect 9198 8385 9226 8414
rect 9198 8359 9199 8385
rect 9225 8359 9226 8385
rect 9198 8353 9226 8359
rect 9254 8330 9282 8335
rect 9254 8283 9282 8302
rect 8862 7793 8890 7798
rect 8974 8105 9002 8111
rect 8974 8079 8975 8105
rect 9001 8079 9002 8105
rect 8974 8050 9002 8079
rect 9142 8050 9170 8055
rect 8974 8049 9170 8050
rect 8974 8023 9143 8049
rect 9169 8023 9170 8049
rect 8974 8022 9170 8023
rect 8806 7658 8834 7663
rect 8750 7657 8834 7658
rect 8750 7631 8807 7657
rect 8833 7631 8834 7657
rect 8750 7630 8834 7631
rect 8470 7266 8498 7518
rect 8694 7546 8722 7551
rect 8582 7266 8610 7271
rect 8470 7265 8610 7266
rect 8470 7239 8583 7265
rect 8609 7239 8610 7265
rect 8470 7238 8610 7239
rect 8582 7233 8610 7238
rect 8638 7153 8666 7159
rect 8638 7127 8639 7153
rect 8665 7127 8666 7153
rect 8638 7042 8666 7127
rect 7350 6903 7351 6929
rect 7377 6903 7378 6929
rect 7350 6897 7378 6903
rect 8526 7014 8666 7042
rect 7014 6873 7098 6874
rect 7014 6847 7015 6873
rect 7041 6847 7098 6873
rect 7014 6846 7098 6847
rect 7014 6841 7042 6846
rect 8414 6818 8442 6823
rect 8526 6818 8554 7014
rect 8694 6986 8722 7518
rect 8750 7209 8778 7630
rect 8806 7625 8834 7630
rect 8918 7658 8946 7663
rect 8918 7611 8946 7630
rect 8974 7266 9002 8022
rect 9142 8017 9170 8022
rect 9310 8049 9338 8414
rect 9422 8409 9450 8414
rect 9310 8023 9311 8049
rect 9337 8023 9338 8049
rect 9310 8017 9338 8023
rect 9366 8274 9394 8279
rect 9366 8049 9394 8246
rect 9422 8106 9450 8111
rect 9422 8059 9450 8078
rect 9366 8023 9367 8049
rect 9393 8023 9394 8049
rect 9366 8017 9394 8023
rect 9478 8049 9506 8526
rect 9534 8498 9562 8503
rect 9534 8451 9562 8470
rect 9590 8497 9618 9086
rect 9814 8834 9842 9198
rect 9870 9179 9898 9198
rect 9926 8945 9954 9310
rect 10038 9310 10122 9338
rect 10206 9505 10234 9511
rect 10206 9479 10207 9505
rect 10233 9479 10234 9505
rect 10206 9338 10234 9479
rect 9926 8919 9927 8945
rect 9953 8919 9954 8945
rect 9926 8913 9954 8919
rect 9982 9170 10010 9175
rect 9870 8834 9898 8839
rect 9814 8833 9898 8834
rect 9814 8807 9871 8833
rect 9897 8807 9898 8833
rect 9814 8806 9898 8807
rect 9870 8801 9898 8806
rect 9590 8471 9591 8497
rect 9617 8471 9618 8497
rect 9590 8465 9618 8471
rect 9702 8778 9730 8783
rect 9702 8442 9730 8750
rect 9926 8778 9954 8783
rect 9982 8778 10010 9142
rect 10038 9002 10066 9310
rect 10206 9305 10234 9310
rect 10094 9114 10122 9119
rect 10094 9067 10122 9086
rect 10038 8974 10122 9002
rect 9926 8777 10010 8778
rect 9926 8751 9927 8777
rect 9953 8751 10010 8777
rect 9926 8750 10010 8751
rect 9926 8745 9954 8750
rect 9918 8638 10050 8643
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 9918 8605 10050 8610
rect 9478 8023 9479 8049
rect 9505 8023 9506 8049
rect 9030 7938 9058 7943
rect 9030 7713 9058 7910
rect 9478 7938 9506 8023
rect 9478 7905 9506 7910
rect 9590 8330 9618 8335
rect 9478 7826 9506 7831
rect 9030 7687 9031 7713
rect 9057 7687 9058 7713
rect 9030 7681 9058 7687
rect 9142 7714 9170 7719
rect 9142 7667 9170 7686
rect 9478 7713 9506 7798
rect 9590 7770 9618 8302
rect 9478 7687 9479 7713
rect 9505 7687 9506 7713
rect 9478 7681 9506 7687
rect 9534 7769 9618 7770
rect 9534 7743 9591 7769
rect 9617 7743 9618 7769
rect 9534 7742 9618 7743
rect 9702 7770 9730 8414
rect 10094 8050 10122 8974
rect 10262 8274 10290 12446
rect 10542 11970 10570 12670
rect 10542 11633 10570 11942
rect 10542 11607 10543 11633
rect 10569 11607 10570 11633
rect 10542 11601 10570 11607
rect 10318 11577 10346 11583
rect 10318 11551 10319 11577
rect 10345 11551 10346 11577
rect 10318 10906 10346 11551
rect 10374 11354 10402 11359
rect 10374 11241 10402 11326
rect 10374 11215 10375 11241
rect 10401 11215 10402 11241
rect 10374 11209 10402 11215
rect 10318 10873 10346 10878
rect 10374 11074 10402 11079
rect 10318 10793 10346 10799
rect 10318 10767 10319 10793
rect 10345 10767 10346 10793
rect 10318 10458 10346 10767
rect 10318 10425 10346 10430
rect 10374 10010 10402 11046
rect 10374 9617 10402 9982
rect 10374 9591 10375 9617
rect 10401 9591 10402 9617
rect 10374 9585 10402 9591
rect 10486 10906 10514 10911
rect 10430 9338 10458 9343
rect 10430 9291 10458 9310
rect 10486 8553 10514 10878
rect 10598 10905 10626 12726
rect 10878 12754 10906 12759
rect 10934 12754 10962 13398
rect 10906 12726 10962 12754
rect 10990 13482 11018 13487
rect 10878 12721 10906 12726
rect 10990 12697 11018 13454
rect 11046 13089 11074 13958
rect 11774 13930 11802 13935
rect 11662 13874 11690 13879
rect 11662 13827 11690 13846
rect 11550 13818 11578 13823
rect 11382 13594 11410 13599
rect 11410 13566 11466 13594
rect 11382 13561 11410 13566
rect 11326 13537 11354 13543
rect 11326 13511 11327 13537
rect 11353 13511 11354 13537
rect 11102 13481 11130 13487
rect 11102 13455 11103 13481
rect 11129 13455 11130 13481
rect 11102 13146 11130 13455
rect 11214 13481 11242 13487
rect 11214 13455 11215 13481
rect 11241 13455 11242 13481
rect 11214 13258 11242 13455
rect 11326 13426 11354 13511
rect 11438 13537 11466 13566
rect 11438 13511 11439 13537
rect 11465 13511 11466 13537
rect 11438 13505 11466 13511
rect 11550 13537 11578 13790
rect 11550 13511 11551 13537
rect 11577 13511 11578 13537
rect 11550 13505 11578 13511
rect 11774 13538 11802 13902
rect 11774 13505 11802 13510
rect 11326 13393 11354 13398
rect 11606 13482 11634 13487
rect 11606 13425 11634 13454
rect 11606 13399 11607 13425
rect 11633 13399 11634 13425
rect 11606 13393 11634 13399
rect 11774 13426 11802 13431
rect 11214 13230 11746 13258
rect 11102 13113 11130 13118
rect 11158 13202 11186 13207
rect 11046 13063 11047 13089
rect 11073 13063 11074 13089
rect 11046 13057 11074 13063
rect 11158 12810 11186 13174
rect 11158 12753 11186 12782
rect 11158 12727 11159 12753
rect 11185 12727 11186 12753
rect 11158 12721 11186 12727
rect 10990 12671 10991 12697
rect 11017 12671 11018 12697
rect 10990 12665 11018 12671
rect 10766 12641 10794 12647
rect 10766 12615 10767 12641
rect 10793 12615 10794 12641
rect 10710 12474 10738 12479
rect 10710 12427 10738 12446
rect 10766 12362 10794 12615
rect 10822 12362 10850 12367
rect 10766 12361 10850 12362
rect 10766 12335 10823 12361
rect 10849 12335 10850 12361
rect 10766 12334 10850 12335
rect 10766 11969 10794 11975
rect 10766 11943 10767 11969
rect 10793 11943 10794 11969
rect 10766 11914 10794 11943
rect 10766 11881 10794 11886
rect 10710 11578 10738 11583
rect 10822 11578 10850 12334
rect 10878 11913 10906 11919
rect 10878 11887 10879 11913
rect 10905 11887 10906 11913
rect 10878 11690 10906 11887
rect 11046 11914 11074 11919
rect 11074 11886 11130 11914
rect 11046 11881 11074 11886
rect 10878 11662 10962 11690
rect 10934 11634 10962 11662
rect 10878 11578 10906 11583
rect 10822 11550 10878 11578
rect 10710 11531 10738 11550
rect 10878 11545 10906 11550
rect 10934 11466 10962 11606
rect 11046 11633 11074 11639
rect 11046 11607 11047 11633
rect 11073 11607 11074 11633
rect 10878 11438 10962 11466
rect 10990 11577 11018 11583
rect 10990 11551 10991 11577
rect 11017 11551 11018 11577
rect 10878 11130 10906 11438
rect 10990 11354 11018 11551
rect 10990 11321 11018 11326
rect 11046 11242 11074 11607
rect 11102 11298 11130 11886
rect 11158 11913 11186 11919
rect 11158 11887 11159 11913
rect 11185 11887 11186 11913
rect 11158 11522 11186 11887
rect 11214 11857 11242 13230
rect 11214 11831 11215 11857
rect 11241 11831 11242 11857
rect 11214 11825 11242 11831
rect 11270 13146 11298 13151
rect 11158 11489 11186 11494
rect 11214 11522 11242 11527
rect 11270 11522 11298 13118
rect 11718 13145 11746 13230
rect 11718 13119 11719 13145
rect 11745 13119 11746 13145
rect 11718 13113 11746 13119
rect 11774 13201 11802 13398
rect 11830 13257 11858 14238
rect 11942 13930 11970 13935
rect 11942 13883 11970 13902
rect 12278 13874 12306 18999
rect 13398 18745 13426 19278
rect 17598 19222 17730 19227
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17598 19189 17730 19194
rect 14686 19138 14714 19143
rect 14686 19091 14714 19110
rect 13398 18719 13399 18745
rect 13425 18719 13426 18745
rect 13398 18713 13426 18719
rect 14294 19025 14322 19031
rect 14294 18999 14295 19025
rect 14321 18999 14322 19025
rect 12950 18633 12978 18639
rect 12950 18607 12951 18633
rect 12977 18607 12978 18633
rect 12950 14042 12978 18607
rect 13118 14042 13146 14047
rect 12670 14041 13090 14042
rect 12670 14015 12951 14041
rect 12977 14015 13090 14041
rect 12670 14014 13090 14015
rect 12670 13985 12698 14014
rect 12950 14009 12978 14014
rect 12670 13959 12671 13985
rect 12697 13959 12698 13985
rect 12670 13953 12698 13959
rect 13062 13930 13090 14014
rect 13118 13995 13146 14014
rect 14294 14042 14322 18999
rect 17598 18438 17730 18443
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17598 18405 17730 18410
rect 17598 17654 17730 17659
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17598 17621 17730 17626
rect 17598 16870 17730 16875
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17598 16837 17730 16842
rect 17598 16086 17730 16091
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17598 16053 17730 16058
rect 17598 15302 17730 15307
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17598 15269 17730 15274
rect 17598 14518 17730 14523
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17598 14485 17730 14490
rect 14294 14009 14322 14014
rect 13062 13902 13202 13930
rect 12222 13846 12278 13874
rect 12110 13482 12138 13487
rect 12110 13435 12138 13454
rect 11830 13231 11831 13257
rect 11857 13231 11858 13257
rect 11830 13225 11858 13231
rect 11774 13175 11775 13201
rect 11801 13175 11802 13201
rect 11774 12810 11802 13175
rect 12110 13202 12138 13207
rect 12110 13155 12138 13174
rect 12222 13145 12250 13846
rect 12278 13841 12306 13846
rect 12614 13818 12642 13823
rect 12614 13771 12642 13790
rect 13174 13593 13202 13902
rect 17598 13734 17730 13739
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17598 13701 17730 13706
rect 13174 13567 13175 13593
rect 13201 13567 13202 13593
rect 13174 13561 13202 13567
rect 20006 13593 20034 13599
rect 20006 13567 20007 13593
rect 20033 13567 20034 13593
rect 12222 13119 12223 13145
rect 12249 13119 12250 13145
rect 12222 13113 12250 13119
rect 12614 13538 12642 13543
rect 12614 13145 12642 13510
rect 13398 13538 13426 13543
rect 13398 13258 13426 13510
rect 18830 13537 18858 13543
rect 18830 13511 18831 13537
rect 18857 13511 18858 13537
rect 13398 13225 13426 13230
rect 13678 13258 13706 13263
rect 12614 13119 12615 13145
rect 12641 13119 12642 13145
rect 12614 13113 12642 13119
rect 13286 13146 13314 13151
rect 12278 13090 12306 13095
rect 11774 12782 12082 12810
rect 12054 12753 12082 12782
rect 12278 12809 12306 13062
rect 13006 13090 13034 13095
rect 13006 13043 13034 13062
rect 12278 12783 12279 12809
rect 12305 12783 12306 12809
rect 12278 12777 12306 12783
rect 12054 12727 12055 12753
rect 12081 12727 12082 12753
rect 12054 12721 12082 12727
rect 12334 12754 12362 12759
rect 12334 12707 12362 12726
rect 13174 12754 13202 12759
rect 13174 12707 13202 12726
rect 12166 12698 12194 12703
rect 12110 12697 12194 12698
rect 12110 12671 12167 12697
rect 12193 12671 12194 12697
rect 12110 12670 12194 12671
rect 12110 12082 12138 12670
rect 12166 12665 12194 12670
rect 13286 12697 13314 13118
rect 13286 12671 13287 12697
rect 13313 12671 13314 12697
rect 13286 12665 13314 12671
rect 13342 12697 13370 12703
rect 13342 12671 13343 12697
rect 13369 12671 13370 12697
rect 11830 12054 12138 12082
rect 13286 12306 13314 12311
rect 11830 12025 11858 12054
rect 11830 11999 11831 12025
rect 11857 11999 11858 12025
rect 11830 11689 11858 11999
rect 11942 11970 11970 11975
rect 11942 11923 11970 11942
rect 12110 11914 12138 11919
rect 12278 11914 12306 11919
rect 12110 11913 12306 11914
rect 12110 11887 12111 11913
rect 12137 11887 12279 11913
rect 12305 11887 12306 11913
rect 12110 11886 12306 11887
rect 12110 11881 12138 11886
rect 12278 11881 12306 11886
rect 11830 11663 11831 11689
rect 11857 11663 11858 11689
rect 11830 11657 11858 11663
rect 12446 11857 12474 11863
rect 12446 11831 12447 11857
rect 12473 11831 12474 11857
rect 11942 11634 11970 11639
rect 11886 11633 11970 11634
rect 11886 11607 11943 11633
rect 11969 11607 11970 11633
rect 11886 11606 11970 11607
rect 11214 11521 11298 11522
rect 11214 11495 11215 11521
rect 11241 11495 11298 11521
rect 11214 11494 11298 11495
rect 11382 11578 11410 11583
rect 11438 11578 11466 11583
rect 11410 11577 11466 11578
rect 11410 11551 11439 11577
rect 11465 11551 11466 11577
rect 11410 11550 11466 11551
rect 11214 11489 11242 11494
rect 11102 11270 11242 11298
rect 10990 11214 11046 11242
rect 10878 11097 10906 11102
rect 10934 11185 10962 11191
rect 10934 11159 10935 11185
rect 10961 11159 10962 11185
rect 10654 11074 10682 11079
rect 10654 11027 10682 11046
rect 10934 11018 10962 11159
rect 10878 10990 10962 11018
rect 10878 10906 10906 10990
rect 10598 10879 10599 10905
rect 10625 10879 10626 10905
rect 10598 10873 10626 10879
rect 10822 10878 10878 10906
rect 10654 10849 10682 10855
rect 10654 10823 10655 10849
rect 10681 10823 10682 10849
rect 10598 10794 10626 10799
rect 10598 10747 10626 10766
rect 10654 10094 10682 10823
rect 10822 10345 10850 10878
rect 10878 10873 10906 10878
rect 10822 10319 10823 10345
rect 10849 10319 10850 10345
rect 10822 10313 10850 10319
rect 10990 10094 11018 11214
rect 11046 11209 11074 11214
rect 11102 11185 11130 11191
rect 11102 11159 11103 11185
rect 11129 11159 11130 11185
rect 11102 10794 11130 11159
rect 10654 10066 10738 10094
rect 10710 9730 10738 10066
rect 10710 9683 10738 9702
rect 10934 10066 11018 10094
rect 11046 10346 11074 10351
rect 11046 10066 11074 10318
rect 11102 10345 11130 10766
rect 11102 10319 11103 10345
rect 11129 10319 11130 10345
rect 11102 10313 11130 10319
rect 11158 10458 11186 10463
rect 10654 9562 10682 9567
rect 10654 9515 10682 9534
rect 10878 9281 10906 9287
rect 10878 9255 10879 9281
rect 10905 9255 10906 9281
rect 10486 8527 10487 8553
rect 10513 8527 10514 8553
rect 10486 8521 10514 8527
rect 10654 9170 10682 9175
rect 10654 8554 10682 9142
rect 10654 8521 10682 8526
rect 10878 8554 10906 9255
rect 10934 9170 10962 10066
rect 11046 10019 11074 10038
rect 10990 9673 11018 9679
rect 10990 9647 10991 9673
rect 11017 9647 11018 9673
rect 10990 9338 11018 9647
rect 10990 9225 11018 9310
rect 10990 9199 10991 9225
rect 11017 9199 11018 9225
rect 10990 9193 11018 9199
rect 11158 9617 11186 10430
rect 11214 10401 11242 11270
rect 11382 11073 11410 11550
rect 11438 11545 11466 11550
rect 11606 11522 11634 11527
rect 11662 11522 11690 11527
rect 11634 11521 11690 11522
rect 11634 11495 11663 11521
rect 11689 11495 11690 11521
rect 11634 11494 11690 11495
rect 11382 11047 11383 11073
rect 11409 11047 11410 11073
rect 11214 10375 11215 10401
rect 11241 10375 11242 10401
rect 11214 10122 11242 10375
rect 11270 10682 11298 10687
rect 11270 10402 11298 10654
rect 11382 10514 11410 11047
rect 11550 11074 11578 11079
rect 11606 11074 11634 11494
rect 11662 11489 11690 11494
rect 11774 11354 11802 11359
rect 11718 11241 11746 11247
rect 11718 11215 11719 11241
rect 11745 11215 11746 11241
rect 11718 11186 11746 11215
rect 11718 11153 11746 11158
rect 11774 11186 11802 11326
rect 11774 11185 11858 11186
rect 11774 11159 11775 11185
rect 11801 11159 11858 11185
rect 11774 11158 11858 11159
rect 11774 11153 11802 11158
rect 11550 11073 11634 11074
rect 11550 11047 11551 11073
rect 11577 11047 11634 11073
rect 11550 11046 11634 11047
rect 11662 11073 11690 11079
rect 11662 11047 11663 11073
rect 11689 11047 11690 11073
rect 11438 10514 11466 10519
rect 11382 10513 11466 10514
rect 11382 10487 11439 10513
rect 11465 10487 11466 10513
rect 11382 10486 11466 10487
rect 11438 10481 11466 10486
rect 11494 10458 11522 10463
rect 11494 10411 11522 10430
rect 11270 10355 11298 10374
rect 11214 10089 11242 10094
rect 11158 9591 11159 9617
rect 11185 9591 11186 9617
rect 10934 9137 10962 9142
rect 11158 9058 11186 9591
rect 11382 9618 11410 9623
rect 11382 9571 11410 9590
rect 11438 9282 11466 9287
rect 11438 9225 11466 9254
rect 11438 9199 11439 9225
rect 11465 9199 11466 9225
rect 11438 9193 11466 9199
rect 11494 9225 11522 9231
rect 11494 9199 11495 9225
rect 11521 9199 11522 9225
rect 11158 9025 11186 9030
rect 11494 9002 11522 9199
rect 11382 8974 11522 9002
rect 11158 8946 11186 8951
rect 11382 8946 11410 8974
rect 11046 8945 11410 8946
rect 11046 8919 11159 8945
rect 11185 8919 11410 8945
rect 11046 8918 11410 8919
rect 11046 8666 11074 8918
rect 11158 8913 11186 8918
rect 11438 8890 11466 8895
rect 11438 8843 11466 8862
rect 10878 8521 10906 8526
rect 10990 8638 11074 8666
rect 11102 8777 11130 8783
rect 11102 8751 11103 8777
rect 11129 8751 11130 8777
rect 10262 8241 10290 8246
rect 10318 8497 10346 8503
rect 10318 8471 10319 8497
rect 10345 8471 10346 8497
rect 10094 8017 10122 8022
rect 9758 7938 9786 7943
rect 9758 7937 9842 7938
rect 9758 7911 9759 7937
rect 9785 7911 9842 7937
rect 9758 7910 9842 7911
rect 9758 7905 9786 7910
rect 9758 7770 9786 7775
rect 9702 7769 9786 7770
rect 9702 7743 9759 7769
rect 9785 7743 9786 7769
rect 9702 7742 9786 7743
rect 9086 7602 9114 7607
rect 8974 7238 9058 7266
rect 8750 7183 8751 7209
rect 8777 7183 8778 7209
rect 8750 7177 8778 7183
rect 8918 7153 8946 7159
rect 8918 7127 8919 7153
rect 8945 7127 8946 7153
rect 8750 6986 8778 6991
rect 8918 6986 8946 7127
rect 8414 6817 8554 6818
rect 8414 6791 8415 6817
rect 8441 6791 8554 6817
rect 8414 6790 8554 6791
rect 8582 6985 8918 6986
rect 8582 6959 8751 6985
rect 8777 6959 8918 6985
rect 8582 6958 8918 6959
rect 2238 6678 2370 6683
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2238 6645 2370 6650
rect 2238 5894 2370 5899
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2238 5861 2370 5866
rect 8414 5866 8442 6790
rect 8582 6481 8610 6958
rect 8750 6953 8778 6958
rect 8918 6939 8946 6958
rect 8974 7154 9002 7159
rect 8974 6985 9002 7126
rect 8974 6959 8975 6985
rect 9001 6959 9002 6985
rect 8974 6953 9002 6959
rect 8918 6761 8946 6767
rect 8918 6735 8919 6761
rect 8945 6735 8946 6761
rect 8918 6537 8946 6735
rect 8918 6511 8919 6537
rect 8945 6511 8946 6537
rect 8918 6505 8946 6511
rect 8582 6455 8583 6481
rect 8609 6455 8610 6481
rect 8582 6449 8610 6455
rect 9030 6426 9058 7238
rect 9086 6929 9114 7574
rect 9534 7377 9562 7742
rect 9590 7737 9618 7742
rect 9758 7737 9786 7742
rect 9702 7658 9730 7663
rect 9702 7611 9730 7630
rect 9646 7602 9674 7607
rect 9646 7555 9674 7574
rect 9758 7546 9786 7551
rect 9702 7518 9758 7546
rect 9702 7378 9730 7518
rect 9758 7513 9786 7518
rect 9534 7351 9535 7377
rect 9561 7351 9562 7377
rect 9534 7345 9562 7351
rect 9646 7350 9730 7378
rect 9590 7154 9618 7159
rect 9590 7107 9618 7126
rect 9086 6903 9087 6929
rect 9113 6903 9114 6929
rect 9086 6897 9114 6903
rect 9254 6986 9282 6991
rect 9254 6873 9282 6958
rect 9646 6929 9674 7350
rect 9646 6903 9647 6929
rect 9673 6903 9674 6929
rect 9646 6897 9674 6903
rect 9702 7265 9730 7271
rect 9702 7239 9703 7265
rect 9729 7239 9730 7265
rect 9254 6847 9255 6873
rect 9281 6847 9282 6873
rect 9254 6841 9282 6847
rect 8750 6398 9058 6426
rect 8470 5866 8498 5871
rect 8414 5838 8470 5866
rect 8470 5833 8498 5838
rect 2238 5110 2370 5115
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2238 5077 2370 5082
rect 2238 4326 2370 4331
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2238 4293 2370 4298
rect 8750 4214 8778 6398
rect 9702 6370 9730 7239
rect 9758 6986 9786 6991
rect 9814 6986 9842 7910
rect 9918 7854 10050 7859
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 9918 7821 10050 7826
rect 10318 7770 10346 8471
rect 10318 7737 10346 7742
rect 10710 8441 10738 8447
rect 10710 8415 10711 8441
rect 10737 8415 10738 8441
rect 10710 8050 10738 8415
rect 10654 7714 10682 7719
rect 10710 7714 10738 8022
rect 10654 7713 10738 7714
rect 10654 7687 10655 7713
rect 10681 7687 10738 7713
rect 10654 7686 10738 7687
rect 10654 7681 10682 7686
rect 10822 7658 10850 7663
rect 10486 7630 10626 7658
rect 10486 7602 10514 7630
rect 10598 7602 10626 7630
rect 10822 7611 10850 7630
rect 10934 7658 10962 7663
rect 10990 7658 11018 8638
rect 11102 8554 11130 8751
rect 11158 8778 11186 8783
rect 11550 8778 11578 11046
rect 11662 10738 11690 11047
rect 11662 10705 11690 10710
rect 11662 10401 11690 10407
rect 11662 10375 11663 10401
rect 11689 10375 11690 10401
rect 11662 10122 11690 10375
rect 11830 10234 11858 11158
rect 11886 10850 11914 11606
rect 11942 11601 11970 11606
rect 11998 11634 12026 11639
rect 11998 11587 12026 11606
rect 12446 11241 12474 11831
rect 13286 11689 13314 12278
rect 13286 11663 13287 11689
rect 13313 11663 13314 11689
rect 13286 11657 13314 11663
rect 13342 11690 13370 12671
rect 13678 12474 13706 13230
rect 14294 13258 14322 13263
rect 14294 13211 14322 13230
rect 14070 13146 14098 13151
rect 14070 13089 14098 13118
rect 18830 13146 18858 13511
rect 18830 13113 18858 13118
rect 20006 13146 20034 13567
rect 20006 13113 20034 13118
rect 14070 13063 14071 13089
rect 14097 13063 14098 13089
rect 14070 13057 14098 13063
rect 17598 12950 17730 12955
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17598 12917 17730 12922
rect 13454 12473 13874 12474
rect 13454 12447 13679 12473
rect 13705 12447 13874 12473
rect 13454 12446 13874 12447
rect 13454 12025 13482 12446
rect 13454 11999 13455 12025
rect 13481 11999 13482 12025
rect 13454 11993 13482 11999
rect 13566 11858 13594 11863
rect 13342 11657 13370 11662
rect 13454 11830 13566 11858
rect 12894 11634 12922 11639
rect 12894 11577 12922 11606
rect 13398 11633 13426 11639
rect 13398 11607 13399 11633
rect 13425 11607 13426 11633
rect 13118 11578 13146 11583
rect 12894 11551 12895 11577
rect 12921 11551 12922 11577
rect 12894 11545 12922 11551
rect 13062 11577 13146 11578
rect 13062 11551 13119 11577
rect 13145 11551 13146 11577
rect 13062 11550 13146 11551
rect 12446 11215 12447 11241
rect 12473 11215 12474 11241
rect 12446 11209 12474 11215
rect 12110 11185 12138 11191
rect 12110 11159 12111 11185
rect 12137 11159 12138 11185
rect 11998 10906 12026 10911
rect 12110 10906 12138 11159
rect 12026 10878 12082 10906
rect 11998 10873 12026 10878
rect 11886 10822 11970 10850
rect 11662 10089 11690 10094
rect 11718 10206 11914 10234
rect 11718 10094 11746 10206
rect 11718 10066 11802 10094
rect 11606 9729 11634 9735
rect 11606 9703 11607 9729
rect 11633 9703 11634 9729
rect 11606 9282 11634 9703
rect 11774 9506 11802 10066
rect 11886 9673 11914 10206
rect 11942 10094 11970 10822
rect 12054 10793 12082 10878
rect 12110 10873 12138 10878
rect 13062 10905 13090 11550
rect 13118 11545 13146 11550
rect 13062 10879 13063 10905
rect 13089 10879 13090 10905
rect 13062 10850 13090 10879
rect 13062 10817 13090 10822
rect 13286 10849 13314 10855
rect 13286 10823 13287 10849
rect 13313 10823 13314 10849
rect 12054 10767 12055 10793
rect 12081 10767 12082 10793
rect 12054 10761 12082 10767
rect 12334 10794 12362 10799
rect 12334 10747 12362 10766
rect 12726 10794 12754 10799
rect 11942 10066 12138 10094
rect 11886 9647 11887 9673
rect 11913 9647 11914 9673
rect 11886 9641 11914 9647
rect 11718 9478 11802 9506
rect 11830 9617 11858 9623
rect 11830 9591 11831 9617
rect 11857 9591 11858 9617
rect 11662 9282 11690 9287
rect 11606 9254 11662 9282
rect 11606 9170 11634 9175
rect 11606 9123 11634 9142
rect 11662 9058 11690 9254
rect 11718 9225 11746 9478
rect 11830 9394 11858 9591
rect 11830 9337 11858 9366
rect 11830 9311 11831 9337
rect 11857 9311 11858 9337
rect 11830 9305 11858 9311
rect 11998 9506 12026 9511
rect 11718 9199 11719 9225
rect 11745 9199 11746 9225
rect 11718 9193 11746 9199
rect 11942 9225 11970 9231
rect 11942 9199 11943 9225
rect 11969 9199 11970 9225
rect 11158 8777 11578 8778
rect 11158 8751 11159 8777
rect 11185 8751 11578 8777
rect 11158 8750 11578 8751
rect 11606 9030 11690 9058
rect 11886 9114 11914 9119
rect 11158 8745 11186 8750
rect 11102 8521 11130 8526
rect 11270 8497 11298 8750
rect 11270 8471 11271 8497
rect 11297 8471 11298 8497
rect 11270 8465 11298 8471
rect 11326 8610 11354 8615
rect 10934 7657 11018 7658
rect 10934 7631 10935 7657
rect 10961 7631 11018 7657
rect 10934 7630 11018 7631
rect 11046 8441 11074 8447
rect 11046 8415 11047 8441
rect 11073 8415 11074 8441
rect 11046 7994 11074 8415
rect 11326 8441 11354 8582
rect 11326 8415 11327 8441
rect 11353 8415 11354 8441
rect 11326 8409 11354 8415
rect 11438 8386 11466 8391
rect 11438 8339 11466 8358
rect 11046 7658 11074 7966
rect 11438 8274 11466 8279
rect 11214 7770 11242 7775
rect 10934 7625 10962 7630
rect 11046 7625 11074 7630
rect 11102 7742 11214 7770
rect 10710 7602 10738 7607
rect 10598 7601 10738 7602
rect 10598 7575 10711 7601
rect 10737 7575 10738 7601
rect 10598 7574 10738 7575
rect 10486 7569 10514 7574
rect 10710 7569 10738 7574
rect 10542 7546 10570 7551
rect 10934 7546 10962 7551
rect 10542 7545 10682 7546
rect 10542 7519 10543 7545
rect 10569 7519 10682 7545
rect 10542 7518 10682 7519
rect 10542 7513 10570 7518
rect 10654 7434 10682 7518
rect 10654 7406 10794 7434
rect 10766 7377 10794 7406
rect 10766 7351 10767 7377
rect 10793 7351 10794 7377
rect 10766 7345 10794 7351
rect 10934 7265 10962 7518
rect 10934 7239 10935 7265
rect 10961 7239 10962 7265
rect 10934 7233 10962 7239
rect 11102 7265 11130 7742
rect 11214 7723 11242 7742
rect 11438 7769 11466 8246
rect 11438 7743 11439 7769
rect 11465 7743 11466 7769
rect 11438 7737 11466 7743
rect 11326 7657 11354 7663
rect 11326 7631 11327 7657
rect 11353 7631 11354 7657
rect 11326 7602 11354 7631
rect 11326 7569 11354 7574
rect 11382 7601 11410 7607
rect 11382 7575 11383 7601
rect 11409 7575 11410 7601
rect 11326 7378 11354 7383
rect 11382 7378 11410 7575
rect 11326 7377 11410 7378
rect 11326 7351 11327 7377
rect 11353 7351 11410 7377
rect 11326 7350 11410 7351
rect 11326 7345 11354 7350
rect 11102 7239 11103 7265
rect 11129 7239 11130 7265
rect 11102 7233 11130 7239
rect 11494 7266 11522 7271
rect 11606 7266 11634 9030
rect 11718 8554 11746 8559
rect 11718 7769 11746 8526
rect 11830 8330 11858 8335
rect 11718 7743 11719 7769
rect 11745 7743 11746 7769
rect 11718 7737 11746 7743
rect 11774 7993 11802 7999
rect 11774 7967 11775 7993
rect 11801 7967 11802 7993
rect 11774 7769 11802 7967
rect 11774 7743 11775 7769
rect 11801 7743 11802 7769
rect 11774 7737 11802 7743
rect 11830 7658 11858 8302
rect 11886 8049 11914 9086
rect 11942 9058 11970 9199
rect 11942 9025 11970 9030
rect 11886 8023 11887 8049
rect 11913 8023 11914 8049
rect 11886 8017 11914 8023
rect 11998 8049 12026 9478
rect 12110 9505 12138 10066
rect 12726 10009 12754 10766
rect 13230 10793 13258 10799
rect 13230 10767 13231 10793
rect 13257 10767 13258 10793
rect 12782 10738 12810 10743
rect 12782 10691 12810 10710
rect 13118 10738 13146 10743
rect 12726 9983 12727 10009
rect 12753 9983 12754 10009
rect 12726 9977 12754 9983
rect 13118 10009 13146 10710
rect 13118 9983 13119 10009
rect 13145 9983 13146 10009
rect 13118 9977 13146 9983
rect 13062 9953 13090 9959
rect 13062 9927 13063 9953
rect 13089 9927 13090 9953
rect 13062 9898 13090 9927
rect 13230 9898 13258 10767
rect 13286 10794 13314 10823
rect 13286 10761 13314 10766
rect 13062 9870 13258 9898
rect 13286 10681 13314 10687
rect 13398 10682 13426 11607
rect 13454 11633 13482 11830
rect 13566 11825 13594 11830
rect 13454 11607 13455 11633
rect 13481 11607 13482 11633
rect 13454 11601 13482 11607
rect 13622 11578 13650 12446
rect 13678 12441 13706 12446
rect 13846 12361 13874 12446
rect 13846 12335 13847 12361
rect 13873 12335 13874 12361
rect 13846 12329 13874 12335
rect 18830 12362 18858 12367
rect 18830 12315 18858 12334
rect 14238 12306 14266 12311
rect 14238 12259 14266 12278
rect 15302 12306 15330 12311
rect 13958 11970 13986 11975
rect 13958 11923 13986 11942
rect 15302 11970 15330 12278
rect 20006 12249 20034 12255
rect 20006 12223 20007 12249
rect 20033 12223 20034 12249
rect 17598 12166 17730 12171
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17598 12133 17730 12138
rect 20006 12138 20034 12223
rect 20006 12105 20034 12110
rect 20006 12025 20034 12031
rect 20006 11999 20007 12025
rect 20033 11999 20034 12025
rect 15302 11937 15330 11942
rect 18830 11969 18858 11975
rect 18830 11943 18831 11969
rect 18857 11943 18858 11969
rect 13846 11857 13874 11863
rect 13846 11831 13847 11857
rect 13873 11831 13874 11857
rect 13846 11634 13874 11831
rect 13902 11858 13930 11863
rect 13902 11811 13930 11830
rect 14070 11857 14098 11863
rect 14070 11831 14071 11857
rect 14097 11831 14098 11857
rect 13846 11601 13874 11606
rect 14070 11690 14098 11831
rect 18830 11746 18858 11943
rect 20006 11802 20034 11999
rect 20006 11769 20034 11774
rect 18830 11713 18858 11718
rect 13622 11577 13762 11578
rect 13622 11551 13623 11577
rect 13649 11551 13762 11577
rect 13622 11550 13762 11551
rect 13622 11545 13650 11550
rect 13510 11242 13538 11247
rect 13510 11241 13594 11242
rect 13510 11215 13511 11241
rect 13537 11215 13594 11241
rect 13510 11214 13594 11215
rect 13510 11209 13538 11214
rect 13566 11074 13594 11214
rect 13678 11130 13706 11135
rect 13510 10850 13538 10855
rect 13510 10803 13538 10822
rect 13566 10849 13594 11046
rect 13566 10823 13567 10849
rect 13593 10823 13594 10849
rect 13566 10817 13594 10823
rect 13622 11129 13706 11130
rect 13622 11103 13679 11129
rect 13705 11103 13706 11129
rect 13622 11102 13706 11103
rect 13286 10655 13287 10681
rect 13313 10655 13314 10681
rect 13062 9786 13090 9870
rect 13062 9753 13090 9758
rect 13286 9730 13314 10655
rect 13286 9683 13314 9702
rect 13342 10654 13426 10682
rect 13342 10402 13370 10654
rect 12110 9479 12111 9505
rect 12137 9479 12138 9505
rect 12110 8330 12138 9479
rect 12222 9617 12250 9623
rect 12222 9591 12223 9617
rect 12249 9591 12250 9617
rect 12222 9394 12250 9591
rect 12950 9618 12978 9623
rect 12950 9571 12978 9590
rect 13174 9618 13202 9623
rect 13174 9571 13202 9590
rect 13342 9562 13370 10374
rect 13510 10458 13538 10463
rect 13398 10066 13426 10071
rect 13398 10019 13426 10038
rect 13454 9618 13482 9637
rect 13454 9585 13482 9590
rect 13342 9529 13370 9534
rect 12838 9506 12866 9511
rect 12838 9459 12866 9478
rect 13454 9506 13482 9511
rect 12222 9361 12250 9366
rect 13454 9282 13482 9478
rect 12502 9170 12530 9175
rect 12502 8889 12530 9142
rect 12502 8863 12503 8889
rect 12529 8863 12530 8889
rect 12502 8857 12530 8863
rect 12894 8833 12922 8839
rect 12894 8807 12895 8833
rect 12921 8807 12922 8833
rect 12894 8722 12922 8807
rect 13454 8834 13482 9254
rect 13510 9170 13538 10430
rect 13622 10094 13650 11102
rect 13678 11097 13706 11102
rect 13734 10906 13762 11550
rect 14014 11522 14042 11527
rect 13902 11521 14042 11522
rect 13902 11495 14015 11521
rect 14041 11495 14042 11521
rect 13902 11494 14042 11495
rect 13902 11241 13930 11494
rect 14014 11489 14042 11494
rect 14070 11298 14098 11662
rect 15414 11634 15442 11639
rect 15414 11587 15442 11606
rect 15246 11578 15274 11583
rect 15078 11522 15106 11527
rect 15246 11522 15274 11550
rect 18830 11578 18858 11583
rect 18830 11531 18858 11550
rect 15078 11521 15274 11522
rect 15078 11495 15079 11521
rect 15105 11495 15274 11521
rect 15078 11494 15274 11495
rect 13902 11215 13903 11241
rect 13929 11215 13930 11241
rect 13902 11209 13930 11215
rect 13958 11270 14098 11298
rect 14182 11298 14210 11303
rect 14182 11297 14266 11298
rect 14182 11271 14183 11297
rect 14209 11271 14266 11297
rect 14182 11270 14266 11271
rect 13790 11186 13818 11191
rect 13790 11139 13818 11158
rect 13958 11074 13986 11270
rect 14182 11265 14210 11270
rect 14014 11186 14042 11191
rect 14014 11139 14042 11158
rect 14238 11186 14266 11270
rect 14238 11153 14266 11158
rect 14126 11129 14154 11135
rect 14126 11103 14127 11129
rect 14153 11103 14154 11129
rect 14126 11074 14154 11103
rect 14182 11130 14210 11135
rect 14182 11083 14210 11102
rect 15078 11130 15106 11494
rect 20006 11466 20034 11471
rect 20006 11419 20034 11438
rect 17598 11382 17730 11387
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17598 11349 17730 11354
rect 15078 11097 15106 11102
rect 13958 11046 14154 11074
rect 13790 10906 13818 10911
rect 14014 10906 14042 10911
rect 13762 10905 14042 10906
rect 13762 10879 13791 10905
rect 13817 10879 14015 10905
rect 14041 10879 14042 10905
rect 13762 10878 14042 10879
rect 13734 10458 13762 10878
rect 13790 10873 13818 10878
rect 13734 10411 13762 10430
rect 13566 10066 13650 10094
rect 13790 10066 13818 10071
rect 13566 9506 13594 10066
rect 13678 10065 13818 10066
rect 13678 10039 13791 10065
rect 13817 10039 13818 10065
rect 13678 10038 13818 10039
rect 13622 9730 13650 9735
rect 13622 9617 13650 9702
rect 13678 9729 13706 10038
rect 13790 10033 13818 10038
rect 13846 10010 13874 10015
rect 13846 10009 13986 10010
rect 13846 9983 13847 10009
rect 13873 9983 13986 10009
rect 13846 9982 13986 9983
rect 13846 9977 13874 9982
rect 13790 9898 13818 9903
rect 13790 9897 13930 9898
rect 13790 9871 13791 9897
rect 13817 9871 13930 9897
rect 13790 9870 13930 9871
rect 13790 9865 13818 9870
rect 13678 9703 13679 9729
rect 13705 9703 13706 9729
rect 13678 9697 13706 9703
rect 13622 9591 13623 9617
rect 13649 9591 13650 9617
rect 13622 9585 13650 9591
rect 13678 9506 13706 9511
rect 13566 9505 13706 9506
rect 13566 9479 13679 9505
rect 13705 9479 13706 9505
rect 13566 9478 13706 9479
rect 13678 9450 13706 9478
rect 13678 9417 13706 9422
rect 13902 9394 13930 9870
rect 13958 9730 13986 9982
rect 14014 10009 14042 10878
rect 17598 10598 17730 10603
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17598 10565 17730 10570
rect 14294 10066 14322 10071
rect 14322 10038 14378 10066
rect 14294 10033 14322 10038
rect 14014 9983 14015 10009
rect 14041 9983 14042 10009
rect 14014 9977 14042 9983
rect 13958 9702 14154 9730
rect 14126 9673 14154 9702
rect 14126 9647 14127 9673
rect 14153 9647 14154 9673
rect 14126 9641 14154 9647
rect 13958 9561 13986 9567
rect 13958 9535 13959 9561
rect 13985 9535 13986 9561
rect 13958 9506 13986 9535
rect 14070 9562 14098 9567
rect 14070 9515 14098 9534
rect 14182 9562 14210 9567
rect 14182 9515 14210 9534
rect 13958 9473 13986 9478
rect 14238 9506 14266 9511
rect 14350 9506 14378 10038
rect 15302 10010 15330 10015
rect 14406 9954 14434 9959
rect 14406 9953 14826 9954
rect 14406 9927 14407 9953
rect 14433 9927 14826 9953
rect 14406 9926 14826 9927
rect 14406 9921 14434 9926
rect 14798 9673 14826 9926
rect 15078 9729 15106 9735
rect 15078 9703 15079 9729
rect 15105 9703 15106 9729
rect 15078 9674 15106 9703
rect 14798 9647 14799 9673
rect 14825 9647 14826 9673
rect 14798 9641 14826 9647
rect 14966 9646 15106 9674
rect 14238 9505 14378 9506
rect 14238 9479 14239 9505
rect 14265 9479 14378 9505
rect 14238 9478 14378 9479
rect 14238 9473 14266 9478
rect 14350 9450 14378 9478
rect 13902 9366 14266 9394
rect 14182 9282 14210 9287
rect 13846 9225 13874 9231
rect 13846 9199 13847 9225
rect 13873 9199 13874 9225
rect 13678 9170 13706 9175
rect 13846 9170 13874 9199
rect 13510 9169 13874 9170
rect 13510 9143 13679 9169
rect 13705 9143 13874 9169
rect 13510 9142 13874 9143
rect 13454 8806 13650 8834
rect 12894 8689 12922 8694
rect 13118 8722 13146 8727
rect 13118 8675 13146 8694
rect 13454 8722 13482 8727
rect 12110 8297 12138 8302
rect 11998 8023 11999 8049
rect 12025 8023 12026 8049
rect 11830 7611 11858 7630
rect 11886 7937 11914 7943
rect 11886 7911 11887 7937
rect 11913 7911 11914 7937
rect 11886 7322 11914 7911
rect 11998 7714 12026 8023
rect 11998 7681 12026 7686
rect 13454 7770 13482 8694
rect 13622 8050 13650 8806
rect 13678 8722 13706 9142
rect 13678 8689 13706 8694
rect 14182 8554 14210 9254
rect 14238 9281 14266 9366
rect 14238 9255 14239 9281
rect 14265 9255 14266 9281
rect 14238 9249 14266 9255
rect 14014 8526 14210 8554
rect 13846 8441 13874 8447
rect 13846 8415 13847 8441
rect 13873 8415 13874 8441
rect 13846 8386 13874 8415
rect 13678 8050 13706 8055
rect 13622 8049 13706 8050
rect 13622 8023 13679 8049
rect 13705 8023 13706 8049
rect 13622 8022 13706 8023
rect 13678 8017 13706 8022
rect 13846 8049 13874 8358
rect 13958 8385 13986 8391
rect 13958 8359 13959 8385
rect 13985 8359 13986 8385
rect 13958 8162 13986 8359
rect 13846 8023 13847 8049
rect 13873 8023 13874 8049
rect 13846 8017 13874 8023
rect 13902 8134 13986 8162
rect 12054 7658 12082 7663
rect 12054 7611 12082 7630
rect 13118 7658 13146 7663
rect 12334 7602 12362 7607
rect 12054 7322 12082 7327
rect 11886 7321 12082 7322
rect 11886 7295 12055 7321
rect 12081 7295 12082 7321
rect 11886 7294 12082 7295
rect 12054 7289 12082 7294
rect 11494 7265 11634 7266
rect 11494 7239 11495 7265
rect 11521 7239 11634 7265
rect 11494 7238 11634 7239
rect 11662 7265 11690 7271
rect 11662 7239 11663 7265
rect 11689 7239 11690 7265
rect 11494 7233 11522 7238
rect 10822 7153 10850 7159
rect 11382 7154 11410 7159
rect 10822 7127 10823 7153
rect 10849 7127 10850 7153
rect 9918 7070 10050 7075
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 9918 7037 10050 7042
rect 9786 6958 9842 6986
rect 9758 6953 9786 6958
rect 10206 6818 10234 6823
rect 9982 6537 10010 6543
rect 9982 6511 9983 6537
rect 10009 6511 10010 6537
rect 9982 6370 10010 6511
rect 10206 6537 10234 6790
rect 10206 6511 10207 6537
rect 10233 6511 10234 6537
rect 10206 6505 10234 6511
rect 10710 6818 10738 6823
rect 10822 6818 10850 7127
rect 11270 7153 11410 7154
rect 11270 7127 11383 7153
rect 11409 7127 11410 7153
rect 11270 7126 11410 7127
rect 11270 6929 11298 7126
rect 11382 7121 11410 7126
rect 11270 6903 11271 6929
rect 11297 6903 11298 6929
rect 11270 6897 11298 6903
rect 10934 6874 10962 6879
rect 10934 6827 10962 6846
rect 11662 6874 11690 7239
rect 11662 6841 11690 6846
rect 10710 6817 10850 6818
rect 10710 6791 10711 6817
rect 10737 6791 10850 6817
rect 10710 6790 10850 6791
rect 12334 6817 12362 7574
rect 13118 7321 13146 7630
rect 13118 7295 13119 7321
rect 13145 7295 13146 7321
rect 12670 6874 12698 6879
rect 12670 6827 12698 6846
rect 12334 6791 12335 6817
rect 12361 6791 12362 6817
rect 9702 6342 10010 6370
rect 8862 5866 8890 5871
rect 8750 4186 8834 4214
rect 2238 3542 2370 3547
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2238 3509 2370 3514
rect 2238 2758 2370 2763
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2238 2725 2370 2730
rect 8750 2618 8778 2623
rect 2238 1974 2370 1979
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2238 1941 2370 1946
rect 8750 400 8778 2590
rect 8806 1777 8834 4186
rect 8862 2561 8890 5838
rect 9366 2618 9394 2623
rect 9366 2571 9394 2590
rect 8862 2535 8863 2561
rect 8889 2535 8890 2561
rect 8862 2529 8890 2535
rect 9814 2170 9842 6342
rect 9918 6286 10050 6291
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 9918 6253 10050 6258
rect 9918 5502 10050 5507
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 9918 5469 10050 5474
rect 9918 4718 10050 4723
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 9918 4685 10050 4690
rect 9918 3934 10050 3939
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 9918 3901 10050 3906
rect 9918 3150 10050 3155
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 9918 3117 10050 3122
rect 9918 2366 10050 2371
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 9918 2333 10050 2338
rect 9870 2170 9898 2175
rect 9814 2169 9898 2170
rect 9814 2143 9871 2169
rect 9897 2143 9898 2169
rect 9814 2142 9898 2143
rect 9870 2137 9898 2142
rect 9758 2058 9786 2063
rect 9310 1834 9338 1839
rect 8806 1751 8807 1777
rect 8833 1751 8834 1777
rect 8806 1745 8834 1751
rect 9086 1833 9338 1834
rect 9086 1807 9311 1833
rect 9337 1807 9338 1833
rect 9086 1806 9338 1807
rect 9086 400 9114 1806
rect 9310 1801 9338 1806
rect 9758 400 9786 2030
rect 10374 2058 10402 2063
rect 10374 2011 10402 2030
rect 10710 1777 10738 6790
rect 12334 4214 12362 6791
rect 13118 4214 13146 7295
rect 13454 7657 13482 7742
rect 13846 7714 13874 7719
rect 13902 7714 13930 8134
rect 13958 8050 13986 8055
rect 14014 8050 14042 8526
rect 14182 8497 14210 8526
rect 14182 8471 14183 8497
rect 14209 8471 14210 8497
rect 14182 8465 14210 8471
rect 14070 8441 14098 8447
rect 14070 8415 14071 8441
rect 14097 8415 14098 8441
rect 14070 8162 14098 8415
rect 14350 8162 14378 9422
rect 14574 9618 14602 9623
rect 14574 9282 14602 9590
rect 14910 9618 14938 9623
rect 14966 9618 14994 9646
rect 14910 9617 14994 9618
rect 14910 9591 14911 9617
rect 14937 9591 14994 9617
rect 14910 9590 14994 9591
rect 14910 9585 14938 9590
rect 14686 9561 14714 9567
rect 14686 9535 14687 9561
rect 14713 9535 14714 9561
rect 14686 9506 14714 9535
rect 14686 9473 14714 9478
rect 15022 9561 15050 9567
rect 15022 9535 15023 9561
rect 15049 9535 15050 9561
rect 15022 9450 15050 9535
rect 15302 9562 15330 9982
rect 18830 10010 18858 10015
rect 18830 9963 18858 9982
rect 15078 9506 15106 9511
rect 15078 9459 15106 9478
rect 15022 9417 15050 9422
rect 14574 9249 14602 9254
rect 15302 9169 15330 9534
rect 15470 9953 15498 9959
rect 15470 9927 15471 9953
rect 15497 9927 15498 9953
rect 15470 9506 15498 9927
rect 20006 9897 20034 9903
rect 20006 9871 20007 9897
rect 20033 9871 20034 9897
rect 17598 9814 17730 9819
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17598 9781 17730 9786
rect 20006 9786 20034 9871
rect 20006 9753 20034 9758
rect 20006 9673 20034 9679
rect 20006 9647 20007 9673
rect 20033 9647 20034 9673
rect 18830 9618 18858 9623
rect 18830 9571 18858 9590
rect 15470 9473 15498 9478
rect 20006 9450 20034 9647
rect 20006 9417 20034 9422
rect 15302 9143 15303 9169
rect 15329 9143 15330 9169
rect 15302 9137 15330 9143
rect 17598 9030 17730 9035
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17598 8997 17730 9002
rect 18942 8441 18970 8447
rect 18942 8415 18943 8441
rect 18969 8415 18970 8441
rect 17598 8246 17730 8251
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17598 8213 17730 8218
rect 14070 8129 14098 8134
rect 14126 8134 14378 8162
rect 13958 8049 14042 8050
rect 13958 8023 13959 8049
rect 13985 8023 14042 8049
rect 13958 8022 14042 8023
rect 14070 8050 14098 8055
rect 14126 8050 14154 8134
rect 14070 8049 14154 8050
rect 14070 8023 14071 8049
rect 14097 8023 14154 8049
rect 14070 8022 14154 8023
rect 14350 8050 14378 8134
rect 13958 8017 13986 8022
rect 14070 8017 14098 8022
rect 14350 8017 14378 8022
rect 14518 8162 14546 8167
rect 14518 8049 14546 8134
rect 14518 8023 14519 8049
rect 14545 8023 14546 8049
rect 14518 8017 14546 8023
rect 14686 8050 14714 8055
rect 14686 8003 14714 8022
rect 14910 8050 14938 8055
rect 14910 8003 14938 8022
rect 15134 8050 15162 8055
rect 18830 8050 18858 8055
rect 15162 8022 15218 8050
rect 15134 8017 15162 8022
rect 14182 7994 14210 7999
rect 14182 7947 14210 7966
rect 14854 7994 14882 7999
rect 14854 7947 14882 7966
rect 13846 7713 13930 7714
rect 13846 7687 13847 7713
rect 13873 7687 13930 7713
rect 13846 7686 13930 7687
rect 14126 7937 14154 7943
rect 14126 7911 14127 7937
rect 14153 7911 14154 7937
rect 13846 7681 13874 7686
rect 13454 7631 13455 7657
rect 13481 7631 13482 7657
rect 13342 7153 13370 7159
rect 13342 7127 13343 7153
rect 13369 7127 13370 7153
rect 13342 6986 13370 7127
rect 13454 6986 13482 7631
rect 13510 6986 13538 6991
rect 13342 6985 13706 6986
rect 13342 6959 13511 6985
rect 13537 6959 13706 6985
rect 13342 6958 13706 6959
rect 13342 6874 13370 6958
rect 13510 6953 13538 6958
rect 13342 6841 13370 6846
rect 13678 6873 13706 6958
rect 14070 6930 14098 6935
rect 14126 6930 14154 7911
rect 14630 7938 14658 7943
rect 14630 7891 14658 7910
rect 14966 7938 14994 7943
rect 14910 7602 14938 7607
rect 14966 7602 14994 7910
rect 15134 7770 15162 7775
rect 15134 7723 15162 7742
rect 14910 7601 14994 7602
rect 14910 7575 14911 7601
rect 14937 7575 14994 7601
rect 14910 7574 14994 7575
rect 14910 7569 14938 7574
rect 14070 6929 14154 6930
rect 14070 6903 14071 6929
rect 14097 6903 14154 6929
rect 14070 6902 14154 6903
rect 14070 6897 14098 6902
rect 13678 6847 13679 6873
rect 13705 6847 13706 6873
rect 13678 6841 13706 6847
rect 15134 6818 15162 6823
rect 15190 6818 15218 8022
rect 18830 8003 18858 8022
rect 18942 7938 18970 8415
rect 19950 8385 19978 8391
rect 19950 8359 19951 8385
rect 19977 8359 19978 8385
rect 19950 8106 19978 8359
rect 19950 8073 19978 8078
rect 20006 8105 20034 8111
rect 20006 8079 20007 8105
rect 20033 8079 20034 8105
rect 18942 7905 18970 7910
rect 20006 7770 20034 8079
rect 20006 7737 20034 7742
rect 17598 7462 17730 7467
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17598 7429 17730 7434
rect 15134 6817 15218 6818
rect 15134 6791 15135 6817
rect 15161 6791 15218 6817
rect 15134 6790 15218 6791
rect 15134 6785 15162 6790
rect 17598 6678 17730 6683
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17598 6645 17730 6650
rect 17598 5894 17730 5899
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17598 5861 17730 5866
rect 17598 5110 17730 5115
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17598 5077 17730 5082
rect 17598 4326 17730 4331
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17598 4293 17730 4298
rect 12278 4186 12362 4214
rect 12614 4186 13146 4214
rect 12110 2058 12138 2063
rect 10710 1751 10711 1777
rect 10737 1751 10738 1777
rect 10710 1745 10738 1751
rect 11438 1834 11466 1839
rect 11214 1666 11242 1671
rect 11102 1665 11242 1666
rect 11102 1639 11215 1665
rect 11241 1639 11242 1665
rect 11102 1638 11242 1639
rect 9918 1582 10050 1587
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 9918 1549 10050 1554
rect 11102 400 11130 1638
rect 11214 1633 11242 1638
rect 11438 400 11466 1806
rect 12110 400 12138 2030
rect 12278 1777 12306 4186
rect 12614 2169 12642 4186
rect 17598 3542 17730 3547
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17598 3509 17730 3514
rect 17598 2758 17730 2763
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17598 2725 17730 2730
rect 12614 2143 12615 2169
rect 12641 2143 12642 2169
rect 12614 2137 12642 2143
rect 13118 2058 13146 2063
rect 13118 2011 13146 2030
rect 17598 1974 17730 1979
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17598 1941 17730 1946
rect 12782 1834 12810 1839
rect 12782 1787 12810 1806
rect 12278 1751 12279 1777
rect 12305 1751 12306 1777
rect 12278 1745 12306 1751
rect 8736 0 8792 400
rect 9072 0 9128 400
rect 9744 0 9800 400
rect 11088 0 11144 400
rect 11424 0 11480 400
rect 12096 0 12152 400
<< via2 >>
rect 2238 19221 2266 19222
rect 2238 19195 2239 19221
rect 2239 19195 2265 19221
rect 2265 19195 2266 19221
rect 2238 19194 2266 19195
rect 2290 19221 2318 19222
rect 2290 19195 2291 19221
rect 2291 19195 2317 19221
rect 2317 19195 2318 19221
rect 2290 19194 2318 19195
rect 2342 19221 2370 19222
rect 2342 19195 2343 19221
rect 2343 19195 2369 19221
rect 2369 19195 2370 19221
rect 2342 19194 2370 19195
rect 2238 18437 2266 18438
rect 2238 18411 2239 18437
rect 2239 18411 2265 18437
rect 2265 18411 2266 18437
rect 2238 18410 2266 18411
rect 2290 18437 2318 18438
rect 2290 18411 2291 18437
rect 2291 18411 2317 18437
rect 2317 18411 2318 18437
rect 2290 18410 2318 18411
rect 2342 18437 2370 18438
rect 2342 18411 2343 18437
rect 2343 18411 2369 18437
rect 2369 18411 2370 18437
rect 2342 18410 2370 18411
rect 8750 19110 8778 19138
rect 9310 19137 9338 19138
rect 9310 19111 9311 19137
rect 9311 19111 9337 19137
rect 9337 19111 9338 19137
rect 9310 19110 9338 19111
rect 7742 18326 7770 18354
rect 8358 18353 8386 18354
rect 8358 18327 8359 18353
rect 8359 18327 8385 18353
rect 8385 18327 8386 18353
rect 8358 18326 8386 18327
rect 2238 17653 2266 17654
rect 2238 17627 2239 17653
rect 2239 17627 2265 17653
rect 2265 17627 2266 17653
rect 2238 17626 2266 17627
rect 2290 17653 2318 17654
rect 2290 17627 2291 17653
rect 2291 17627 2317 17653
rect 2317 17627 2318 17653
rect 2290 17626 2318 17627
rect 2342 17653 2370 17654
rect 2342 17627 2343 17653
rect 2343 17627 2369 17653
rect 2369 17627 2370 17653
rect 2342 17626 2370 17627
rect 2238 16869 2266 16870
rect 2238 16843 2239 16869
rect 2239 16843 2265 16869
rect 2265 16843 2266 16869
rect 2238 16842 2266 16843
rect 2290 16869 2318 16870
rect 2290 16843 2291 16869
rect 2291 16843 2317 16869
rect 2317 16843 2318 16869
rect 2290 16842 2318 16843
rect 2342 16869 2370 16870
rect 2342 16843 2343 16869
rect 2343 16843 2369 16869
rect 2369 16843 2370 16869
rect 2342 16842 2370 16843
rect 2238 16085 2266 16086
rect 2238 16059 2239 16085
rect 2239 16059 2265 16085
rect 2265 16059 2266 16085
rect 2238 16058 2266 16059
rect 2290 16085 2318 16086
rect 2290 16059 2291 16085
rect 2291 16059 2317 16085
rect 2317 16059 2318 16085
rect 2290 16058 2318 16059
rect 2342 16085 2370 16086
rect 2342 16059 2343 16085
rect 2343 16059 2369 16085
rect 2369 16059 2370 16085
rect 2342 16058 2370 16059
rect 2238 15301 2266 15302
rect 2238 15275 2239 15301
rect 2239 15275 2265 15301
rect 2265 15275 2266 15301
rect 2238 15274 2266 15275
rect 2290 15301 2318 15302
rect 2290 15275 2291 15301
rect 2291 15275 2317 15301
rect 2317 15275 2318 15301
rect 2290 15274 2318 15275
rect 2342 15301 2370 15302
rect 2342 15275 2343 15301
rect 2343 15275 2369 15301
rect 2369 15275 2370 15301
rect 2342 15274 2370 15275
rect 2238 14517 2266 14518
rect 2238 14491 2239 14517
rect 2239 14491 2265 14517
rect 2265 14491 2266 14517
rect 2238 14490 2266 14491
rect 2290 14517 2318 14518
rect 2290 14491 2291 14517
rect 2291 14491 2317 14517
rect 2317 14491 2318 14517
rect 2290 14490 2318 14491
rect 2342 14517 2370 14518
rect 2342 14491 2343 14517
rect 2343 14491 2369 14517
rect 2369 14491 2370 14517
rect 2342 14490 2370 14491
rect 2086 13790 2114 13818
rect 966 12782 994 12810
rect 966 11774 994 11802
rect 966 11465 994 11466
rect 966 11439 967 11465
rect 967 11439 993 11465
rect 993 11439 994 11465
rect 966 11438 994 11439
rect 2238 13733 2266 13734
rect 2238 13707 2239 13733
rect 2239 13707 2265 13733
rect 2265 13707 2266 13733
rect 2238 13706 2266 13707
rect 2290 13733 2318 13734
rect 2290 13707 2291 13733
rect 2291 13707 2317 13733
rect 2317 13707 2318 13733
rect 2290 13706 2318 13707
rect 2342 13733 2370 13734
rect 2342 13707 2343 13733
rect 2343 13707 2369 13733
rect 2369 13707 2370 13733
rect 2342 13706 2370 13707
rect 6566 13873 6594 13874
rect 6566 13847 6567 13873
rect 6567 13847 6593 13873
rect 6593 13847 6594 13873
rect 6566 13846 6594 13847
rect 7126 13846 7154 13874
rect 6230 13510 6258 13538
rect 7462 13537 7490 13538
rect 7462 13511 7463 13537
rect 7463 13511 7489 13537
rect 7489 13511 7490 13537
rect 7462 13510 7490 13511
rect 5614 13398 5642 13426
rect 7182 13174 7210 13202
rect 2142 13062 2170 13090
rect 2238 12949 2266 12950
rect 2238 12923 2239 12949
rect 2239 12923 2265 12949
rect 2265 12923 2266 12949
rect 2238 12922 2266 12923
rect 2290 12949 2318 12950
rect 2290 12923 2291 12949
rect 2291 12923 2317 12949
rect 2317 12923 2318 12949
rect 2290 12922 2318 12923
rect 2342 12949 2370 12950
rect 2342 12923 2343 12949
rect 2343 12923 2369 12949
rect 2369 12923 2370 12949
rect 2342 12922 2370 12923
rect 7014 13089 7042 13090
rect 7014 13063 7015 13089
rect 7015 13063 7041 13089
rect 7041 13063 7042 13089
rect 7014 13062 7042 13063
rect 7910 13510 7938 13538
rect 12782 19278 12810 19306
rect 11438 19110 11466 19138
rect 12782 19137 12810 19138
rect 12782 19111 12783 19137
rect 12783 19111 12809 19137
rect 12809 19111 12810 19137
rect 12782 19110 12810 19111
rect 13118 19110 13146 19138
rect 13398 19278 13426 19306
rect 9918 18829 9946 18830
rect 9918 18803 9919 18829
rect 9919 18803 9945 18829
rect 9945 18803 9946 18829
rect 9918 18802 9946 18803
rect 9970 18829 9998 18830
rect 9970 18803 9971 18829
rect 9971 18803 9997 18829
rect 9997 18803 9998 18829
rect 9970 18802 9998 18803
rect 10022 18829 10050 18830
rect 10022 18803 10023 18829
rect 10023 18803 10049 18829
rect 10049 18803 10050 18829
rect 10022 18802 10050 18803
rect 9422 18718 9450 18746
rect 10038 18745 10066 18746
rect 10038 18719 10039 18745
rect 10039 18719 10065 18745
rect 10065 18719 10066 18745
rect 10038 18718 10066 18719
rect 9918 18045 9946 18046
rect 9918 18019 9919 18045
rect 9919 18019 9945 18045
rect 9945 18019 9946 18045
rect 9918 18018 9946 18019
rect 9970 18045 9998 18046
rect 9970 18019 9971 18045
rect 9971 18019 9997 18045
rect 9997 18019 9998 18045
rect 9970 18018 9998 18019
rect 10022 18045 10050 18046
rect 10022 18019 10023 18045
rect 10023 18019 10049 18045
rect 10049 18019 10050 18045
rect 10022 18018 10050 18019
rect 9918 17261 9946 17262
rect 9918 17235 9919 17261
rect 9919 17235 9945 17261
rect 9945 17235 9946 17261
rect 9918 17234 9946 17235
rect 9970 17261 9998 17262
rect 9970 17235 9971 17261
rect 9971 17235 9997 17261
rect 9997 17235 9998 17261
rect 9970 17234 9998 17235
rect 10022 17261 10050 17262
rect 10022 17235 10023 17261
rect 10023 17235 10049 17261
rect 10049 17235 10050 17261
rect 10022 17234 10050 17235
rect 9918 16477 9946 16478
rect 9918 16451 9919 16477
rect 9919 16451 9945 16477
rect 9945 16451 9946 16477
rect 9918 16450 9946 16451
rect 9970 16477 9998 16478
rect 9970 16451 9971 16477
rect 9971 16451 9997 16477
rect 9997 16451 9998 16477
rect 9970 16450 9998 16451
rect 10022 16477 10050 16478
rect 10022 16451 10023 16477
rect 10023 16451 10049 16477
rect 10049 16451 10050 16477
rect 10022 16450 10050 16451
rect 8190 13566 8218 13594
rect 7798 13062 7826 13090
rect 6398 12697 6426 12698
rect 6398 12671 6399 12697
rect 6399 12671 6425 12697
rect 6425 12671 6426 12697
rect 6398 12670 6426 12671
rect 7574 13006 7602 13034
rect 7518 12950 7546 12978
rect 7294 12697 7322 12698
rect 7294 12671 7295 12697
rect 7295 12671 7321 12697
rect 7321 12671 7322 12697
rect 7294 12670 7322 12671
rect 7238 12614 7266 12642
rect 7462 12446 7490 12474
rect 7742 12950 7770 12978
rect 8078 13201 8106 13202
rect 8078 13175 8079 13201
rect 8079 13175 8105 13201
rect 8105 13175 8106 13201
rect 8078 13174 8106 13175
rect 7910 13062 7938 13090
rect 7574 12473 7602 12474
rect 7574 12447 7575 12473
rect 7575 12447 7601 12473
rect 7601 12447 7602 12473
rect 7574 12446 7602 12447
rect 7686 12614 7714 12642
rect 2238 12165 2266 12166
rect 2238 12139 2239 12165
rect 2239 12139 2265 12165
rect 2265 12139 2266 12165
rect 2238 12138 2266 12139
rect 2290 12165 2318 12166
rect 2290 12139 2291 12165
rect 2291 12139 2317 12165
rect 2317 12139 2318 12165
rect 2290 12138 2318 12139
rect 2342 12165 2370 12166
rect 2342 12139 2343 12165
rect 2343 12139 2369 12165
rect 2369 12139 2370 12165
rect 2342 12138 2370 12139
rect 2142 11969 2170 11970
rect 2142 11943 2143 11969
rect 2143 11943 2169 11969
rect 2169 11943 2170 11969
rect 2142 11942 2170 11943
rect 5558 11942 5586 11970
rect 2142 11577 2170 11578
rect 2142 11551 2143 11577
rect 2143 11551 2169 11577
rect 2169 11551 2170 11577
rect 2142 11550 2170 11551
rect 2238 11381 2266 11382
rect 2238 11355 2239 11381
rect 2239 11355 2265 11381
rect 2265 11355 2266 11381
rect 2238 11354 2266 11355
rect 2290 11381 2318 11382
rect 2290 11355 2291 11381
rect 2291 11355 2317 11381
rect 2317 11355 2318 11381
rect 2290 11354 2318 11355
rect 2342 11381 2370 11382
rect 2342 11355 2343 11381
rect 2343 11355 2369 11381
rect 2369 11355 2370 11381
rect 2342 11354 2370 11355
rect 6062 11550 6090 11578
rect 7014 11942 7042 11970
rect 6958 11326 6986 11354
rect 7518 11129 7546 11130
rect 7518 11103 7519 11129
rect 7519 11103 7545 11129
rect 7545 11103 7546 11129
rect 7518 11102 7546 11103
rect 7070 11073 7098 11074
rect 7070 11047 7071 11073
rect 7071 11047 7097 11073
rect 7097 11047 7098 11073
rect 7070 11046 7098 11047
rect 7798 11577 7826 11578
rect 7798 11551 7799 11577
rect 7799 11551 7825 11577
rect 7825 11551 7826 11577
rect 7798 11550 7826 11551
rect 7686 11438 7714 11466
rect 7854 11214 7882 11242
rect 8414 13145 8442 13146
rect 8414 13119 8415 13145
rect 8415 13119 8441 13145
rect 8441 13119 8442 13145
rect 8414 13118 8442 13119
rect 9198 13566 9226 13594
rect 9918 15693 9946 15694
rect 9918 15667 9919 15693
rect 9919 15667 9945 15693
rect 9945 15667 9946 15693
rect 9918 15666 9946 15667
rect 9970 15693 9998 15694
rect 9970 15667 9971 15693
rect 9971 15667 9997 15693
rect 9997 15667 9998 15693
rect 9970 15666 9998 15667
rect 10022 15693 10050 15694
rect 10022 15667 10023 15693
rect 10023 15667 10049 15693
rect 10049 15667 10050 15693
rect 10022 15666 10050 15667
rect 9918 14909 9946 14910
rect 9918 14883 9919 14909
rect 9919 14883 9945 14909
rect 9945 14883 9946 14909
rect 9918 14882 9946 14883
rect 9970 14909 9998 14910
rect 9970 14883 9971 14909
rect 9971 14883 9997 14909
rect 9997 14883 9998 14909
rect 9970 14882 9998 14883
rect 10022 14909 10050 14910
rect 10022 14883 10023 14909
rect 10023 14883 10049 14909
rect 10049 14883 10050 14909
rect 10022 14882 10050 14883
rect 10934 14238 10962 14266
rect 9918 14125 9946 14126
rect 9918 14099 9919 14125
rect 9919 14099 9945 14125
rect 9945 14099 9946 14125
rect 9918 14098 9946 14099
rect 9970 14125 9998 14126
rect 9970 14099 9971 14125
rect 9971 14099 9997 14125
rect 9997 14099 9998 14125
rect 9970 14098 9998 14099
rect 10022 14125 10050 14126
rect 10022 14099 10023 14125
rect 10023 14099 10049 14125
rect 10049 14099 10050 14125
rect 10022 14098 10050 14099
rect 11830 14238 11858 14266
rect 10262 13929 10290 13930
rect 10262 13903 10263 13929
rect 10263 13903 10289 13929
rect 10289 13903 10290 13929
rect 10262 13902 10290 13903
rect 8582 13062 8610 13090
rect 8246 12614 8274 12642
rect 8918 13062 8946 13090
rect 8750 12950 8778 12978
rect 8638 12697 8666 12698
rect 8638 12671 8639 12697
rect 8639 12671 8665 12697
rect 8665 12671 8666 12697
rect 8638 12670 8666 12671
rect 9086 13145 9114 13146
rect 9086 13119 9087 13145
rect 9087 13119 9113 13145
rect 9113 13119 9114 13145
rect 9086 13118 9114 13119
rect 9030 12838 9058 12866
rect 9030 12670 9058 12698
rect 7630 11046 7658 11074
rect 2238 10597 2266 10598
rect 2238 10571 2239 10597
rect 2239 10571 2265 10597
rect 2265 10571 2266 10597
rect 2238 10570 2266 10571
rect 2290 10597 2318 10598
rect 2290 10571 2291 10597
rect 2291 10571 2317 10597
rect 2317 10571 2318 10597
rect 2290 10570 2318 10571
rect 2342 10597 2370 10598
rect 2342 10571 2343 10597
rect 2343 10571 2369 10597
rect 2369 10571 2370 10597
rect 2342 10570 2370 10571
rect 6006 10374 6034 10402
rect 7350 10457 7378 10458
rect 7350 10431 7351 10457
rect 7351 10431 7377 10457
rect 7377 10431 7378 10457
rect 7350 10430 7378 10431
rect 7070 10374 7098 10402
rect 2086 9926 2114 9954
rect 2238 9813 2266 9814
rect 2238 9787 2239 9813
rect 2239 9787 2265 9813
rect 2265 9787 2266 9813
rect 2238 9786 2266 9787
rect 2290 9813 2318 9814
rect 2290 9787 2291 9813
rect 2291 9787 2317 9813
rect 2317 9787 2318 9813
rect 2290 9786 2318 9787
rect 2342 9813 2370 9814
rect 2342 9787 2343 9813
rect 2343 9787 2369 9813
rect 2369 9787 2370 9813
rect 2342 9786 2370 9787
rect 7070 9982 7098 10010
rect 5558 9225 5586 9226
rect 5558 9199 5559 9225
rect 5559 9199 5585 9225
rect 5585 9199 5586 9225
rect 5558 9198 5586 9199
rect 2238 9029 2266 9030
rect 2238 9003 2239 9029
rect 2239 9003 2265 9029
rect 2265 9003 2266 9029
rect 2238 9002 2266 9003
rect 2290 9029 2318 9030
rect 2290 9003 2291 9029
rect 2291 9003 2317 9029
rect 2317 9003 2318 9029
rect 2290 9002 2318 9003
rect 2342 9029 2370 9030
rect 2342 9003 2343 9029
rect 2343 9003 2369 9029
rect 2369 9003 2370 9029
rect 2342 9002 2370 9003
rect 2238 8245 2266 8246
rect 2238 8219 2239 8245
rect 2239 8219 2265 8245
rect 2265 8219 2266 8245
rect 2238 8218 2266 8219
rect 2290 8245 2318 8246
rect 2290 8219 2291 8245
rect 2291 8219 2317 8245
rect 2317 8219 2318 8245
rect 2290 8218 2318 8219
rect 2342 8245 2370 8246
rect 2342 8219 2343 8245
rect 2343 8219 2369 8245
rect 2369 8219 2370 8245
rect 2342 8218 2370 8219
rect 2142 8134 2170 8162
rect 966 8078 994 8106
rect 2142 8049 2170 8050
rect 2142 8023 2143 8049
rect 2143 8023 2169 8049
rect 2169 8023 2170 8049
rect 2142 8022 2170 8023
rect 5614 8022 5642 8050
rect 5614 7798 5642 7826
rect 5670 8134 5698 8162
rect 1022 7742 1050 7770
rect 7518 10430 7546 10458
rect 7406 10065 7434 10066
rect 7406 10039 7407 10065
rect 7407 10039 7433 10065
rect 7433 10039 7434 10065
rect 7406 10038 7434 10039
rect 7574 10009 7602 10010
rect 7574 9983 7575 10009
rect 7575 9983 7601 10009
rect 7601 9983 7602 10009
rect 7574 9982 7602 9983
rect 7182 9225 7210 9226
rect 7182 9199 7183 9225
rect 7183 9199 7209 9225
rect 7209 9199 7210 9225
rect 7182 9198 7210 9199
rect 7014 8526 7042 8554
rect 5894 8022 5922 8050
rect 6902 8049 6930 8050
rect 6902 8023 6903 8049
rect 6903 8023 6929 8049
rect 6929 8023 6930 8049
rect 6902 8022 6930 8023
rect 8582 11438 8610 11466
rect 8246 11073 8274 11074
rect 8246 11047 8247 11073
rect 8247 11047 8273 11073
rect 8273 11047 8274 11073
rect 8246 11046 8274 11047
rect 8358 10934 8386 10962
rect 7966 10878 7994 10906
rect 8414 10849 8442 10850
rect 8414 10823 8415 10849
rect 8415 10823 8441 10849
rect 8441 10823 8442 10849
rect 8414 10822 8442 10823
rect 7854 10457 7882 10458
rect 7854 10431 7855 10457
rect 7855 10431 7881 10457
rect 7881 10431 7882 10457
rect 7854 10430 7882 10431
rect 7742 9814 7770 9842
rect 7910 10038 7938 10066
rect 8190 10065 8218 10066
rect 8190 10039 8191 10065
rect 8191 10039 8217 10065
rect 8217 10039 8218 10065
rect 8190 10038 8218 10039
rect 8022 10009 8050 10010
rect 8022 9983 8023 10009
rect 8023 9983 8049 10009
rect 8049 9983 8050 10009
rect 8022 9982 8050 9983
rect 8414 9814 8442 9842
rect 7910 9534 7938 9562
rect 7966 9422 7994 9450
rect 8190 9142 8218 9170
rect 8302 8694 8330 8722
rect 7630 8526 7658 8554
rect 8190 8553 8218 8554
rect 8190 8527 8191 8553
rect 8191 8527 8217 8553
rect 8217 8527 8218 8553
rect 8190 8526 8218 8527
rect 7070 8078 7098 8106
rect 5670 7742 5698 7770
rect 6790 7686 6818 7714
rect 2238 7461 2266 7462
rect 2238 7435 2239 7461
rect 2239 7435 2265 7461
rect 2265 7435 2266 7461
rect 2238 7434 2266 7435
rect 2290 7461 2318 7462
rect 2290 7435 2291 7461
rect 2291 7435 2317 7461
rect 2317 7435 2318 7461
rect 2290 7434 2318 7435
rect 2342 7461 2370 7462
rect 2342 7435 2343 7461
rect 2343 7435 2369 7461
rect 2369 7435 2370 7461
rect 2342 7434 2370 7435
rect 6902 7798 6930 7826
rect 7406 8441 7434 8442
rect 7406 8415 7407 8441
rect 7407 8415 7433 8441
rect 7433 8415 7434 8441
rect 7406 8414 7434 8415
rect 7294 7769 7322 7770
rect 7294 7743 7295 7769
rect 7295 7743 7321 7769
rect 7321 7743 7322 7769
rect 7294 7742 7322 7743
rect 7518 8078 7546 8106
rect 8414 8078 8442 8106
rect 7462 7686 7490 7714
rect 7518 7742 7546 7770
rect 7014 7518 7042 7546
rect 7350 7630 7378 7658
rect 7182 7574 7210 7602
rect 7518 7574 7546 7602
rect 7742 7574 7770 7602
rect 7406 7518 7434 7546
rect 8638 11214 8666 11242
rect 8582 10878 8610 10906
rect 8526 9590 8554 9618
rect 8750 11185 8778 11186
rect 8750 11159 8751 11185
rect 8751 11159 8777 11185
rect 8777 11159 8778 11185
rect 8750 11158 8778 11159
rect 9142 12473 9170 12474
rect 9142 12447 9143 12473
rect 9143 12447 9169 12473
rect 9169 12447 9170 12473
rect 9142 12446 9170 12447
rect 9030 11718 9058 11746
rect 9422 12614 9450 12642
rect 9534 12838 9562 12866
rect 9310 11689 9338 11690
rect 9310 11663 9311 11689
rect 9311 11663 9337 11689
rect 9337 11663 9338 11689
rect 9310 11662 9338 11663
rect 9478 11577 9506 11578
rect 9478 11551 9479 11577
rect 9479 11551 9505 11577
rect 9505 11551 9506 11577
rect 9478 11550 9506 11551
rect 9198 11241 9226 11242
rect 9198 11215 9199 11241
rect 9199 11215 9225 11241
rect 9225 11215 9226 11241
rect 9198 11214 9226 11215
rect 9478 11185 9506 11186
rect 9478 11159 9479 11185
rect 9479 11159 9505 11185
rect 9505 11159 9506 11185
rect 9478 11158 9506 11159
rect 8750 10934 8778 10962
rect 9422 10934 9450 10962
rect 8750 9953 8778 9954
rect 8750 9927 8751 9953
rect 8751 9927 8777 9953
rect 8777 9927 8778 9953
rect 8750 9926 8778 9927
rect 8862 10822 8890 10850
rect 8750 9590 8778 9618
rect 8694 9505 8722 9506
rect 8694 9479 8695 9505
rect 8695 9479 8721 9505
rect 8721 9479 8722 9505
rect 8694 9478 8722 9479
rect 9366 10849 9394 10850
rect 9366 10823 9367 10849
rect 9367 10823 9393 10849
rect 9393 10823 9394 10849
rect 9366 10822 9394 10823
rect 8750 9198 8778 9226
rect 8862 9422 8890 9450
rect 9086 10793 9114 10794
rect 9086 10767 9087 10793
rect 9087 10767 9113 10793
rect 9113 10767 9114 10793
rect 9086 10766 9114 10767
rect 9366 10374 9394 10402
rect 9366 10094 9394 10122
rect 9086 9982 9114 10010
rect 9142 9814 9170 9842
rect 9254 9897 9282 9898
rect 9254 9871 9255 9897
rect 9255 9871 9281 9897
rect 9281 9871 9282 9897
rect 9254 9870 9282 9871
rect 8974 9617 9002 9618
rect 8974 9591 8975 9617
rect 8975 9591 9001 9617
rect 9001 9591 9002 9617
rect 8974 9590 9002 9591
rect 8918 9310 8946 9338
rect 8974 9478 9002 9506
rect 8918 8721 8946 8722
rect 8918 8695 8919 8721
rect 8919 8695 8945 8721
rect 8945 8695 8946 8721
rect 8918 8694 8946 8695
rect 9254 9534 9282 9562
rect 9310 9310 9338 9338
rect 9198 8777 9226 8778
rect 9198 8751 9199 8777
rect 9199 8751 9225 8777
rect 9225 8751 9226 8777
rect 9198 8750 9226 8751
rect 9310 8526 9338 8554
rect 10766 13566 10794 13594
rect 9918 13341 9946 13342
rect 9918 13315 9919 13341
rect 9919 13315 9945 13341
rect 9945 13315 9946 13341
rect 9918 13314 9946 13315
rect 9970 13341 9998 13342
rect 9970 13315 9971 13341
rect 9971 13315 9997 13341
rect 9997 13315 9998 13341
rect 9970 13314 9998 13315
rect 10022 13341 10050 13342
rect 10022 13315 10023 13341
rect 10023 13315 10049 13341
rect 10049 13315 10050 13341
rect 10022 13314 10050 13315
rect 10934 13398 10962 13426
rect 10654 12865 10682 12866
rect 10654 12839 10655 12865
rect 10655 12839 10681 12865
rect 10681 12839 10682 12865
rect 10654 12838 10682 12839
rect 10822 12809 10850 12810
rect 10822 12783 10823 12809
rect 10823 12783 10849 12809
rect 10849 12783 10850 12809
rect 10822 12782 10850 12783
rect 10598 12726 10626 12754
rect 9926 12641 9954 12642
rect 9926 12615 9927 12641
rect 9927 12615 9953 12641
rect 9953 12615 9954 12641
rect 9926 12614 9954 12615
rect 9918 12557 9946 12558
rect 9918 12531 9919 12557
rect 9919 12531 9945 12557
rect 9945 12531 9946 12557
rect 9918 12530 9946 12531
rect 9970 12557 9998 12558
rect 9970 12531 9971 12557
rect 9971 12531 9997 12557
rect 9997 12531 9998 12557
rect 9970 12530 9998 12531
rect 10022 12557 10050 12558
rect 10022 12531 10023 12557
rect 10023 12531 10049 12557
rect 10049 12531 10050 12557
rect 10022 12530 10050 12531
rect 10262 12446 10290 12474
rect 9918 11773 9946 11774
rect 9758 11718 9786 11746
rect 9918 11747 9919 11773
rect 9919 11747 9945 11773
rect 9945 11747 9946 11773
rect 9918 11746 9946 11747
rect 9970 11773 9998 11774
rect 9970 11747 9971 11773
rect 9971 11747 9997 11773
rect 9997 11747 9998 11773
rect 9970 11746 9998 11747
rect 10022 11773 10050 11774
rect 10022 11747 10023 11773
rect 10023 11747 10049 11773
rect 10049 11747 10050 11773
rect 10022 11746 10050 11747
rect 9590 11326 9618 11354
rect 9646 11270 9674 11298
rect 9758 10934 9786 10962
rect 9534 9870 9562 9898
rect 9478 9505 9506 9506
rect 9478 9479 9479 9505
rect 9479 9479 9505 9505
rect 9505 9479 9506 9505
rect 9478 9478 9506 9479
rect 10150 11550 10178 11578
rect 9918 10989 9946 10990
rect 9918 10963 9919 10989
rect 9919 10963 9945 10989
rect 9945 10963 9946 10989
rect 9918 10962 9946 10963
rect 9970 10989 9998 10990
rect 9970 10963 9971 10989
rect 9971 10963 9997 10989
rect 9997 10963 9998 10989
rect 9970 10962 9998 10963
rect 10022 10989 10050 10990
rect 10022 10963 10023 10989
rect 10023 10963 10049 10989
rect 10049 10963 10050 10989
rect 10022 10962 10050 10963
rect 9758 10793 9786 10794
rect 9758 10767 9759 10793
rect 9759 10767 9785 10793
rect 9785 10767 9786 10793
rect 9758 10766 9786 10767
rect 9870 10654 9898 10682
rect 10038 10318 10066 10346
rect 9918 10205 9946 10206
rect 9918 10179 9919 10205
rect 9919 10179 9945 10205
rect 9945 10179 9946 10205
rect 9918 10178 9946 10179
rect 9970 10205 9998 10206
rect 9970 10179 9971 10205
rect 9971 10179 9997 10205
rect 9997 10179 9998 10205
rect 9970 10178 9998 10179
rect 10022 10205 10050 10206
rect 10022 10179 10023 10205
rect 10023 10179 10049 10205
rect 10049 10179 10050 10205
rect 10022 10178 10050 10179
rect 10094 10038 10122 10066
rect 9702 9926 9730 9954
rect 9870 9758 9898 9786
rect 10038 9702 10066 9730
rect 9918 9421 9946 9422
rect 9918 9395 9919 9421
rect 9919 9395 9945 9421
rect 9945 9395 9946 9421
rect 9918 9394 9946 9395
rect 9970 9421 9998 9422
rect 9970 9395 9971 9421
rect 9971 9395 9997 9421
rect 9997 9395 9998 9421
rect 9970 9394 9998 9395
rect 10022 9421 10050 9422
rect 10022 9395 10023 9421
rect 10023 9395 10049 9421
rect 10049 9395 10050 9421
rect 10022 9394 10050 9395
rect 9758 9225 9786 9226
rect 9758 9199 9759 9225
rect 9759 9199 9785 9225
rect 9785 9199 9786 9225
rect 9758 9198 9786 9199
rect 9646 9169 9674 9170
rect 9646 9143 9647 9169
rect 9647 9143 9673 9169
rect 9673 9143 9674 9169
rect 9646 9142 9674 9143
rect 9590 9086 9618 9114
rect 9142 8470 9170 8498
rect 8974 8441 9002 8442
rect 8974 8415 8975 8441
rect 8975 8415 9001 8441
rect 9001 8415 9002 8441
rect 8974 8414 9002 8415
rect 9254 8329 9282 8330
rect 9254 8303 9255 8329
rect 9255 8303 9281 8329
rect 9281 8303 9282 8329
rect 9254 8302 9282 8303
rect 8862 7798 8890 7826
rect 8470 7518 8498 7546
rect 8694 7518 8722 7546
rect 8918 7657 8946 7658
rect 8918 7631 8919 7657
rect 8919 7631 8945 7657
rect 8945 7631 8946 7657
rect 8918 7630 8946 7631
rect 9366 8246 9394 8274
rect 9422 8105 9450 8106
rect 9422 8079 9423 8105
rect 9423 8079 9449 8105
rect 9449 8079 9450 8105
rect 9422 8078 9450 8079
rect 9534 8497 9562 8498
rect 9534 8471 9535 8497
rect 9535 8471 9561 8497
rect 9561 8471 9562 8497
rect 9534 8470 9562 8471
rect 9870 9225 9898 9226
rect 9870 9199 9871 9225
rect 9871 9199 9897 9225
rect 9897 9199 9898 9225
rect 9870 9198 9898 9199
rect 10206 9310 10234 9338
rect 9982 9142 10010 9170
rect 9702 8750 9730 8778
rect 10094 9113 10122 9114
rect 10094 9087 10095 9113
rect 10095 9087 10121 9113
rect 10121 9087 10122 9113
rect 10094 9086 10122 9087
rect 9918 8637 9946 8638
rect 9918 8611 9919 8637
rect 9919 8611 9945 8637
rect 9945 8611 9946 8637
rect 9918 8610 9946 8611
rect 9970 8637 9998 8638
rect 9970 8611 9971 8637
rect 9971 8611 9997 8637
rect 9997 8611 9998 8637
rect 9970 8610 9998 8611
rect 10022 8637 10050 8638
rect 10022 8611 10023 8637
rect 10023 8611 10049 8637
rect 10049 8611 10050 8637
rect 10022 8610 10050 8611
rect 9702 8414 9730 8442
rect 9030 7910 9058 7938
rect 9478 7910 9506 7938
rect 9590 8302 9618 8330
rect 9478 7798 9506 7826
rect 9142 7713 9170 7714
rect 9142 7687 9143 7713
rect 9143 7687 9169 7713
rect 9169 7687 9170 7713
rect 9142 7686 9170 7687
rect 10542 11942 10570 11970
rect 10374 11326 10402 11354
rect 10318 10878 10346 10906
rect 10374 11046 10402 11074
rect 10318 10430 10346 10458
rect 10374 9982 10402 10010
rect 10486 10878 10514 10906
rect 10430 9337 10458 9338
rect 10430 9311 10431 9337
rect 10431 9311 10457 9337
rect 10457 9311 10458 9337
rect 10430 9310 10458 9311
rect 10878 12726 10906 12754
rect 10990 13454 11018 13482
rect 11774 13902 11802 13930
rect 11662 13873 11690 13874
rect 11662 13847 11663 13873
rect 11663 13847 11689 13873
rect 11689 13847 11690 13873
rect 11662 13846 11690 13847
rect 11550 13790 11578 13818
rect 11382 13566 11410 13594
rect 11774 13537 11802 13538
rect 11774 13511 11775 13537
rect 11775 13511 11801 13537
rect 11801 13511 11802 13537
rect 11774 13510 11802 13511
rect 11326 13398 11354 13426
rect 11606 13454 11634 13482
rect 11774 13398 11802 13426
rect 11102 13118 11130 13146
rect 11158 13174 11186 13202
rect 11158 12782 11186 12810
rect 10710 12473 10738 12474
rect 10710 12447 10711 12473
rect 10711 12447 10737 12473
rect 10737 12447 10738 12473
rect 10710 12446 10738 12447
rect 10766 11886 10794 11914
rect 10710 11577 10738 11578
rect 10710 11551 10711 11577
rect 10711 11551 10737 11577
rect 10737 11551 10738 11577
rect 10710 11550 10738 11551
rect 11046 11886 11074 11914
rect 10934 11606 10962 11634
rect 10878 11550 10906 11578
rect 10990 11326 11018 11354
rect 11270 13145 11298 13146
rect 11270 13119 11271 13145
rect 11271 13119 11297 13145
rect 11297 13119 11298 13145
rect 11270 13118 11298 13119
rect 11158 11494 11186 11522
rect 11942 13929 11970 13930
rect 11942 13903 11943 13929
rect 11943 13903 11969 13929
rect 11969 13903 11970 13929
rect 11942 13902 11970 13903
rect 17598 19221 17626 19222
rect 17598 19195 17599 19221
rect 17599 19195 17625 19221
rect 17625 19195 17626 19221
rect 17598 19194 17626 19195
rect 17650 19221 17678 19222
rect 17650 19195 17651 19221
rect 17651 19195 17677 19221
rect 17677 19195 17678 19221
rect 17650 19194 17678 19195
rect 17702 19221 17730 19222
rect 17702 19195 17703 19221
rect 17703 19195 17729 19221
rect 17729 19195 17730 19221
rect 17702 19194 17730 19195
rect 14686 19137 14714 19138
rect 14686 19111 14687 19137
rect 14687 19111 14713 19137
rect 14713 19111 14714 19137
rect 14686 19110 14714 19111
rect 13118 14041 13146 14042
rect 13118 14015 13119 14041
rect 13119 14015 13145 14041
rect 13145 14015 13146 14041
rect 13118 14014 13146 14015
rect 17598 18437 17626 18438
rect 17598 18411 17599 18437
rect 17599 18411 17625 18437
rect 17625 18411 17626 18437
rect 17598 18410 17626 18411
rect 17650 18437 17678 18438
rect 17650 18411 17651 18437
rect 17651 18411 17677 18437
rect 17677 18411 17678 18437
rect 17650 18410 17678 18411
rect 17702 18437 17730 18438
rect 17702 18411 17703 18437
rect 17703 18411 17729 18437
rect 17729 18411 17730 18437
rect 17702 18410 17730 18411
rect 17598 17653 17626 17654
rect 17598 17627 17599 17653
rect 17599 17627 17625 17653
rect 17625 17627 17626 17653
rect 17598 17626 17626 17627
rect 17650 17653 17678 17654
rect 17650 17627 17651 17653
rect 17651 17627 17677 17653
rect 17677 17627 17678 17653
rect 17650 17626 17678 17627
rect 17702 17653 17730 17654
rect 17702 17627 17703 17653
rect 17703 17627 17729 17653
rect 17729 17627 17730 17653
rect 17702 17626 17730 17627
rect 17598 16869 17626 16870
rect 17598 16843 17599 16869
rect 17599 16843 17625 16869
rect 17625 16843 17626 16869
rect 17598 16842 17626 16843
rect 17650 16869 17678 16870
rect 17650 16843 17651 16869
rect 17651 16843 17677 16869
rect 17677 16843 17678 16869
rect 17650 16842 17678 16843
rect 17702 16869 17730 16870
rect 17702 16843 17703 16869
rect 17703 16843 17729 16869
rect 17729 16843 17730 16869
rect 17702 16842 17730 16843
rect 17598 16085 17626 16086
rect 17598 16059 17599 16085
rect 17599 16059 17625 16085
rect 17625 16059 17626 16085
rect 17598 16058 17626 16059
rect 17650 16085 17678 16086
rect 17650 16059 17651 16085
rect 17651 16059 17677 16085
rect 17677 16059 17678 16085
rect 17650 16058 17678 16059
rect 17702 16085 17730 16086
rect 17702 16059 17703 16085
rect 17703 16059 17729 16085
rect 17729 16059 17730 16085
rect 17702 16058 17730 16059
rect 17598 15301 17626 15302
rect 17598 15275 17599 15301
rect 17599 15275 17625 15301
rect 17625 15275 17626 15301
rect 17598 15274 17626 15275
rect 17650 15301 17678 15302
rect 17650 15275 17651 15301
rect 17651 15275 17677 15301
rect 17677 15275 17678 15301
rect 17650 15274 17678 15275
rect 17702 15301 17730 15302
rect 17702 15275 17703 15301
rect 17703 15275 17729 15301
rect 17729 15275 17730 15301
rect 17702 15274 17730 15275
rect 17598 14517 17626 14518
rect 17598 14491 17599 14517
rect 17599 14491 17625 14517
rect 17625 14491 17626 14517
rect 17598 14490 17626 14491
rect 17650 14517 17678 14518
rect 17650 14491 17651 14517
rect 17651 14491 17677 14517
rect 17677 14491 17678 14517
rect 17650 14490 17678 14491
rect 17702 14517 17730 14518
rect 17702 14491 17703 14517
rect 17703 14491 17729 14517
rect 17729 14491 17730 14517
rect 17702 14490 17730 14491
rect 14294 14014 14322 14042
rect 12278 13846 12306 13874
rect 12110 13481 12138 13482
rect 12110 13455 12111 13481
rect 12111 13455 12137 13481
rect 12137 13455 12138 13481
rect 12110 13454 12138 13455
rect 12110 13201 12138 13202
rect 12110 13175 12111 13201
rect 12111 13175 12137 13201
rect 12137 13175 12138 13201
rect 12110 13174 12138 13175
rect 12614 13817 12642 13818
rect 12614 13791 12615 13817
rect 12615 13791 12641 13817
rect 12641 13791 12642 13817
rect 12614 13790 12642 13791
rect 17598 13733 17626 13734
rect 17598 13707 17599 13733
rect 17599 13707 17625 13733
rect 17625 13707 17626 13733
rect 17598 13706 17626 13707
rect 17650 13733 17678 13734
rect 17650 13707 17651 13733
rect 17651 13707 17677 13733
rect 17677 13707 17678 13733
rect 17650 13706 17678 13707
rect 17702 13733 17730 13734
rect 17702 13707 17703 13733
rect 17703 13707 17729 13733
rect 17729 13707 17730 13733
rect 17702 13706 17730 13707
rect 12614 13510 12642 13538
rect 13398 13537 13426 13538
rect 13398 13511 13399 13537
rect 13399 13511 13425 13537
rect 13425 13511 13426 13537
rect 13398 13510 13426 13511
rect 13398 13230 13426 13258
rect 13678 13230 13706 13258
rect 13286 13118 13314 13146
rect 12278 13062 12306 13090
rect 13006 13089 13034 13090
rect 13006 13063 13007 13089
rect 13007 13063 13033 13089
rect 13033 13063 13034 13089
rect 13006 13062 13034 13063
rect 12334 12753 12362 12754
rect 12334 12727 12335 12753
rect 12335 12727 12361 12753
rect 12361 12727 12362 12753
rect 12334 12726 12362 12727
rect 13174 12753 13202 12754
rect 13174 12727 13175 12753
rect 13175 12727 13201 12753
rect 13201 12727 13202 12753
rect 13174 12726 13202 12727
rect 13286 12278 13314 12306
rect 11942 11969 11970 11970
rect 11942 11943 11943 11969
rect 11943 11943 11969 11969
rect 11969 11943 11970 11969
rect 11942 11942 11970 11943
rect 11382 11550 11410 11578
rect 11046 11214 11074 11242
rect 10878 11102 10906 11130
rect 10654 11073 10682 11074
rect 10654 11047 10655 11073
rect 10655 11047 10681 11073
rect 10681 11047 10682 11073
rect 10654 11046 10682 11047
rect 10878 10878 10906 10906
rect 10598 10793 10626 10794
rect 10598 10767 10599 10793
rect 10599 10767 10625 10793
rect 10625 10767 10626 10793
rect 10598 10766 10626 10767
rect 11102 10766 11130 10794
rect 10710 9729 10738 9730
rect 10710 9703 10711 9729
rect 10711 9703 10737 9729
rect 10737 9703 10738 9729
rect 10710 9702 10738 9703
rect 11046 10318 11074 10346
rect 11158 10430 11186 10458
rect 10654 9561 10682 9562
rect 10654 9535 10655 9561
rect 10655 9535 10681 9561
rect 10681 9535 10682 9561
rect 10654 9534 10682 9535
rect 10654 9169 10682 9170
rect 10654 9143 10655 9169
rect 10655 9143 10681 9169
rect 10681 9143 10682 9169
rect 10654 9142 10682 9143
rect 10654 8526 10682 8554
rect 11046 10065 11074 10066
rect 11046 10039 11047 10065
rect 11047 10039 11073 10065
rect 11073 10039 11074 10065
rect 11046 10038 11074 10039
rect 10990 9310 11018 9338
rect 11606 11494 11634 11522
rect 11270 10654 11298 10682
rect 11774 11326 11802 11354
rect 11718 11158 11746 11186
rect 11494 10457 11522 10458
rect 11494 10431 11495 10457
rect 11495 10431 11521 10457
rect 11521 10431 11522 10457
rect 11494 10430 11522 10431
rect 11270 10401 11298 10402
rect 11270 10375 11271 10401
rect 11271 10375 11297 10401
rect 11297 10375 11298 10401
rect 11270 10374 11298 10375
rect 11214 10094 11242 10122
rect 10934 9142 10962 9170
rect 11382 9617 11410 9618
rect 11382 9591 11383 9617
rect 11383 9591 11409 9617
rect 11409 9591 11410 9617
rect 11382 9590 11410 9591
rect 11438 9254 11466 9282
rect 11158 9030 11186 9058
rect 11438 8889 11466 8890
rect 11438 8863 11439 8889
rect 11439 8863 11465 8889
rect 11465 8863 11466 8889
rect 11438 8862 11466 8863
rect 10878 8526 10906 8554
rect 10262 8246 10290 8274
rect 10094 8022 10122 8050
rect 9086 7574 9114 7602
rect 8918 6958 8946 6986
rect 2238 6677 2266 6678
rect 2238 6651 2239 6677
rect 2239 6651 2265 6677
rect 2265 6651 2266 6677
rect 2238 6650 2266 6651
rect 2290 6677 2318 6678
rect 2290 6651 2291 6677
rect 2291 6651 2317 6677
rect 2317 6651 2318 6677
rect 2290 6650 2318 6651
rect 2342 6677 2370 6678
rect 2342 6651 2343 6677
rect 2343 6651 2369 6677
rect 2369 6651 2370 6677
rect 2342 6650 2370 6651
rect 2238 5893 2266 5894
rect 2238 5867 2239 5893
rect 2239 5867 2265 5893
rect 2265 5867 2266 5893
rect 2238 5866 2266 5867
rect 2290 5893 2318 5894
rect 2290 5867 2291 5893
rect 2291 5867 2317 5893
rect 2317 5867 2318 5893
rect 2290 5866 2318 5867
rect 2342 5893 2370 5894
rect 2342 5867 2343 5893
rect 2343 5867 2369 5893
rect 2369 5867 2370 5893
rect 2342 5866 2370 5867
rect 8974 7126 9002 7154
rect 9702 7657 9730 7658
rect 9702 7631 9703 7657
rect 9703 7631 9729 7657
rect 9729 7631 9730 7657
rect 9702 7630 9730 7631
rect 9646 7601 9674 7602
rect 9646 7575 9647 7601
rect 9647 7575 9673 7601
rect 9673 7575 9674 7601
rect 9646 7574 9674 7575
rect 9758 7518 9786 7546
rect 9590 7153 9618 7154
rect 9590 7127 9591 7153
rect 9591 7127 9617 7153
rect 9617 7127 9618 7153
rect 9590 7126 9618 7127
rect 9254 6958 9282 6986
rect 8470 5838 8498 5866
rect 2238 5109 2266 5110
rect 2238 5083 2239 5109
rect 2239 5083 2265 5109
rect 2265 5083 2266 5109
rect 2238 5082 2266 5083
rect 2290 5109 2318 5110
rect 2290 5083 2291 5109
rect 2291 5083 2317 5109
rect 2317 5083 2318 5109
rect 2290 5082 2318 5083
rect 2342 5109 2370 5110
rect 2342 5083 2343 5109
rect 2343 5083 2369 5109
rect 2369 5083 2370 5109
rect 2342 5082 2370 5083
rect 2238 4325 2266 4326
rect 2238 4299 2239 4325
rect 2239 4299 2265 4325
rect 2265 4299 2266 4325
rect 2238 4298 2266 4299
rect 2290 4325 2318 4326
rect 2290 4299 2291 4325
rect 2291 4299 2317 4325
rect 2317 4299 2318 4325
rect 2290 4298 2318 4299
rect 2342 4325 2370 4326
rect 2342 4299 2343 4325
rect 2343 4299 2369 4325
rect 2369 4299 2370 4325
rect 2342 4298 2370 4299
rect 9918 7853 9946 7854
rect 9918 7827 9919 7853
rect 9919 7827 9945 7853
rect 9945 7827 9946 7853
rect 9918 7826 9946 7827
rect 9970 7853 9998 7854
rect 9970 7827 9971 7853
rect 9971 7827 9997 7853
rect 9997 7827 9998 7853
rect 9970 7826 9998 7827
rect 10022 7853 10050 7854
rect 10022 7827 10023 7853
rect 10023 7827 10049 7853
rect 10049 7827 10050 7853
rect 10022 7826 10050 7827
rect 10318 7742 10346 7770
rect 10710 8022 10738 8050
rect 10486 7574 10514 7602
rect 10822 7657 10850 7658
rect 10822 7631 10823 7657
rect 10823 7631 10849 7657
rect 10849 7631 10850 7657
rect 10822 7630 10850 7631
rect 11662 10710 11690 10738
rect 11998 11633 12026 11634
rect 11998 11607 11999 11633
rect 11999 11607 12025 11633
rect 12025 11607 12026 11633
rect 11998 11606 12026 11607
rect 14294 13257 14322 13258
rect 14294 13231 14295 13257
rect 14295 13231 14321 13257
rect 14321 13231 14322 13257
rect 14294 13230 14322 13231
rect 14070 13118 14098 13146
rect 18830 13118 18858 13146
rect 20006 13118 20034 13146
rect 17598 12949 17626 12950
rect 17598 12923 17599 12949
rect 17599 12923 17625 12949
rect 17625 12923 17626 12949
rect 17598 12922 17626 12923
rect 17650 12949 17678 12950
rect 17650 12923 17651 12949
rect 17651 12923 17677 12949
rect 17677 12923 17678 12949
rect 17650 12922 17678 12923
rect 17702 12949 17730 12950
rect 17702 12923 17703 12949
rect 17703 12923 17729 12949
rect 17729 12923 17730 12949
rect 17702 12922 17730 12923
rect 13342 11662 13370 11690
rect 13566 11830 13594 11858
rect 12894 11606 12922 11634
rect 11998 10878 12026 10906
rect 11662 10094 11690 10122
rect 12110 10878 12138 10906
rect 13062 10822 13090 10850
rect 12334 10793 12362 10794
rect 12334 10767 12335 10793
rect 12335 10767 12361 10793
rect 12361 10767 12362 10793
rect 12334 10766 12362 10767
rect 12726 10766 12754 10794
rect 11662 9254 11690 9282
rect 11606 9169 11634 9170
rect 11606 9143 11607 9169
rect 11607 9143 11633 9169
rect 11633 9143 11634 9169
rect 11606 9142 11634 9143
rect 11830 9366 11858 9394
rect 11998 9478 12026 9506
rect 11886 9086 11914 9114
rect 11102 8526 11130 8554
rect 11326 8582 11354 8610
rect 11438 8385 11466 8386
rect 11438 8359 11439 8385
rect 11439 8359 11465 8385
rect 11465 8359 11466 8385
rect 11438 8358 11466 8359
rect 11046 7966 11074 7994
rect 11438 8246 11466 8274
rect 11046 7630 11074 7658
rect 11214 7769 11242 7770
rect 11214 7743 11215 7769
rect 11215 7743 11241 7769
rect 11241 7743 11242 7769
rect 11214 7742 11242 7743
rect 10934 7518 10962 7546
rect 11326 7574 11354 7602
rect 11718 8526 11746 8554
rect 11830 8302 11858 8330
rect 11942 9030 11970 9058
rect 12782 10737 12810 10738
rect 12782 10711 12783 10737
rect 12783 10711 12809 10737
rect 12809 10711 12810 10737
rect 12782 10710 12810 10711
rect 13118 10710 13146 10738
rect 13286 10766 13314 10794
rect 18830 12361 18858 12362
rect 18830 12335 18831 12361
rect 18831 12335 18857 12361
rect 18857 12335 18858 12361
rect 18830 12334 18858 12335
rect 14238 12305 14266 12306
rect 14238 12279 14239 12305
rect 14239 12279 14265 12305
rect 14265 12279 14266 12305
rect 14238 12278 14266 12279
rect 15302 12305 15330 12306
rect 15302 12279 15303 12305
rect 15303 12279 15329 12305
rect 15329 12279 15330 12305
rect 15302 12278 15330 12279
rect 13958 11969 13986 11970
rect 13958 11943 13959 11969
rect 13959 11943 13985 11969
rect 13985 11943 13986 11969
rect 13958 11942 13986 11943
rect 17598 12165 17626 12166
rect 17598 12139 17599 12165
rect 17599 12139 17625 12165
rect 17625 12139 17626 12165
rect 17598 12138 17626 12139
rect 17650 12165 17678 12166
rect 17650 12139 17651 12165
rect 17651 12139 17677 12165
rect 17677 12139 17678 12165
rect 17650 12138 17678 12139
rect 17702 12165 17730 12166
rect 17702 12139 17703 12165
rect 17703 12139 17729 12165
rect 17729 12139 17730 12165
rect 17702 12138 17730 12139
rect 20006 12110 20034 12138
rect 15302 11942 15330 11970
rect 13902 11857 13930 11858
rect 13902 11831 13903 11857
rect 13903 11831 13929 11857
rect 13929 11831 13930 11857
rect 13902 11830 13930 11831
rect 13846 11606 13874 11634
rect 20006 11774 20034 11802
rect 18830 11718 18858 11746
rect 14070 11662 14098 11690
rect 13566 11046 13594 11074
rect 13510 10849 13538 10850
rect 13510 10823 13511 10849
rect 13511 10823 13537 10849
rect 13537 10823 13538 10849
rect 13510 10822 13538 10823
rect 13062 9758 13090 9786
rect 13286 9729 13314 9730
rect 13286 9703 13287 9729
rect 13287 9703 13313 9729
rect 13313 9703 13314 9729
rect 13286 9702 13314 9703
rect 13342 10374 13370 10402
rect 12950 9617 12978 9618
rect 12950 9591 12951 9617
rect 12951 9591 12977 9617
rect 12977 9591 12978 9617
rect 12950 9590 12978 9591
rect 13174 9617 13202 9618
rect 13174 9591 13175 9617
rect 13175 9591 13201 9617
rect 13201 9591 13202 9617
rect 13174 9590 13202 9591
rect 13510 10430 13538 10458
rect 13398 10065 13426 10066
rect 13398 10039 13399 10065
rect 13399 10039 13425 10065
rect 13425 10039 13426 10065
rect 13398 10038 13426 10039
rect 13454 9617 13482 9618
rect 13454 9591 13455 9617
rect 13455 9591 13481 9617
rect 13481 9591 13482 9617
rect 13454 9590 13482 9591
rect 13342 9534 13370 9562
rect 12838 9505 12866 9506
rect 12838 9479 12839 9505
rect 12839 9479 12865 9505
rect 12865 9479 12866 9505
rect 12838 9478 12866 9479
rect 13454 9478 13482 9506
rect 12222 9366 12250 9394
rect 13454 9254 13482 9282
rect 12502 9142 12530 9170
rect 15414 11633 15442 11634
rect 15414 11607 15415 11633
rect 15415 11607 15441 11633
rect 15441 11607 15442 11633
rect 15414 11606 15442 11607
rect 15246 11577 15274 11578
rect 15246 11551 15247 11577
rect 15247 11551 15273 11577
rect 15273 11551 15274 11577
rect 15246 11550 15274 11551
rect 18830 11577 18858 11578
rect 18830 11551 18831 11577
rect 18831 11551 18857 11577
rect 18857 11551 18858 11577
rect 18830 11550 18858 11551
rect 13790 11185 13818 11186
rect 13790 11159 13791 11185
rect 13791 11159 13817 11185
rect 13817 11159 13818 11185
rect 13790 11158 13818 11159
rect 14014 11185 14042 11186
rect 14014 11159 14015 11185
rect 14015 11159 14041 11185
rect 14041 11159 14042 11185
rect 14014 11158 14042 11159
rect 14238 11158 14266 11186
rect 14182 11129 14210 11130
rect 14182 11103 14183 11129
rect 14183 11103 14209 11129
rect 14209 11103 14210 11129
rect 14182 11102 14210 11103
rect 20006 11465 20034 11466
rect 20006 11439 20007 11465
rect 20007 11439 20033 11465
rect 20033 11439 20034 11465
rect 20006 11438 20034 11439
rect 17598 11381 17626 11382
rect 17598 11355 17599 11381
rect 17599 11355 17625 11381
rect 17625 11355 17626 11381
rect 17598 11354 17626 11355
rect 17650 11381 17678 11382
rect 17650 11355 17651 11381
rect 17651 11355 17677 11381
rect 17677 11355 17678 11381
rect 17650 11354 17678 11355
rect 17702 11381 17730 11382
rect 17702 11355 17703 11381
rect 17703 11355 17729 11381
rect 17729 11355 17730 11381
rect 17702 11354 17730 11355
rect 15078 11102 15106 11130
rect 13734 10878 13762 10906
rect 13734 10457 13762 10458
rect 13734 10431 13735 10457
rect 13735 10431 13761 10457
rect 13761 10431 13762 10457
rect 13734 10430 13762 10431
rect 13622 9702 13650 9730
rect 13678 9422 13706 9450
rect 17598 10597 17626 10598
rect 17598 10571 17599 10597
rect 17599 10571 17625 10597
rect 17625 10571 17626 10597
rect 17598 10570 17626 10571
rect 17650 10597 17678 10598
rect 17650 10571 17651 10597
rect 17651 10571 17677 10597
rect 17677 10571 17678 10597
rect 17650 10570 17678 10571
rect 17702 10597 17730 10598
rect 17702 10571 17703 10597
rect 17703 10571 17729 10597
rect 17729 10571 17730 10597
rect 17702 10570 17730 10571
rect 14294 10038 14322 10066
rect 14070 9561 14098 9562
rect 14070 9535 14071 9561
rect 14071 9535 14097 9561
rect 14097 9535 14098 9561
rect 14070 9534 14098 9535
rect 14182 9561 14210 9562
rect 14182 9535 14183 9561
rect 14183 9535 14209 9561
rect 14209 9535 14210 9561
rect 14182 9534 14210 9535
rect 13958 9478 13986 9506
rect 15302 9982 15330 10010
rect 14350 9422 14378 9450
rect 14182 9254 14210 9282
rect 12894 8694 12922 8722
rect 13118 8721 13146 8722
rect 13118 8695 13119 8721
rect 13119 8695 13145 8721
rect 13145 8695 13146 8721
rect 13118 8694 13146 8695
rect 13454 8694 13482 8722
rect 12110 8302 12138 8330
rect 11830 7657 11858 7658
rect 11830 7631 11831 7657
rect 11831 7631 11857 7657
rect 11857 7631 11858 7657
rect 11830 7630 11858 7631
rect 11998 7686 12026 7714
rect 13678 8694 13706 8722
rect 13846 8358 13874 8386
rect 13454 7742 13482 7770
rect 12054 7657 12082 7658
rect 12054 7631 12055 7657
rect 12055 7631 12081 7657
rect 12081 7631 12082 7657
rect 12054 7630 12082 7631
rect 13118 7630 13146 7658
rect 12334 7574 12362 7602
rect 9918 7069 9946 7070
rect 9918 7043 9919 7069
rect 9919 7043 9945 7069
rect 9945 7043 9946 7069
rect 9918 7042 9946 7043
rect 9970 7069 9998 7070
rect 9970 7043 9971 7069
rect 9971 7043 9997 7069
rect 9997 7043 9998 7069
rect 9970 7042 9998 7043
rect 10022 7069 10050 7070
rect 10022 7043 10023 7069
rect 10023 7043 10049 7069
rect 10049 7043 10050 7069
rect 10022 7042 10050 7043
rect 9758 6958 9786 6986
rect 10206 6790 10234 6818
rect 10934 6873 10962 6874
rect 10934 6847 10935 6873
rect 10935 6847 10961 6873
rect 10961 6847 10962 6873
rect 10934 6846 10962 6847
rect 11662 6846 11690 6874
rect 12670 6873 12698 6874
rect 12670 6847 12671 6873
rect 12671 6847 12697 6873
rect 12697 6847 12698 6873
rect 12670 6846 12698 6847
rect 8862 5838 8890 5866
rect 2238 3541 2266 3542
rect 2238 3515 2239 3541
rect 2239 3515 2265 3541
rect 2265 3515 2266 3541
rect 2238 3514 2266 3515
rect 2290 3541 2318 3542
rect 2290 3515 2291 3541
rect 2291 3515 2317 3541
rect 2317 3515 2318 3541
rect 2290 3514 2318 3515
rect 2342 3541 2370 3542
rect 2342 3515 2343 3541
rect 2343 3515 2369 3541
rect 2369 3515 2370 3541
rect 2342 3514 2370 3515
rect 2238 2757 2266 2758
rect 2238 2731 2239 2757
rect 2239 2731 2265 2757
rect 2265 2731 2266 2757
rect 2238 2730 2266 2731
rect 2290 2757 2318 2758
rect 2290 2731 2291 2757
rect 2291 2731 2317 2757
rect 2317 2731 2318 2757
rect 2290 2730 2318 2731
rect 2342 2757 2370 2758
rect 2342 2731 2343 2757
rect 2343 2731 2369 2757
rect 2369 2731 2370 2757
rect 2342 2730 2370 2731
rect 8750 2590 8778 2618
rect 2238 1973 2266 1974
rect 2238 1947 2239 1973
rect 2239 1947 2265 1973
rect 2265 1947 2266 1973
rect 2238 1946 2266 1947
rect 2290 1973 2318 1974
rect 2290 1947 2291 1973
rect 2291 1947 2317 1973
rect 2317 1947 2318 1973
rect 2290 1946 2318 1947
rect 2342 1973 2370 1974
rect 2342 1947 2343 1973
rect 2343 1947 2369 1973
rect 2369 1947 2370 1973
rect 2342 1946 2370 1947
rect 9366 2617 9394 2618
rect 9366 2591 9367 2617
rect 9367 2591 9393 2617
rect 9393 2591 9394 2617
rect 9366 2590 9394 2591
rect 9918 6285 9946 6286
rect 9918 6259 9919 6285
rect 9919 6259 9945 6285
rect 9945 6259 9946 6285
rect 9918 6258 9946 6259
rect 9970 6285 9998 6286
rect 9970 6259 9971 6285
rect 9971 6259 9997 6285
rect 9997 6259 9998 6285
rect 9970 6258 9998 6259
rect 10022 6285 10050 6286
rect 10022 6259 10023 6285
rect 10023 6259 10049 6285
rect 10049 6259 10050 6285
rect 10022 6258 10050 6259
rect 9918 5501 9946 5502
rect 9918 5475 9919 5501
rect 9919 5475 9945 5501
rect 9945 5475 9946 5501
rect 9918 5474 9946 5475
rect 9970 5501 9998 5502
rect 9970 5475 9971 5501
rect 9971 5475 9997 5501
rect 9997 5475 9998 5501
rect 9970 5474 9998 5475
rect 10022 5501 10050 5502
rect 10022 5475 10023 5501
rect 10023 5475 10049 5501
rect 10049 5475 10050 5501
rect 10022 5474 10050 5475
rect 9918 4717 9946 4718
rect 9918 4691 9919 4717
rect 9919 4691 9945 4717
rect 9945 4691 9946 4717
rect 9918 4690 9946 4691
rect 9970 4717 9998 4718
rect 9970 4691 9971 4717
rect 9971 4691 9997 4717
rect 9997 4691 9998 4717
rect 9970 4690 9998 4691
rect 10022 4717 10050 4718
rect 10022 4691 10023 4717
rect 10023 4691 10049 4717
rect 10049 4691 10050 4717
rect 10022 4690 10050 4691
rect 9918 3933 9946 3934
rect 9918 3907 9919 3933
rect 9919 3907 9945 3933
rect 9945 3907 9946 3933
rect 9918 3906 9946 3907
rect 9970 3933 9998 3934
rect 9970 3907 9971 3933
rect 9971 3907 9997 3933
rect 9997 3907 9998 3933
rect 9970 3906 9998 3907
rect 10022 3933 10050 3934
rect 10022 3907 10023 3933
rect 10023 3907 10049 3933
rect 10049 3907 10050 3933
rect 10022 3906 10050 3907
rect 9918 3149 9946 3150
rect 9918 3123 9919 3149
rect 9919 3123 9945 3149
rect 9945 3123 9946 3149
rect 9918 3122 9946 3123
rect 9970 3149 9998 3150
rect 9970 3123 9971 3149
rect 9971 3123 9997 3149
rect 9997 3123 9998 3149
rect 9970 3122 9998 3123
rect 10022 3149 10050 3150
rect 10022 3123 10023 3149
rect 10023 3123 10049 3149
rect 10049 3123 10050 3149
rect 10022 3122 10050 3123
rect 9918 2365 9946 2366
rect 9918 2339 9919 2365
rect 9919 2339 9945 2365
rect 9945 2339 9946 2365
rect 9918 2338 9946 2339
rect 9970 2365 9998 2366
rect 9970 2339 9971 2365
rect 9971 2339 9997 2365
rect 9997 2339 9998 2365
rect 9970 2338 9998 2339
rect 10022 2365 10050 2366
rect 10022 2339 10023 2365
rect 10023 2339 10049 2365
rect 10049 2339 10050 2365
rect 10022 2338 10050 2339
rect 9758 2030 9786 2058
rect 10374 2057 10402 2058
rect 10374 2031 10375 2057
rect 10375 2031 10401 2057
rect 10401 2031 10402 2057
rect 10374 2030 10402 2031
rect 14574 9617 14602 9618
rect 14574 9591 14575 9617
rect 14575 9591 14601 9617
rect 14601 9591 14602 9617
rect 14574 9590 14602 9591
rect 14686 9478 14714 9506
rect 18830 10009 18858 10010
rect 18830 9983 18831 10009
rect 18831 9983 18857 10009
rect 18857 9983 18858 10009
rect 18830 9982 18858 9983
rect 15302 9534 15330 9562
rect 15078 9505 15106 9506
rect 15078 9479 15079 9505
rect 15079 9479 15105 9505
rect 15105 9479 15106 9505
rect 15078 9478 15106 9479
rect 15022 9422 15050 9450
rect 14574 9254 14602 9282
rect 17598 9813 17626 9814
rect 17598 9787 17599 9813
rect 17599 9787 17625 9813
rect 17625 9787 17626 9813
rect 17598 9786 17626 9787
rect 17650 9813 17678 9814
rect 17650 9787 17651 9813
rect 17651 9787 17677 9813
rect 17677 9787 17678 9813
rect 17650 9786 17678 9787
rect 17702 9813 17730 9814
rect 17702 9787 17703 9813
rect 17703 9787 17729 9813
rect 17729 9787 17730 9813
rect 17702 9786 17730 9787
rect 20006 9758 20034 9786
rect 18830 9617 18858 9618
rect 18830 9591 18831 9617
rect 18831 9591 18857 9617
rect 18857 9591 18858 9617
rect 18830 9590 18858 9591
rect 15470 9478 15498 9506
rect 20006 9422 20034 9450
rect 17598 9029 17626 9030
rect 17598 9003 17599 9029
rect 17599 9003 17625 9029
rect 17625 9003 17626 9029
rect 17598 9002 17626 9003
rect 17650 9029 17678 9030
rect 17650 9003 17651 9029
rect 17651 9003 17677 9029
rect 17677 9003 17678 9029
rect 17650 9002 17678 9003
rect 17702 9029 17730 9030
rect 17702 9003 17703 9029
rect 17703 9003 17729 9029
rect 17729 9003 17730 9029
rect 17702 9002 17730 9003
rect 17598 8245 17626 8246
rect 17598 8219 17599 8245
rect 17599 8219 17625 8245
rect 17625 8219 17626 8245
rect 17598 8218 17626 8219
rect 17650 8245 17678 8246
rect 17650 8219 17651 8245
rect 17651 8219 17677 8245
rect 17677 8219 17678 8245
rect 17650 8218 17678 8219
rect 17702 8245 17730 8246
rect 17702 8219 17703 8245
rect 17703 8219 17729 8245
rect 17729 8219 17730 8245
rect 17702 8218 17730 8219
rect 14070 8134 14098 8162
rect 14350 8022 14378 8050
rect 14518 8134 14546 8162
rect 14686 8049 14714 8050
rect 14686 8023 14687 8049
rect 14687 8023 14713 8049
rect 14713 8023 14714 8049
rect 14686 8022 14714 8023
rect 14910 8049 14938 8050
rect 14910 8023 14911 8049
rect 14911 8023 14937 8049
rect 14937 8023 14938 8049
rect 14910 8022 14938 8023
rect 15134 8022 15162 8050
rect 14182 7993 14210 7994
rect 14182 7967 14183 7993
rect 14183 7967 14209 7993
rect 14209 7967 14210 7993
rect 14182 7966 14210 7967
rect 14854 7993 14882 7994
rect 14854 7967 14855 7993
rect 14855 7967 14881 7993
rect 14881 7967 14882 7993
rect 14854 7966 14882 7967
rect 13342 6846 13370 6874
rect 14630 7937 14658 7938
rect 14630 7911 14631 7937
rect 14631 7911 14657 7937
rect 14657 7911 14658 7937
rect 14630 7910 14658 7911
rect 14966 7910 14994 7938
rect 15134 7769 15162 7770
rect 15134 7743 15135 7769
rect 15135 7743 15161 7769
rect 15161 7743 15162 7769
rect 15134 7742 15162 7743
rect 18830 8049 18858 8050
rect 18830 8023 18831 8049
rect 18831 8023 18857 8049
rect 18857 8023 18858 8049
rect 18830 8022 18858 8023
rect 19950 8078 19978 8106
rect 18942 7910 18970 7938
rect 20006 7742 20034 7770
rect 17598 7461 17626 7462
rect 17598 7435 17599 7461
rect 17599 7435 17625 7461
rect 17625 7435 17626 7461
rect 17598 7434 17626 7435
rect 17650 7461 17678 7462
rect 17650 7435 17651 7461
rect 17651 7435 17677 7461
rect 17677 7435 17678 7461
rect 17650 7434 17678 7435
rect 17702 7461 17730 7462
rect 17702 7435 17703 7461
rect 17703 7435 17729 7461
rect 17729 7435 17730 7461
rect 17702 7434 17730 7435
rect 17598 6677 17626 6678
rect 17598 6651 17599 6677
rect 17599 6651 17625 6677
rect 17625 6651 17626 6677
rect 17598 6650 17626 6651
rect 17650 6677 17678 6678
rect 17650 6651 17651 6677
rect 17651 6651 17677 6677
rect 17677 6651 17678 6677
rect 17650 6650 17678 6651
rect 17702 6677 17730 6678
rect 17702 6651 17703 6677
rect 17703 6651 17729 6677
rect 17729 6651 17730 6677
rect 17702 6650 17730 6651
rect 17598 5893 17626 5894
rect 17598 5867 17599 5893
rect 17599 5867 17625 5893
rect 17625 5867 17626 5893
rect 17598 5866 17626 5867
rect 17650 5893 17678 5894
rect 17650 5867 17651 5893
rect 17651 5867 17677 5893
rect 17677 5867 17678 5893
rect 17650 5866 17678 5867
rect 17702 5893 17730 5894
rect 17702 5867 17703 5893
rect 17703 5867 17729 5893
rect 17729 5867 17730 5893
rect 17702 5866 17730 5867
rect 17598 5109 17626 5110
rect 17598 5083 17599 5109
rect 17599 5083 17625 5109
rect 17625 5083 17626 5109
rect 17598 5082 17626 5083
rect 17650 5109 17678 5110
rect 17650 5083 17651 5109
rect 17651 5083 17677 5109
rect 17677 5083 17678 5109
rect 17650 5082 17678 5083
rect 17702 5109 17730 5110
rect 17702 5083 17703 5109
rect 17703 5083 17729 5109
rect 17729 5083 17730 5109
rect 17702 5082 17730 5083
rect 17598 4325 17626 4326
rect 17598 4299 17599 4325
rect 17599 4299 17625 4325
rect 17625 4299 17626 4325
rect 17598 4298 17626 4299
rect 17650 4325 17678 4326
rect 17650 4299 17651 4325
rect 17651 4299 17677 4325
rect 17677 4299 17678 4325
rect 17650 4298 17678 4299
rect 17702 4325 17730 4326
rect 17702 4299 17703 4325
rect 17703 4299 17729 4325
rect 17729 4299 17730 4325
rect 17702 4298 17730 4299
rect 12110 2030 12138 2058
rect 11438 1806 11466 1834
rect 9918 1581 9946 1582
rect 9918 1555 9919 1581
rect 9919 1555 9945 1581
rect 9945 1555 9946 1581
rect 9918 1554 9946 1555
rect 9970 1581 9998 1582
rect 9970 1555 9971 1581
rect 9971 1555 9997 1581
rect 9997 1555 9998 1581
rect 9970 1554 9998 1555
rect 10022 1581 10050 1582
rect 10022 1555 10023 1581
rect 10023 1555 10049 1581
rect 10049 1555 10050 1581
rect 10022 1554 10050 1555
rect 17598 3541 17626 3542
rect 17598 3515 17599 3541
rect 17599 3515 17625 3541
rect 17625 3515 17626 3541
rect 17598 3514 17626 3515
rect 17650 3541 17678 3542
rect 17650 3515 17651 3541
rect 17651 3515 17677 3541
rect 17677 3515 17678 3541
rect 17650 3514 17678 3515
rect 17702 3541 17730 3542
rect 17702 3515 17703 3541
rect 17703 3515 17729 3541
rect 17729 3515 17730 3541
rect 17702 3514 17730 3515
rect 17598 2757 17626 2758
rect 17598 2731 17599 2757
rect 17599 2731 17625 2757
rect 17625 2731 17626 2757
rect 17598 2730 17626 2731
rect 17650 2757 17678 2758
rect 17650 2731 17651 2757
rect 17651 2731 17677 2757
rect 17677 2731 17678 2757
rect 17650 2730 17678 2731
rect 17702 2757 17730 2758
rect 17702 2731 17703 2757
rect 17703 2731 17729 2757
rect 17729 2731 17730 2757
rect 17702 2730 17730 2731
rect 13118 2057 13146 2058
rect 13118 2031 13119 2057
rect 13119 2031 13145 2057
rect 13145 2031 13146 2057
rect 13118 2030 13146 2031
rect 17598 1973 17626 1974
rect 17598 1947 17599 1973
rect 17599 1947 17625 1973
rect 17625 1947 17626 1973
rect 17598 1946 17626 1947
rect 17650 1973 17678 1974
rect 17650 1947 17651 1973
rect 17651 1947 17677 1973
rect 17677 1947 17678 1973
rect 17650 1946 17678 1947
rect 17702 1973 17730 1974
rect 17702 1947 17703 1973
rect 17703 1947 17729 1973
rect 17729 1947 17730 1973
rect 17702 1946 17730 1947
rect 12782 1833 12810 1834
rect 12782 1807 12783 1833
rect 12783 1807 12809 1833
rect 12809 1807 12810 1833
rect 12782 1806 12810 1807
<< metal3 >>
rect 12777 19278 12782 19306
rect 12810 19278 13398 19306
rect 13426 19278 13431 19306
rect 2233 19194 2238 19222
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2370 19194 2375 19222
rect 17593 19194 17598 19222
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17730 19194 17735 19222
rect 8745 19110 8750 19138
rect 8778 19110 9310 19138
rect 9338 19110 9343 19138
rect 11433 19110 11438 19138
rect 11466 19110 12782 19138
rect 12810 19110 12815 19138
rect 13113 19110 13118 19138
rect 13146 19110 14686 19138
rect 14714 19110 14719 19138
rect 9913 18802 9918 18830
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 10050 18802 10055 18830
rect 9417 18718 9422 18746
rect 9450 18718 10038 18746
rect 10066 18718 10071 18746
rect 2233 18410 2238 18438
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2370 18410 2375 18438
rect 17593 18410 17598 18438
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17730 18410 17735 18438
rect 7737 18326 7742 18354
rect 7770 18326 8358 18354
rect 8386 18326 8391 18354
rect 9913 18018 9918 18046
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 10050 18018 10055 18046
rect 2233 17626 2238 17654
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2370 17626 2375 17654
rect 17593 17626 17598 17654
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17730 17626 17735 17654
rect 9913 17234 9918 17262
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 10050 17234 10055 17262
rect 2233 16842 2238 16870
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2370 16842 2375 16870
rect 17593 16842 17598 16870
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17730 16842 17735 16870
rect 9913 16450 9918 16478
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 10050 16450 10055 16478
rect 2233 16058 2238 16086
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2370 16058 2375 16086
rect 17593 16058 17598 16086
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17730 16058 17735 16086
rect 9913 15666 9918 15694
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 10050 15666 10055 15694
rect 2233 15274 2238 15302
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2370 15274 2375 15302
rect 17593 15274 17598 15302
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17730 15274 17735 15302
rect 9913 14882 9918 14910
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 10050 14882 10055 14910
rect 2233 14490 2238 14518
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2370 14490 2375 14518
rect 17593 14490 17598 14518
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17730 14490 17735 14518
rect 10929 14238 10934 14266
rect 10962 14238 11830 14266
rect 11858 14238 11863 14266
rect 9913 14098 9918 14126
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 10050 14098 10055 14126
rect 13113 14014 13118 14042
rect 13146 14014 14294 14042
rect 14322 14014 14327 14042
rect 10257 13902 10262 13930
rect 10290 13902 11774 13930
rect 11802 13902 11942 13930
rect 11970 13902 11975 13930
rect 6561 13846 6566 13874
rect 6594 13846 7126 13874
rect 7154 13846 7159 13874
rect 11657 13846 11662 13874
rect 11690 13846 12278 13874
rect 12306 13846 12311 13874
rect 0 13818 400 13832
rect 0 13790 2086 13818
rect 2114 13790 2119 13818
rect 11545 13790 11550 13818
rect 11578 13790 12614 13818
rect 12642 13790 12647 13818
rect 0 13776 400 13790
rect 2233 13706 2238 13734
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2370 13706 2375 13734
rect 17593 13706 17598 13734
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17730 13706 17735 13734
rect 8185 13566 8190 13594
rect 8218 13566 9198 13594
rect 9226 13566 10766 13594
rect 10794 13566 11382 13594
rect 11410 13566 11415 13594
rect 6225 13510 6230 13538
rect 6258 13510 7462 13538
rect 7490 13510 7910 13538
rect 7938 13510 7943 13538
rect 6230 13426 6258 13510
rect 10990 13482 11018 13566
rect 11769 13510 11774 13538
rect 11802 13510 12614 13538
rect 12642 13510 13398 13538
rect 13426 13510 13431 13538
rect 10985 13454 10990 13482
rect 11018 13454 11023 13482
rect 11601 13454 11606 13482
rect 11634 13454 12110 13482
rect 12138 13454 12143 13482
rect 5609 13398 5614 13426
rect 5642 13398 6258 13426
rect 10929 13398 10934 13426
rect 10962 13398 11326 13426
rect 11354 13398 11774 13426
rect 11802 13398 11807 13426
rect 9913 13314 9918 13342
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 10050 13314 10055 13342
rect 13393 13230 13398 13258
rect 13426 13230 13678 13258
rect 13706 13230 14294 13258
rect 14322 13230 14327 13258
rect 7177 13174 7182 13202
rect 7210 13174 8078 13202
rect 8106 13174 8111 13202
rect 11153 13174 11158 13202
rect 11186 13174 12110 13202
rect 12138 13174 12143 13202
rect 20600 13146 21000 13160
rect 8409 13118 8414 13146
rect 8442 13118 9086 13146
rect 9114 13118 9119 13146
rect 11097 13118 11102 13146
rect 11130 13118 11270 13146
rect 11298 13118 11303 13146
rect 13281 13118 13286 13146
rect 13314 13118 14070 13146
rect 14098 13118 18830 13146
rect 18858 13118 18863 13146
rect 20001 13118 20006 13146
rect 20034 13118 21000 13146
rect 20600 13104 21000 13118
rect 2137 13062 2142 13090
rect 2170 13062 7014 13090
rect 7042 13062 7798 13090
rect 7826 13062 7831 13090
rect 7905 13062 7910 13090
rect 7938 13062 8582 13090
rect 8610 13062 8918 13090
rect 8946 13062 8951 13090
rect 12273 13062 12278 13090
rect 12306 13062 13006 13090
rect 13034 13062 13039 13090
rect 7910 13034 7938 13062
rect 7569 13006 7574 13034
rect 7602 13006 7938 13034
rect 7513 12950 7518 12978
rect 7546 12950 7742 12978
rect 7770 12950 8750 12978
rect 8778 12950 8783 12978
rect 2233 12922 2238 12950
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2370 12922 2375 12950
rect 17593 12922 17598 12950
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17730 12922 17735 12950
rect 9025 12838 9030 12866
rect 9058 12838 9534 12866
rect 9562 12838 10654 12866
rect 10682 12838 10687 12866
rect 0 12810 400 12824
rect 0 12782 966 12810
rect 994 12782 999 12810
rect 10817 12782 10822 12810
rect 10850 12782 11158 12810
rect 11186 12782 11191 12810
rect 0 12768 400 12782
rect 10593 12726 10598 12754
rect 10626 12726 10878 12754
rect 10906 12726 10911 12754
rect 12329 12726 12334 12754
rect 12362 12726 13174 12754
rect 13202 12726 13207 12754
rect 6393 12670 6398 12698
rect 6426 12670 7294 12698
rect 7322 12670 7327 12698
rect 8633 12670 8638 12698
rect 8666 12670 9030 12698
rect 9058 12670 9063 12698
rect 7233 12614 7238 12642
rect 7266 12614 7686 12642
rect 7714 12614 8246 12642
rect 8274 12614 9422 12642
rect 9450 12614 9926 12642
rect 9954 12614 9959 12642
rect 9913 12530 9918 12558
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 10050 12530 10055 12558
rect 7457 12446 7462 12474
rect 7490 12446 7574 12474
rect 7602 12446 7607 12474
rect 9137 12446 9142 12474
rect 9170 12446 10262 12474
rect 10290 12446 10710 12474
rect 10738 12446 10743 12474
rect 15946 12334 18830 12362
rect 18858 12334 18863 12362
rect 15946 12306 15974 12334
rect 13281 12278 13286 12306
rect 13314 12278 14238 12306
rect 14266 12278 14271 12306
rect 15297 12278 15302 12306
rect 15330 12278 15974 12306
rect 2233 12138 2238 12166
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2370 12138 2375 12166
rect 17593 12138 17598 12166
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17730 12138 17735 12166
rect 20600 12138 21000 12152
rect 20001 12110 20006 12138
rect 20034 12110 21000 12138
rect 20600 12096 21000 12110
rect 2137 11942 2142 11970
rect 2170 11942 5558 11970
rect 5586 11942 7014 11970
rect 7042 11942 7047 11970
rect 10537 11942 10542 11970
rect 10570 11942 11942 11970
rect 11970 11942 11975 11970
rect 13953 11942 13958 11970
rect 13986 11942 15302 11970
rect 15330 11942 15335 11970
rect 10761 11886 10766 11914
rect 10794 11886 11046 11914
rect 11074 11886 11079 11914
rect 13561 11830 13566 11858
rect 13594 11830 13902 11858
rect 13930 11830 13935 11858
rect 0 11802 400 11816
rect 20600 11802 21000 11816
rect 0 11774 966 11802
rect 994 11774 999 11802
rect 20001 11774 20006 11802
rect 20034 11774 21000 11802
rect 0 11760 400 11774
rect 9913 11746 9918 11774
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 10050 11746 10055 11774
rect 20600 11760 21000 11774
rect 9025 11718 9030 11746
rect 9058 11718 9758 11746
rect 9786 11718 9791 11746
rect 15946 11718 18830 11746
rect 18858 11718 18863 11746
rect 9305 11662 9310 11690
rect 9338 11662 13342 11690
rect 13370 11662 14070 11690
rect 14098 11662 14103 11690
rect 15946 11634 15974 11718
rect 10929 11606 10934 11634
rect 10962 11606 11998 11634
rect 12026 11606 12894 11634
rect 12922 11606 13846 11634
rect 13874 11606 13879 11634
rect 15409 11606 15414 11634
rect 15442 11606 15974 11634
rect 2137 11550 2142 11578
rect 2170 11550 6062 11578
rect 6090 11550 7798 11578
rect 7826 11550 7831 11578
rect 9473 11550 9478 11578
rect 9506 11550 10150 11578
rect 10178 11550 10710 11578
rect 10738 11550 10743 11578
rect 10873 11550 10878 11578
rect 10906 11550 11382 11578
rect 11410 11550 11415 11578
rect 15241 11550 15246 11578
rect 15274 11550 18830 11578
rect 18858 11550 18863 11578
rect 11153 11494 11158 11522
rect 11186 11494 11606 11522
rect 11634 11494 11639 11522
rect 0 11466 400 11480
rect 20600 11466 21000 11480
rect 0 11438 966 11466
rect 994 11438 999 11466
rect 7681 11438 7686 11466
rect 7714 11438 8582 11466
rect 8610 11438 8615 11466
rect 20001 11438 20006 11466
rect 20034 11438 21000 11466
rect 0 11424 400 11438
rect 20600 11424 21000 11438
rect 2233 11354 2238 11382
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2370 11354 2375 11382
rect 17593 11354 17598 11382
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17730 11354 17735 11382
rect 6953 11326 6958 11354
rect 6986 11326 9590 11354
rect 9618 11326 9623 11354
rect 10369 11326 10374 11354
rect 10402 11326 10990 11354
rect 11018 11326 11774 11354
rect 11802 11326 11807 11354
rect 9641 11270 9646 11298
rect 9674 11270 11746 11298
rect 7849 11214 7854 11242
rect 7882 11214 8638 11242
rect 8666 11214 8671 11242
rect 9193 11214 9198 11242
rect 9226 11214 11046 11242
rect 11074 11214 11079 11242
rect 11718 11186 11746 11270
rect 8745 11158 8750 11186
rect 8778 11158 9478 11186
rect 9506 11158 9511 11186
rect 11713 11158 11718 11186
rect 11746 11158 13790 11186
rect 13818 11158 13823 11186
rect 14009 11158 14014 11186
rect 14042 11158 14238 11186
rect 14266 11158 14271 11186
rect 7513 11102 7518 11130
rect 7546 11102 10878 11130
rect 10906 11102 10911 11130
rect 14177 11102 14182 11130
rect 14210 11102 15078 11130
rect 15106 11102 15111 11130
rect 7065 11046 7070 11074
rect 7098 11046 7630 11074
rect 7658 11046 8246 11074
rect 8274 11046 8279 11074
rect 10369 11046 10374 11074
rect 10402 11046 10654 11074
rect 10682 11046 13566 11074
rect 13594 11046 13599 11074
rect 9913 10962 9918 10990
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 10050 10962 10055 10990
rect 8353 10934 8358 10962
rect 8386 10934 8750 10962
rect 8778 10934 8783 10962
rect 9417 10934 9422 10962
rect 9450 10934 9758 10962
rect 9786 10934 9791 10962
rect 7961 10878 7966 10906
rect 7994 10878 8582 10906
rect 8610 10878 8615 10906
rect 10313 10878 10318 10906
rect 10346 10878 10486 10906
rect 10514 10878 10878 10906
rect 10906 10878 11998 10906
rect 12026 10878 12031 10906
rect 12105 10878 12110 10906
rect 12138 10878 13734 10906
rect 13762 10878 13767 10906
rect 8409 10822 8414 10850
rect 8442 10822 8862 10850
rect 8890 10822 9366 10850
rect 9394 10822 10626 10850
rect 13057 10822 13062 10850
rect 13090 10822 13510 10850
rect 13538 10822 13543 10850
rect 10598 10794 10626 10822
rect 9081 10766 9086 10794
rect 9114 10766 9758 10794
rect 9786 10766 10514 10794
rect 10593 10766 10598 10794
rect 10626 10766 10631 10794
rect 11097 10766 11102 10794
rect 11130 10766 12334 10794
rect 12362 10766 12726 10794
rect 12754 10766 13286 10794
rect 13314 10766 13319 10794
rect 10486 10738 10514 10766
rect 10486 10710 11662 10738
rect 11690 10710 12782 10738
rect 12810 10710 13118 10738
rect 13146 10710 13151 10738
rect 9865 10654 9870 10682
rect 9898 10654 11270 10682
rect 11298 10654 11303 10682
rect 2233 10570 2238 10598
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2370 10570 2375 10598
rect 17593 10570 17598 10598
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17730 10570 17735 10598
rect 7345 10430 7350 10458
rect 7378 10430 7518 10458
rect 7546 10430 7854 10458
rect 7882 10430 7887 10458
rect 10313 10430 10318 10458
rect 10346 10430 11158 10458
rect 11186 10430 11494 10458
rect 11522 10430 11527 10458
rect 13505 10430 13510 10458
rect 13538 10430 13734 10458
rect 13762 10430 13767 10458
rect 6001 10374 6006 10402
rect 6034 10374 7070 10402
rect 7098 10374 9366 10402
rect 9394 10374 9399 10402
rect 11265 10374 11270 10402
rect 11298 10374 13342 10402
rect 13370 10374 13375 10402
rect 10033 10318 10038 10346
rect 10066 10318 11046 10346
rect 11074 10318 11079 10346
rect 9913 10178 9918 10206
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 10050 10178 10055 10206
rect 9361 10094 9366 10122
rect 9394 10094 11214 10122
rect 11242 10094 11247 10122
rect 11657 10094 11662 10122
rect 11690 10094 11802 10122
rect 11774 10066 11802 10094
rect 7401 10038 7406 10066
rect 7434 10038 7910 10066
rect 7938 10038 7943 10066
rect 8185 10038 8190 10066
rect 8218 10038 10094 10066
rect 10122 10038 10127 10066
rect 11041 10038 11046 10066
rect 11074 10038 11802 10066
rect 13393 10038 13398 10066
rect 13426 10038 14294 10066
rect 14322 10038 14327 10066
rect 7065 9982 7070 10010
rect 7098 9982 7574 10010
rect 7602 9982 8022 10010
rect 8050 9982 8055 10010
rect 9081 9982 9086 10010
rect 9114 9982 10374 10010
rect 10402 9982 10407 10010
rect 15297 9982 15302 10010
rect 15330 9982 18830 10010
rect 18858 9982 18863 10010
rect 2081 9926 2086 9954
rect 2114 9926 8750 9954
rect 8778 9926 9702 9954
rect 9730 9926 9735 9954
rect 9249 9870 9254 9898
rect 9282 9870 9534 9898
rect 9562 9870 9567 9898
rect 7737 9814 7742 9842
rect 7770 9814 8414 9842
rect 8442 9814 9142 9842
rect 9170 9814 9175 9842
rect 2233 9786 2238 9814
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2370 9786 2375 9814
rect 17593 9786 17598 9814
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17730 9786 17735 9814
rect 20600 9786 21000 9800
rect 9865 9758 9870 9786
rect 9898 9758 13062 9786
rect 13090 9758 13095 9786
rect 20001 9758 20006 9786
rect 20034 9758 21000 9786
rect 20600 9744 21000 9758
rect 10033 9702 10038 9730
rect 10066 9702 10710 9730
rect 10738 9702 10743 9730
rect 13281 9702 13286 9730
rect 13314 9702 13622 9730
rect 13650 9702 13655 9730
rect 8521 9590 8526 9618
rect 8554 9590 8750 9618
rect 8778 9590 8783 9618
rect 8969 9590 8974 9618
rect 9002 9590 11382 9618
rect 11410 9590 12950 9618
rect 12978 9590 13174 9618
rect 13202 9590 13207 9618
rect 13449 9590 13454 9618
rect 13482 9590 14574 9618
rect 14602 9590 14607 9618
rect 15946 9590 18830 9618
rect 18858 9590 18863 9618
rect 7905 9534 7910 9562
rect 7938 9534 9254 9562
rect 9282 9534 10654 9562
rect 10682 9534 10687 9562
rect 13337 9534 13342 9562
rect 13370 9534 14070 9562
rect 14098 9534 14103 9562
rect 14177 9534 14182 9562
rect 14210 9534 15302 9562
rect 15330 9534 15335 9562
rect 14070 9506 14098 9534
rect 15946 9506 15974 9590
rect 8689 9478 8694 9506
rect 8722 9478 8974 9506
rect 9002 9478 9478 9506
rect 9506 9478 9511 9506
rect 11993 9478 11998 9506
rect 12026 9478 12838 9506
rect 12866 9478 12871 9506
rect 13449 9478 13454 9506
rect 13482 9478 13958 9506
rect 13986 9478 13991 9506
rect 14070 9478 14686 9506
rect 14714 9478 14719 9506
rect 15073 9478 15078 9506
rect 15106 9478 15470 9506
rect 15498 9478 15974 9506
rect 12838 9450 12866 9478
rect 20600 9450 21000 9464
rect 7961 9422 7966 9450
rect 7994 9422 8862 9450
rect 8890 9422 8895 9450
rect 12838 9422 13678 9450
rect 13706 9422 13711 9450
rect 14345 9422 14350 9450
rect 14378 9422 15022 9450
rect 15050 9422 15055 9450
rect 20001 9422 20006 9450
rect 20034 9422 21000 9450
rect 9913 9394 9918 9422
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 10050 9394 10055 9422
rect 20600 9408 21000 9422
rect 10094 9366 11830 9394
rect 11858 9366 12222 9394
rect 12250 9366 12255 9394
rect 10094 9338 10122 9366
rect 8913 9310 8918 9338
rect 8946 9310 9310 9338
rect 9338 9310 10122 9338
rect 10201 9310 10206 9338
rect 10234 9310 10430 9338
rect 10458 9310 10990 9338
rect 11018 9310 11023 9338
rect 10206 9226 10234 9310
rect 11433 9254 11438 9282
rect 11466 9254 11662 9282
rect 11690 9254 13454 9282
rect 13482 9254 13487 9282
rect 14177 9254 14182 9282
rect 14210 9254 14574 9282
rect 14602 9254 14607 9282
rect 5553 9198 5558 9226
rect 5586 9198 7182 9226
rect 7210 9198 7215 9226
rect 8745 9198 8750 9226
rect 8778 9198 9758 9226
rect 9786 9198 9791 9226
rect 9865 9198 9870 9226
rect 9898 9198 10234 9226
rect 8185 9142 8190 9170
rect 8218 9142 9646 9170
rect 9674 9142 9982 9170
rect 10010 9142 10015 9170
rect 10649 9142 10654 9170
rect 10682 9142 10934 9170
rect 10962 9142 10967 9170
rect 11601 9142 11606 9170
rect 11634 9142 12502 9170
rect 12530 9142 12535 9170
rect 9585 9086 9590 9114
rect 9618 9086 10094 9114
rect 10122 9086 11886 9114
rect 11914 9086 11919 9114
rect 11153 9030 11158 9058
rect 11186 9030 11942 9058
rect 11970 9030 11975 9058
rect 2233 9002 2238 9030
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2370 9002 2375 9030
rect 11438 8890 11466 9030
rect 17593 9002 17598 9030
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17730 9002 17735 9030
rect 11433 8862 11438 8890
rect 11466 8862 11471 8890
rect 9193 8750 9198 8778
rect 9226 8750 9702 8778
rect 9730 8750 9735 8778
rect 8297 8694 8302 8722
rect 8330 8694 8918 8722
rect 8946 8694 8951 8722
rect 12889 8694 12894 8722
rect 12922 8694 13118 8722
rect 13146 8694 13454 8722
rect 13482 8694 13678 8722
rect 13706 8694 13711 8722
rect 9913 8610 9918 8638
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 10050 8610 10055 8638
rect 10654 8582 11326 8610
rect 11354 8582 11359 8610
rect 10654 8554 10682 8582
rect 7009 8526 7014 8554
rect 7042 8526 7630 8554
rect 7658 8526 8190 8554
rect 8218 8526 8223 8554
rect 9305 8526 9310 8554
rect 9338 8526 10654 8554
rect 10682 8526 10687 8554
rect 10873 8526 10878 8554
rect 10906 8526 11102 8554
rect 11130 8526 11718 8554
rect 11746 8526 11751 8554
rect 9137 8470 9142 8498
rect 9170 8470 9534 8498
rect 9562 8470 9567 8498
rect 10878 8442 10906 8526
rect 7401 8414 7406 8442
rect 7434 8414 8974 8442
rect 9002 8414 9007 8442
rect 9697 8414 9702 8442
rect 9730 8414 10906 8442
rect 11433 8358 11438 8386
rect 11466 8358 13846 8386
rect 13874 8358 13879 8386
rect 9249 8302 9254 8330
rect 9282 8302 9590 8330
rect 9618 8302 9623 8330
rect 11825 8302 11830 8330
rect 11858 8302 12110 8330
rect 12138 8302 12143 8330
rect 9361 8246 9366 8274
rect 9394 8246 10262 8274
rect 10290 8246 11438 8274
rect 11466 8246 11471 8274
rect 2233 8218 2238 8246
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2370 8218 2375 8246
rect 17593 8218 17598 8246
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17730 8218 17735 8246
rect 2137 8134 2142 8162
rect 2170 8134 5670 8162
rect 5698 8134 5703 8162
rect 14065 8134 14070 8162
rect 14098 8134 14518 8162
rect 14546 8134 14551 8162
rect 0 8106 400 8120
rect 20600 8106 21000 8120
rect 0 8078 966 8106
rect 994 8078 999 8106
rect 7065 8078 7070 8106
rect 7098 8078 7518 8106
rect 7546 8078 7551 8106
rect 8409 8078 8414 8106
rect 8442 8078 9422 8106
rect 9450 8078 9455 8106
rect 19945 8078 19950 8106
rect 19978 8078 21000 8106
rect 0 8064 400 8078
rect 20600 8064 21000 8078
rect 2137 8022 2142 8050
rect 2170 8022 5614 8050
rect 5642 8022 5647 8050
rect 5889 8022 5894 8050
rect 5922 8022 6902 8050
rect 6930 8022 10094 8050
rect 10122 8022 10710 8050
rect 10738 8022 10743 8050
rect 14345 8022 14350 8050
rect 14378 8022 14686 8050
rect 14714 8022 14719 8050
rect 14905 8022 14910 8050
rect 14938 8022 15134 8050
rect 15162 8022 18830 8050
rect 18858 8022 18863 8050
rect 9814 7966 11046 7994
rect 11074 7966 11079 7994
rect 14177 7966 14182 7994
rect 14210 7966 14854 7994
rect 14882 7966 14887 7994
rect 9025 7910 9030 7938
rect 9058 7910 9478 7938
rect 9506 7910 9511 7938
rect 9814 7826 9842 7966
rect 14625 7910 14630 7938
rect 14658 7910 14966 7938
rect 14994 7910 18942 7938
rect 18970 7910 18975 7938
rect 9913 7826 9918 7854
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 10050 7826 10055 7854
rect 5609 7798 5614 7826
rect 5642 7798 6902 7826
rect 6930 7798 6935 7826
rect 8857 7798 8862 7826
rect 8890 7798 9478 7826
rect 9506 7798 9842 7826
rect 0 7770 400 7784
rect 20600 7770 21000 7784
rect 0 7742 1022 7770
rect 1050 7742 1055 7770
rect 5665 7742 5670 7770
rect 5698 7742 7294 7770
rect 7322 7742 7327 7770
rect 7513 7742 7518 7770
rect 7546 7742 10318 7770
rect 10346 7742 11214 7770
rect 11242 7742 11247 7770
rect 13449 7742 13454 7770
rect 13482 7742 15134 7770
rect 15162 7742 15167 7770
rect 20001 7742 20006 7770
rect 20034 7742 21000 7770
rect 0 7728 400 7742
rect 20600 7728 21000 7742
rect 6785 7686 6790 7714
rect 6818 7686 7462 7714
rect 7490 7686 7495 7714
rect 9137 7686 9142 7714
rect 9170 7686 11998 7714
rect 12026 7686 12031 7714
rect 7345 7630 7350 7658
rect 7378 7630 8918 7658
rect 8946 7630 8951 7658
rect 9697 7630 9702 7658
rect 9730 7630 10738 7658
rect 10817 7630 10822 7658
rect 10850 7630 11046 7658
rect 11074 7630 11079 7658
rect 11214 7630 11830 7658
rect 11858 7630 11863 7658
rect 12049 7630 12054 7658
rect 12082 7630 13118 7658
rect 13146 7630 13151 7658
rect 7177 7574 7182 7602
rect 7210 7574 7518 7602
rect 7546 7574 7551 7602
rect 7737 7574 7742 7602
rect 7770 7574 8722 7602
rect 9081 7574 9086 7602
rect 9114 7574 9646 7602
rect 9674 7574 9679 7602
rect 9758 7574 10486 7602
rect 10514 7574 10519 7602
rect 8694 7546 8722 7574
rect 9758 7546 9786 7574
rect 10710 7546 10738 7630
rect 11214 7602 11242 7630
rect 10934 7574 11242 7602
rect 11321 7574 11326 7602
rect 11354 7574 12334 7602
rect 12362 7574 12367 7602
rect 10934 7546 10962 7574
rect 7009 7518 7014 7546
rect 7042 7518 7406 7546
rect 7434 7518 8470 7546
rect 8498 7518 8503 7546
rect 8689 7518 8694 7546
rect 8722 7518 8727 7546
rect 9753 7518 9758 7546
rect 9786 7518 9791 7546
rect 10710 7518 10934 7546
rect 10962 7518 10967 7546
rect 2233 7434 2238 7462
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2370 7434 2375 7462
rect 17593 7434 17598 7462
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17730 7434 17735 7462
rect 8969 7126 8974 7154
rect 9002 7126 9590 7154
rect 9618 7126 9623 7154
rect 9913 7042 9918 7070
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 10050 7042 10055 7070
rect 8913 6958 8918 6986
rect 8946 6958 9254 6986
rect 9282 6958 9758 6986
rect 9786 6958 10094 6986
rect 10066 6818 10094 6958
rect 10929 6846 10934 6874
rect 10962 6846 11662 6874
rect 11690 6846 12670 6874
rect 12698 6846 13342 6874
rect 13370 6846 13375 6874
rect 10066 6790 10206 6818
rect 10234 6790 10239 6818
rect 2233 6650 2238 6678
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2370 6650 2375 6678
rect 17593 6650 17598 6678
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17730 6650 17735 6678
rect 9913 6258 9918 6286
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 10050 6258 10055 6286
rect 2233 5866 2238 5894
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2370 5866 2375 5894
rect 17593 5866 17598 5894
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17730 5866 17735 5894
rect 8465 5838 8470 5866
rect 8498 5838 8862 5866
rect 8890 5838 8895 5866
rect 9913 5474 9918 5502
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 10050 5474 10055 5502
rect 2233 5082 2238 5110
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2370 5082 2375 5110
rect 17593 5082 17598 5110
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17730 5082 17735 5110
rect 9913 4690 9918 4718
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 10050 4690 10055 4718
rect 2233 4298 2238 4326
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2370 4298 2375 4326
rect 17593 4298 17598 4326
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17730 4298 17735 4326
rect 9913 3906 9918 3934
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 10050 3906 10055 3934
rect 2233 3514 2238 3542
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2370 3514 2375 3542
rect 17593 3514 17598 3542
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17730 3514 17735 3542
rect 9913 3122 9918 3150
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 10050 3122 10055 3150
rect 2233 2730 2238 2758
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2370 2730 2375 2758
rect 17593 2730 17598 2758
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17730 2730 17735 2758
rect 8745 2590 8750 2618
rect 8778 2590 9366 2618
rect 9394 2590 9399 2618
rect 9913 2338 9918 2366
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 10050 2338 10055 2366
rect 9753 2030 9758 2058
rect 9786 2030 10374 2058
rect 10402 2030 10407 2058
rect 12105 2030 12110 2058
rect 12138 2030 13118 2058
rect 13146 2030 13151 2058
rect 2233 1946 2238 1974
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2370 1946 2375 1974
rect 17593 1946 17598 1974
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17730 1946 17735 1974
rect 11433 1806 11438 1834
rect 11466 1806 12782 1834
rect 12810 1806 12815 1834
rect 9913 1554 9918 1582
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 10050 1554 10055 1582
<< via3 >>
rect 2238 19194 2266 19222
rect 2290 19194 2318 19222
rect 2342 19194 2370 19222
rect 17598 19194 17626 19222
rect 17650 19194 17678 19222
rect 17702 19194 17730 19222
rect 9918 18802 9946 18830
rect 9970 18802 9998 18830
rect 10022 18802 10050 18830
rect 2238 18410 2266 18438
rect 2290 18410 2318 18438
rect 2342 18410 2370 18438
rect 17598 18410 17626 18438
rect 17650 18410 17678 18438
rect 17702 18410 17730 18438
rect 9918 18018 9946 18046
rect 9970 18018 9998 18046
rect 10022 18018 10050 18046
rect 2238 17626 2266 17654
rect 2290 17626 2318 17654
rect 2342 17626 2370 17654
rect 17598 17626 17626 17654
rect 17650 17626 17678 17654
rect 17702 17626 17730 17654
rect 9918 17234 9946 17262
rect 9970 17234 9998 17262
rect 10022 17234 10050 17262
rect 2238 16842 2266 16870
rect 2290 16842 2318 16870
rect 2342 16842 2370 16870
rect 17598 16842 17626 16870
rect 17650 16842 17678 16870
rect 17702 16842 17730 16870
rect 9918 16450 9946 16478
rect 9970 16450 9998 16478
rect 10022 16450 10050 16478
rect 2238 16058 2266 16086
rect 2290 16058 2318 16086
rect 2342 16058 2370 16086
rect 17598 16058 17626 16086
rect 17650 16058 17678 16086
rect 17702 16058 17730 16086
rect 9918 15666 9946 15694
rect 9970 15666 9998 15694
rect 10022 15666 10050 15694
rect 2238 15274 2266 15302
rect 2290 15274 2318 15302
rect 2342 15274 2370 15302
rect 17598 15274 17626 15302
rect 17650 15274 17678 15302
rect 17702 15274 17730 15302
rect 9918 14882 9946 14910
rect 9970 14882 9998 14910
rect 10022 14882 10050 14910
rect 2238 14490 2266 14518
rect 2290 14490 2318 14518
rect 2342 14490 2370 14518
rect 17598 14490 17626 14518
rect 17650 14490 17678 14518
rect 17702 14490 17730 14518
rect 9918 14098 9946 14126
rect 9970 14098 9998 14126
rect 10022 14098 10050 14126
rect 2238 13706 2266 13734
rect 2290 13706 2318 13734
rect 2342 13706 2370 13734
rect 17598 13706 17626 13734
rect 17650 13706 17678 13734
rect 17702 13706 17730 13734
rect 9918 13314 9946 13342
rect 9970 13314 9998 13342
rect 10022 13314 10050 13342
rect 2238 12922 2266 12950
rect 2290 12922 2318 12950
rect 2342 12922 2370 12950
rect 17598 12922 17626 12950
rect 17650 12922 17678 12950
rect 17702 12922 17730 12950
rect 9918 12530 9946 12558
rect 9970 12530 9998 12558
rect 10022 12530 10050 12558
rect 2238 12138 2266 12166
rect 2290 12138 2318 12166
rect 2342 12138 2370 12166
rect 17598 12138 17626 12166
rect 17650 12138 17678 12166
rect 17702 12138 17730 12166
rect 9918 11746 9946 11774
rect 9970 11746 9998 11774
rect 10022 11746 10050 11774
rect 2238 11354 2266 11382
rect 2290 11354 2318 11382
rect 2342 11354 2370 11382
rect 17598 11354 17626 11382
rect 17650 11354 17678 11382
rect 17702 11354 17730 11382
rect 9918 10962 9946 10990
rect 9970 10962 9998 10990
rect 10022 10962 10050 10990
rect 2238 10570 2266 10598
rect 2290 10570 2318 10598
rect 2342 10570 2370 10598
rect 17598 10570 17626 10598
rect 17650 10570 17678 10598
rect 17702 10570 17730 10598
rect 9918 10178 9946 10206
rect 9970 10178 9998 10206
rect 10022 10178 10050 10206
rect 2238 9786 2266 9814
rect 2290 9786 2318 9814
rect 2342 9786 2370 9814
rect 17598 9786 17626 9814
rect 17650 9786 17678 9814
rect 17702 9786 17730 9814
rect 9918 9394 9946 9422
rect 9970 9394 9998 9422
rect 10022 9394 10050 9422
rect 2238 9002 2266 9030
rect 2290 9002 2318 9030
rect 2342 9002 2370 9030
rect 17598 9002 17626 9030
rect 17650 9002 17678 9030
rect 17702 9002 17730 9030
rect 9918 8610 9946 8638
rect 9970 8610 9998 8638
rect 10022 8610 10050 8638
rect 2238 8218 2266 8246
rect 2290 8218 2318 8246
rect 2342 8218 2370 8246
rect 17598 8218 17626 8246
rect 17650 8218 17678 8246
rect 17702 8218 17730 8246
rect 9918 7826 9946 7854
rect 9970 7826 9998 7854
rect 10022 7826 10050 7854
rect 2238 7434 2266 7462
rect 2290 7434 2318 7462
rect 2342 7434 2370 7462
rect 17598 7434 17626 7462
rect 17650 7434 17678 7462
rect 17702 7434 17730 7462
rect 9918 7042 9946 7070
rect 9970 7042 9998 7070
rect 10022 7042 10050 7070
rect 2238 6650 2266 6678
rect 2290 6650 2318 6678
rect 2342 6650 2370 6678
rect 17598 6650 17626 6678
rect 17650 6650 17678 6678
rect 17702 6650 17730 6678
rect 9918 6258 9946 6286
rect 9970 6258 9998 6286
rect 10022 6258 10050 6286
rect 2238 5866 2266 5894
rect 2290 5866 2318 5894
rect 2342 5866 2370 5894
rect 17598 5866 17626 5894
rect 17650 5866 17678 5894
rect 17702 5866 17730 5894
rect 9918 5474 9946 5502
rect 9970 5474 9998 5502
rect 10022 5474 10050 5502
rect 2238 5082 2266 5110
rect 2290 5082 2318 5110
rect 2342 5082 2370 5110
rect 17598 5082 17626 5110
rect 17650 5082 17678 5110
rect 17702 5082 17730 5110
rect 9918 4690 9946 4718
rect 9970 4690 9998 4718
rect 10022 4690 10050 4718
rect 2238 4298 2266 4326
rect 2290 4298 2318 4326
rect 2342 4298 2370 4326
rect 17598 4298 17626 4326
rect 17650 4298 17678 4326
rect 17702 4298 17730 4326
rect 9918 3906 9946 3934
rect 9970 3906 9998 3934
rect 10022 3906 10050 3934
rect 2238 3514 2266 3542
rect 2290 3514 2318 3542
rect 2342 3514 2370 3542
rect 17598 3514 17626 3542
rect 17650 3514 17678 3542
rect 17702 3514 17730 3542
rect 9918 3122 9946 3150
rect 9970 3122 9998 3150
rect 10022 3122 10050 3150
rect 2238 2730 2266 2758
rect 2290 2730 2318 2758
rect 2342 2730 2370 2758
rect 17598 2730 17626 2758
rect 17650 2730 17678 2758
rect 17702 2730 17730 2758
rect 9918 2338 9946 2366
rect 9970 2338 9998 2366
rect 10022 2338 10050 2366
rect 2238 1946 2266 1974
rect 2290 1946 2318 1974
rect 2342 1946 2370 1974
rect 17598 1946 17626 1974
rect 17650 1946 17678 1974
rect 17702 1946 17730 1974
rect 9918 1554 9946 1582
rect 9970 1554 9998 1582
rect 10022 1554 10050 1582
<< metal4 >>
rect 2224 19222 2384 19238
rect 2224 19194 2238 19222
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2370 19194 2384 19222
rect 2224 18438 2384 19194
rect 2224 18410 2238 18438
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2370 18410 2384 18438
rect 2224 17654 2384 18410
rect 2224 17626 2238 17654
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2370 17626 2384 17654
rect 2224 16870 2384 17626
rect 2224 16842 2238 16870
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2370 16842 2384 16870
rect 2224 16086 2384 16842
rect 2224 16058 2238 16086
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2370 16058 2384 16086
rect 2224 15302 2384 16058
rect 2224 15274 2238 15302
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2370 15274 2384 15302
rect 2224 14518 2384 15274
rect 2224 14490 2238 14518
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2370 14490 2384 14518
rect 2224 13734 2384 14490
rect 2224 13706 2238 13734
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2370 13706 2384 13734
rect 2224 12950 2384 13706
rect 2224 12922 2238 12950
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2370 12922 2384 12950
rect 2224 12166 2384 12922
rect 2224 12138 2238 12166
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2370 12138 2384 12166
rect 2224 11382 2384 12138
rect 2224 11354 2238 11382
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2370 11354 2384 11382
rect 2224 10598 2384 11354
rect 2224 10570 2238 10598
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2370 10570 2384 10598
rect 2224 9814 2384 10570
rect 2224 9786 2238 9814
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2370 9786 2384 9814
rect 2224 9030 2384 9786
rect 2224 9002 2238 9030
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2370 9002 2384 9030
rect 2224 8246 2384 9002
rect 2224 8218 2238 8246
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2370 8218 2384 8246
rect 2224 7462 2384 8218
rect 2224 7434 2238 7462
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2370 7434 2384 7462
rect 2224 6678 2384 7434
rect 2224 6650 2238 6678
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2370 6650 2384 6678
rect 2224 5894 2384 6650
rect 2224 5866 2238 5894
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2370 5866 2384 5894
rect 2224 5110 2384 5866
rect 2224 5082 2238 5110
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2370 5082 2384 5110
rect 2224 4326 2384 5082
rect 2224 4298 2238 4326
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2370 4298 2384 4326
rect 2224 3542 2384 4298
rect 2224 3514 2238 3542
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2370 3514 2384 3542
rect 2224 2758 2384 3514
rect 2224 2730 2238 2758
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2370 2730 2384 2758
rect 2224 1974 2384 2730
rect 2224 1946 2238 1974
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2370 1946 2384 1974
rect 2224 1538 2384 1946
rect 9904 18830 10064 19238
rect 9904 18802 9918 18830
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 10050 18802 10064 18830
rect 9904 18046 10064 18802
rect 9904 18018 9918 18046
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 10050 18018 10064 18046
rect 9904 17262 10064 18018
rect 9904 17234 9918 17262
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 10050 17234 10064 17262
rect 9904 16478 10064 17234
rect 9904 16450 9918 16478
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 10050 16450 10064 16478
rect 9904 15694 10064 16450
rect 9904 15666 9918 15694
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 10050 15666 10064 15694
rect 9904 14910 10064 15666
rect 9904 14882 9918 14910
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 10050 14882 10064 14910
rect 9904 14126 10064 14882
rect 9904 14098 9918 14126
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 10050 14098 10064 14126
rect 9904 13342 10064 14098
rect 9904 13314 9918 13342
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 10050 13314 10064 13342
rect 9904 12558 10064 13314
rect 9904 12530 9918 12558
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 10050 12530 10064 12558
rect 9904 11774 10064 12530
rect 9904 11746 9918 11774
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 10050 11746 10064 11774
rect 9904 10990 10064 11746
rect 9904 10962 9918 10990
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 10050 10962 10064 10990
rect 9904 10206 10064 10962
rect 9904 10178 9918 10206
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 10050 10178 10064 10206
rect 9904 9422 10064 10178
rect 9904 9394 9918 9422
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 10050 9394 10064 9422
rect 9904 8638 10064 9394
rect 9904 8610 9918 8638
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 10050 8610 10064 8638
rect 9904 7854 10064 8610
rect 9904 7826 9918 7854
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 10050 7826 10064 7854
rect 9904 7070 10064 7826
rect 9904 7042 9918 7070
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 10050 7042 10064 7070
rect 9904 6286 10064 7042
rect 9904 6258 9918 6286
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 10050 6258 10064 6286
rect 9904 5502 10064 6258
rect 9904 5474 9918 5502
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 10050 5474 10064 5502
rect 9904 4718 10064 5474
rect 9904 4690 9918 4718
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 10050 4690 10064 4718
rect 9904 3934 10064 4690
rect 9904 3906 9918 3934
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 10050 3906 10064 3934
rect 9904 3150 10064 3906
rect 9904 3122 9918 3150
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 10050 3122 10064 3150
rect 9904 2366 10064 3122
rect 9904 2338 9918 2366
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 10050 2338 10064 2366
rect 9904 1582 10064 2338
rect 9904 1554 9918 1582
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 10050 1554 10064 1582
rect 9904 1538 10064 1554
rect 17584 19222 17744 19238
rect 17584 19194 17598 19222
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17730 19194 17744 19222
rect 17584 18438 17744 19194
rect 17584 18410 17598 18438
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17730 18410 17744 18438
rect 17584 17654 17744 18410
rect 17584 17626 17598 17654
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17730 17626 17744 17654
rect 17584 16870 17744 17626
rect 17584 16842 17598 16870
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17730 16842 17744 16870
rect 17584 16086 17744 16842
rect 17584 16058 17598 16086
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17730 16058 17744 16086
rect 17584 15302 17744 16058
rect 17584 15274 17598 15302
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17730 15274 17744 15302
rect 17584 14518 17744 15274
rect 17584 14490 17598 14518
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17730 14490 17744 14518
rect 17584 13734 17744 14490
rect 17584 13706 17598 13734
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17730 13706 17744 13734
rect 17584 12950 17744 13706
rect 17584 12922 17598 12950
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17730 12922 17744 12950
rect 17584 12166 17744 12922
rect 17584 12138 17598 12166
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17730 12138 17744 12166
rect 17584 11382 17744 12138
rect 17584 11354 17598 11382
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17730 11354 17744 11382
rect 17584 10598 17744 11354
rect 17584 10570 17598 10598
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17730 10570 17744 10598
rect 17584 9814 17744 10570
rect 17584 9786 17598 9814
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17730 9786 17744 9814
rect 17584 9030 17744 9786
rect 17584 9002 17598 9030
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17730 9002 17744 9030
rect 17584 8246 17744 9002
rect 17584 8218 17598 8246
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17730 8218 17744 8246
rect 17584 7462 17744 8218
rect 17584 7434 17598 7462
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17730 7434 17744 7462
rect 17584 6678 17744 7434
rect 17584 6650 17598 6678
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17730 6650 17744 6678
rect 17584 5894 17744 6650
rect 17584 5866 17598 5894
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17730 5866 17744 5894
rect 17584 5110 17744 5866
rect 17584 5082 17598 5110
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17730 5082 17744 5110
rect 17584 4326 17744 5082
rect 17584 4298 17598 4326
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17730 4298 17744 4326
rect 17584 3542 17744 4298
rect 17584 3514 17598 3542
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17730 3514 17744 3542
rect 17584 2758 17744 3514
rect 17584 2730 17598 2758
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17730 2730 17744 2758
rect 17584 1974 17744 2730
rect 17584 1946 17598 1974
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17730 1946 17744 1974
rect 17584 1538 17744 1946
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _118_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 12096 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _119_
timestamp 1698175906
transform -1 0 12376 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _120_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 13664 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _121_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 13272 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _122_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 12096 0 -1 11760
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _123_
timestamp 1698175906
transform -1 0 10416 0 -1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _124_
timestamp 1698175906
transform -1 0 9576 0 -1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _125_
timestamp 1698175906
transform -1 0 13440 0 1 12544
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _126_
timestamp 1698175906
transform 1 0 7168 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _127_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10584 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _128_
timestamp 1698175906
transform 1 0 7504 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _129_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8176 0 -1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _130_
timestamp 1698175906
transform -1 0 11592 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _131_
timestamp 1698175906
transform -1 0 11480 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _132_
timestamp 1698175906
transform 1 0 10584 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _133_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10416 0 -1 10976
box -43 -43 2059 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _134_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 12432 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _135_
timestamp 1698175906
transform -1 0 13160 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _136_
timestamp 1698175906
transform 1 0 7952 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _137_
timestamp 1698175906
transform 1 0 8288 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _138_
timestamp 1698175906
transform 1 0 9800 0 1 8624
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _139_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 12712 0 -1 10192
box -43 -43 883 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _140_
timestamp 1698175906
transform -1 0 14784 0 1 7840
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _141_
timestamp 1698175906
transform -1 0 10136 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _142_
timestamp 1698175906
transform 1 0 7616 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _143_
timestamp 1698175906
transform 1 0 11368 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _144_
timestamp 1698175906
transform -1 0 10472 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _145_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10360 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _146_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10584 0 -1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _147_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10808 0 1 9408
box -43 -43 715 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _148_
timestamp 1698175906
transform 1 0 13160 0 -1 10976
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _149_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 13104 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _150_
timestamp 1698175906
transform 1 0 13832 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _151_
timestamp 1698175906
transform 1 0 7840 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _152_
timestamp 1698175906
transform 1 0 10024 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _153_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 11872 0 1 10976
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _154_
timestamp 1698175906
transform 1 0 14056 0 1 10976
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _155_
timestamp 1698175906
transform -1 0 13104 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _156_
timestamp 1698175906
transform -1 0 14056 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _157_
timestamp 1698175906
transform -1 0 11144 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _158_
timestamp 1698175906
transform 1 0 11032 0 1 8624
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _159_
timestamp 1698175906
transform -1 0 10584 0 -1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _160_
timestamp 1698175906
transform -1 0 11144 0 1 7056
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _161_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10472 0 -1 7840
box -43 -43 659 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _162_
timestamp 1698175906
transform -1 0 10976 0 -1 12544
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _163_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 9856 0 -1 10976
box -43 -43 771 435
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _164_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 9632 0 -1 10192
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _165_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10584 0 1 12544
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _166_
timestamp 1698175906
transform -1 0 11256 0 1 12544
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _167_
timestamp 1698175906
transform -1 0 9128 0 -1 10976
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _168_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 8848 0 1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _169_
timestamp 1698175906
transform 1 0 9016 0 1 13328
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _170_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8960 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _171_
timestamp 1698175906
transform -1 0 7336 0 1 9408
box -43 -43 715 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _172_
timestamp 1698175906
transform 1 0 6776 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _173_
timestamp 1698175906
transform 1 0 9968 0 -1 11760
box -43 -43 715 435
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _174_
timestamp 1698175906
transform 1 0 11760 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _175_
timestamp 1698175906
transform 1 0 12208 0 1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _176_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 12040 0 1 9408
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _177_
timestamp 1698175906
transform -1 0 11760 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _178_
timestamp 1698175906
transform -1 0 8848 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _179_
timestamp 1698175906
transform -1 0 9744 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _180_
timestamp 1698175906
transform -1 0 9408 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _181_
timestamp 1698175906
transform 1 0 8624 0 -1 9408
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _182_
timestamp 1698175906
transform 1 0 7616 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _183_
timestamp 1698175906
transform -1 0 7728 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _184_
timestamp 1698175906
transform -1 0 9408 0 -1 8624
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _185_
timestamp 1698175906
transform 1 0 9464 0 1 7056
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _186_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9408 0 -1 7840
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _187_
timestamp 1698175906
transform -1 0 9184 0 -1 7056
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _188_
timestamp 1698175906
transform 1 0 8512 0 1 7056
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _189_
timestamp 1698175906
transform 1 0 8792 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _190_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9576 0 -1 9408
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _191_
timestamp 1698175906
transform 1 0 11648 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _192_
timestamp 1698175906
transform 1 0 11704 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _193_
timestamp 1698175906
transform -1 0 12768 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _194_
timestamp 1698175906
transform -1 0 11368 0 1 11760
box -43 -43 771 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _195_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10640 0 -1 11760
box -43 -43 771 435
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _196_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 11032 0 1 13328
box -43 -43 659 435
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _197_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 11144 0 -1 13328
box -43 -43 1331 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _198_
timestamp 1698175906
transform -1 0 11032 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _199_
timestamp 1698175906
transform -1 0 10472 0 1 12544
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _200_
timestamp 1698175906
transform 1 0 10584 0 1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _201_
timestamp 1698175906
transform -1 0 10472 0 1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _202_
timestamp 1698175906
transform -1 0 11312 0 1 10192
box -43 -43 771 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _203_
timestamp 1698175906
transform 1 0 13776 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _204_
timestamp 1698175906
transform -1 0 13552 0 -1 11760
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _205_
timestamp 1698175906
transform -1 0 15008 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _206_
timestamp 1698175906
transform 1 0 13664 0 1 7840
box -43 -43 659 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _207_
timestamp 1698175906
transform 1 0 14952 0 1 9408
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _208_
timestamp 1698175906
transform -1 0 14952 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _209_
timestamp 1698175906
transform 1 0 13552 0 1 9408
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _210_
timestamp 1698175906
transform 1 0 13888 0 1 9408
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _211_
timestamp 1698175906
transform -1 0 13944 0 -1 10192
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _212_
timestamp 1698175906
transform -1 0 11536 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _213_
timestamp 1698175906
transform 1 0 11256 0 1 7056
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _214_
timestamp 1698175906
transform -1 0 8512 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _215_
timestamp 1698175906
transform -1 0 7616 0 -1 7840
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _216_
timestamp 1698175906
transform -1 0 7616 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _217_
timestamp 1698175906
transform -1 0 7224 0 1 7056
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _218_
timestamp 1698175906
transform -1 0 7112 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _219_
timestamp 1698175906
transform -1 0 7896 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _220_
timestamp 1698175906
transform -1 0 9688 0 1 10976
box -43 -43 883 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _221_
timestamp 1698175906
transform -1 0 9016 0 1 9408
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _222_
timestamp 1698175906
transform 1 0 7448 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _223_
timestamp 1698175906
transform -1 0 7672 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _224_
timestamp 1698175906
transform -1 0 6496 0 1 12544
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _225_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8624 0 -1 13328
box -43 -43 715 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _226_
timestamp 1698175906
transform -1 0 8512 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _227_
timestamp 1698175906
transform 1 0 7616 0 -1 13328
box -43 -43 715 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _228_
timestamp 1698175906
transform -1 0 7280 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _229_
timestamp 1698175906
transform -1 0 9968 0 -1 11760
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _230_
timestamp 1698175906
transform -1 0 7224 0 1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _231_
timestamp 1698175906
transform 1 0 6776 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _232_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 9408 0 1 8624
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _233_
timestamp 1698175906
transform -1 0 9688 0 -1 8624
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _234_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9072 0 1 7840
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _235_
timestamp 1698175906
transform -1 0 8512 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _236_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 12544 0 -1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _237_
timestamp 1698175906
transform 1 0 13384 0 -1 7840
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _238_
timestamp 1698175906
transform 1 0 13552 0 -1 11760
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _239_
timestamp 1698175906
transform 1 0 9184 0 -1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _240_
timestamp 1698175906
transform 1 0 8176 0 1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _241_
timestamp 1698175906
transform 1 0 5432 0 -1 9408
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _242_
timestamp 1698175906
transform 1 0 5544 0 -1 10192
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _243_
timestamp 1698175906
transform 1 0 11984 0 1 10976
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _244_
timestamp 1698175906
transform -1 0 12992 0 1 8624
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _245_
timestamp 1698175906
transform -1 0 7616 0 -1 11760
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _246_
timestamp 1698175906
transform 1 0 8456 0 1 6272
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _247_
timestamp 1698175906
transform 1 0 6888 0 -1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _248_
timestamp 1698175906
transform 1 0 11592 0 1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _249_
timestamp 1698175906
transform 1 0 11648 0 1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _250_
timestamp 1698175906
transform 1 0 10136 0 -1 14112
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _251_
timestamp 1698175906
transform 1 0 9520 0 -1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _252_
timestamp 1698175906
transform 1 0 13776 0 -1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _253_
timestamp 1698175906
transform 1 0 13608 0 -1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _254_
timestamp 1698175906
transform 1 0 13944 0 -1 10192
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _255_
timestamp 1698175906
transform 1 0 13776 0 -1 9408
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _256_
timestamp 1698175906
transform 1 0 10808 0 -1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _257_
timestamp 1698175906
transform -1 0 7224 0 -1 7840
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _258_
timestamp 1698175906
transform -1 0 7168 0 -1 8624
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _259_
timestamp 1698175906
transform 1 0 5488 0 -1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _260_
timestamp 1698175906
transform 1 0 7392 0 1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _261_
timestamp 1698175906
transform 1 0 6104 0 -1 14112
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _262_
timestamp 1698175906
transform -1 0 7112 0 -1 10976
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _263_
timestamp 1698175906
transform 1 0 7448 0 1 7840
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _264_
timestamp 1698175906
transform 1 0 12880 0 -1 14112
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _265_
timestamp 1698175906
transform 1 0 15176 0 -1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__236__CLK dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 14280 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__237__CLK
timestamp 1698175906
transform 1 0 15120 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__238__CLK
timestamp 1698175906
transform 1 0 13440 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__239__CLK
timestamp 1698175906
transform 1 0 8736 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__240__CLK
timestamp 1698175906
transform 1 0 9912 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__241__CLK
timestamp 1698175906
transform 1 0 7168 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__242__CLK
timestamp 1698175906
transform 1 0 7336 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__243__CLK
timestamp 1698175906
transform 1 0 13776 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__244__CLK
timestamp 1698175906
transform 1 0 13104 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__245__CLK
timestamp 1698175906
transform 1 0 7616 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__246__CLK
timestamp 1698175906
transform 1 0 10192 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__247__CLK
timestamp 1698175906
transform 1 0 8904 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__248__CLK
timestamp 1698175906
transform 1 0 13328 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__249__CLK
timestamp 1698175906
transform 1 0 13384 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__250__CLK
timestamp 1698175906
transform -1 0 11984 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__251__CLK
timestamp 1698175906
transform 1 0 9408 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__252__CLK
timestamp 1698175906
transform 1 0 13664 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__253__CLK
timestamp 1698175906
transform 1 0 13496 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__254__CLK
timestamp 1698175906
transform 1 0 14000 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__255__CLK
timestamp 1698175906
transform 1 0 13664 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__256__CLK
timestamp 1698175906
transform 1 0 12656 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__257__CLK
timestamp 1698175906
transform 1 0 7728 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__258__CLK
timestamp 1698175906
transform 1 0 7168 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__259__CLK
timestamp 1698175906
transform 1 0 7224 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__260__CLK
timestamp 1698175906
transform 1 0 9520 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__261__CLK
timestamp 1698175906
transform -1 0 7952 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__262__CLK
timestamp 1698175906
transform 1 0 7224 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__263__CLK
timestamp 1698175906
transform 1 0 9744 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1698175906
transform 1 0 8736 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9632 0 -1 10192
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1698175906
transform -1 0 10472 0 1 10192
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1698175906
transform 1 0 11592 0 1 10192
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 784 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698175906
transform 1 0 2688 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698175906
transform 1 0 4592 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698175906
transform 1 0 6496 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_138 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8400 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_142 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8624 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_172
timestamp 1698175906
transform 1 0 10304 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_176
timestamp 1698175906
transform 1 0 10528 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_232
timestamp 1698175906
transform 1 0 13664 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_236
timestamp 1698175906
transform 1 0 13888 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_240
timestamp 1698175906
transform 1 0 14112 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_274
timestamp 1698175906
transform 1 0 16016 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_308
timestamp 1698175906
transform 1 0 17920 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_342
timestamp 1698175906
transform 1 0 19824 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_346
timestamp 1698175906
transform 1 0 20048 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_348 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 20160 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 784 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698175906
transform 1 0 4368 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698175906
transform 1 0 4704 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698175906
transform 1 0 8288 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_142 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8624 0 -1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_158
timestamp 1698175906
transform 1 0 9520 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_162
timestamp 1698175906
transform 1 0 9744 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_189
timestamp 1698175906
transform 1 0 11256 0 -1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_205
timestamp 1698175906
transform 1 0 12152 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_209
timestamp 1698175906
transform 1 0 12376 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_238
timestamp 1698175906
transform 1 0 14000 0 -1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_270 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 15792 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_278
timestamp 1698175906
transform 1 0 16240 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_282
timestamp 1698175906
transform 1 0 16464 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_346
timestamp 1698175906
transform 1 0 20048 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_348
timestamp 1698175906
transform 1 0 20160 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698175906
transform 1 0 784 0 1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698175906
transform 1 0 2576 0 1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698175906
transform 1 0 2744 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698175906
transform 1 0 6328 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_107
timestamp 1698175906
transform 1 0 6664 0 1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_139
timestamp 1698175906
transform 1 0 8456 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_143
timestamp 1698175906
transform 1 0 8680 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_171
timestamp 1698175906
transform 1 0 10248 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_177
timestamp 1698175906
transform 1 0 10584 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_241
timestamp 1698175906
transform 1 0 14168 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698175906
transform 1 0 14504 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698175906
transform 1 0 18088 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_317
timestamp 1698175906
transform 1 0 18424 0 1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698175906
transform 1 0 784 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698175906
transform 1 0 4368 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698175906
transform 1 0 4704 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698175906
transform 1 0 8288 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_142
timestamp 1698175906
transform 1 0 8624 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_206
timestamp 1698175906
transform 1 0 12208 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_212
timestamp 1698175906
transform 1 0 12544 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_276
timestamp 1698175906
transform 1 0 16128 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_282
timestamp 1698175906
transform 1 0 16464 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_346
timestamp 1698175906
transform 1 0 20048 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_348
timestamp 1698175906
transform 1 0 20160 0 -1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698175906
transform 1 0 784 0 1 3136
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698175906
transform 1 0 2576 0 1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698175906
transform 1 0 2744 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698175906
transform 1 0 6328 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_107
timestamp 1698175906
transform 1 0 6664 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698175906
transform 1 0 10248 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_177
timestamp 1698175906
transform 1 0 10584 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_241
timestamp 1698175906
transform 1 0 14168 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698175906
transform 1 0 14504 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698175906
transform 1 0 18088 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_317
timestamp 1698175906
transform 1 0 18424 0 1 3136
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698175906
transform 1 0 784 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698175906
transform 1 0 4368 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698175906
transform 1 0 4704 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698175906
transform 1 0 8288 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_142
timestamp 1698175906
transform 1 0 8624 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_206
timestamp 1698175906
transform 1 0 12208 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_212
timestamp 1698175906
transform 1 0 12544 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698175906
transform 1 0 16128 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_282
timestamp 1698175906
transform 1 0 16464 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_346
timestamp 1698175906
transform 1 0 20048 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_348
timestamp 1698175906
transform 1 0 20160 0 -1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698175906
transform 1 0 784 0 1 3920
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698175906
transform 1 0 2576 0 1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698175906
transform 1 0 2744 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698175906
transform 1 0 6328 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_107
timestamp 1698175906
transform 1 0 6664 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_171
timestamp 1698175906
transform 1 0 10248 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_177
timestamp 1698175906
transform 1 0 10584 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_241
timestamp 1698175906
transform 1 0 14168 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_247
timestamp 1698175906
transform 1 0 14504 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_311
timestamp 1698175906
transform 1 0 18088 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_317
timestamp 1698175906
transform 1 0 18424 0 1 3920
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698175906
transform 1 0 784 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698175906
transform 1 0 4368 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_72
timestamp 1698175906
transform 1 0 4704 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698175906
transform 1 0 8288 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_142
timestamp 1698175906
transform 1 0 8624 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_206
timestamp 1698175906
transform 1 0 12208 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_212
timestamp 1698175906
transform 1 0 12544 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_276
timestamp 1698175906
transform 1 0 16128 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_282
timestamp 1698175906
transform 1 0 16464 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_346
timestamp 1698175906
transform 1 0 20048 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_348
timestamp 1698175906
transform 1 0 20160 0 -1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698175906
transform 1 0 784 0 1 4704
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698175906
transform 1 0 2576 0 1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_37
timestamp 1698175906
transform 1 0 2744 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_101
timestamp 1698175906
transform 1 0 6328 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_107
timestamp 1698175906
transform 1 0 6664 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_171
timestamp 1698175906
transform 1 0 10248 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_177
timestamp 1698175906
transform 1 0 10584 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_241
timestamp 1698175906
transform 1 0 14168 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_247
timestamp 1698175906
transform 1 0 14504 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_311
timestamp 1698175906
transform 1 0 18088 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_317
timestamp 1698175906
transform 1 0 18424 0 1 4704
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698175906
transform 1 0 784 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698175906
transform 1 0 4368 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_72
timestamp 1698175906
transform 1 0 4704 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_136
timestamp 1698175906
transform 1 0 8288 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_142
timestamp 1698175906
transform 1 0 8624 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_206
timestamp 1698175906
transform 1 0 12208 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_212
timestamp 1698175906
transform 1 0 12544 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_276
timestamp 1698175906
transform 1 0 16128 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_282
timestamp 1698175906
transform 1 0 16464 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_346
timestamp 1698175906
transform 1 0 20048 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_348
timestamp 1698175906
transform 1 0 20160 0 -1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698175906
transform 1 0 784 0 1 5488
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698175906
transform 1 0 2576 0 1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_37
timestamp 1698175906
transform 1 0 2744 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698175906
transform 1 0 6328 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_107
timestamp 1698175906
transform 1 0 6664 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_171
timestamp 1698175906
transform 1 0 10248 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_177
timestamp 1698175906
transform 1 0 10584 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_241
timestamp 1698175906
transform 1 0 14168 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_247
timestamp 1698175906
transform 1 0 14504 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_311
timestamp 1698175906
transform 1 0 18088 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_317
timestamp 1698175906
transform 1 0 18424 0 1 5488
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2
timestamp 1698175906
transform 1 0 784 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698175906
transform 1 0 4368 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_72
timestamp 1698175906
transform 1 0 4704 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698175906
transform 1 0 8288 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_142
timestamp 1698175906
transform 1 0 8624 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_206
timestamp 1698175906
transform 1 0 12208 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_212
timestamp 1698175906
transform 1 0 12544 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_276
timestamp 1698175906
transform 1 0 16128 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_282
timestamp 1698175906
transform 1 0 16464 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_346
timestamp 1698175906
transform 1 0 20048 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_348
timestamp 1698175906
transform 1 0 20160 0 -1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698175906
transform 1 0 784 0 1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698175906
transform 1 0 2576 0 1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_37
timestamp 1698175906
transform 1 0 2744 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698175906
transform 1 0 6328 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_107
timestamp 1698175906
transform 1 0 6664 0 1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_168
timestamp 1698175906
transform 1 0 10080 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_172
timestamp 1698175906
transform 1 0 10304 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_174
timestamp 1698175906
transform 1 0 10416 0 1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_177
timestamp 1698175906
transform 1 0 10584 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_241
timestamp 1698175906
transform 1 0 14168 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_247
timestamp 1698175906
transform 1 0 14504 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_311
timestamp 1698175906
transform 1 0 18088 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_317
timestamp 1698175906
transform 1 0 18424 0 1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_2
timestamp 1698175906
transform 1 0 784 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_66
timestamp 1698175906
transform 1 0 4368 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_72
timestamp 1698175906
transform 1 0 4704 0 -1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_104
timestamp 1698175906
transform 1 0 6496 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_108
timestamp 1698175906
transform 1 0 6720 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_110
timestamp 1698175906
transform 1 0 6832 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_142
timestamp 1698175906
transform 1 0 8624 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_212
timestamp 1698175906
transform 1 0 12544 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_216
timestamp 1698175906
transform 1 0 12768 0 -1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_224
timestamp 1698175906
transform 1 0 13216 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_228
timestamp 1698175906
transform 1 0 13440 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_260
timestamp 1698175906
transform 1 0 15232 0 -1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_276
timestamp 1698175906
transform 1 0 16128 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_282
timestamp 1698175906
transform 1 0 16464 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_346
timestamp 1698175906
transform 1 0 20048 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_348
timestamp 1698175906
transform 1 0 20160 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698175906
transform 1 0 784 0 1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698175906
transform 1 0 2576 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_37
timestamp 1698175906
transform 1 0 2744 0 1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_101
timestamp 1698175906
transform 1 0 6328 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_107
timestamp 1698175906
transform 1 0 6664 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_109
timestamp 1698175906
transform 1 0 6776 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_117
timestamp 1698175906
transform 1 0 7224 0 1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_133
timestamp 1698175906
transform 1 0 8120 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_137
timestamp 1698175906
transform 1 0 8344 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_139
timestamp 1698175906
transform 1 0 8456 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_145
timestamp 1698175906
transform 1 0 8792 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_149
timestamp 1698175906
transform 1 0 9016 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_163
timestamp 1698175906
transform 1 0 9800 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_171
timestamp 1698175906
transform 1 0 10248 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_177
timestamp 1698175906
transform 1 0 10584 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_179
timestamp 1698175906
transform 1 0 10696 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_187
timestamp 1698175906
transform 1 0 11144 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_224
timestamp 1698175906
transform 1 0 13216 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_228
timestamp 1698175906
transform 1 0 13440 0 1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_244
timestamp 1698175906
transform 1 0 14336 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_247
timestamp 1698175906
transform 1 0 14504 0 1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_311
timestamp 1698175906
transform 1 0 18088 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_317
timestamp 1698175906
transform 1 0 18424 0 1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_2
timestamp 1698175906
transform 1 0 784 0 -1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_66
timestamp 1698175906
transform 1 0 4368 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_72
timestamp 1698175906
transform 1 0 4704 0 -1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_124
timestamp 1698175906
transform 1 0 7616 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_128
timestamp 1698175906
transform 1 0 7840 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_136
timestamp 1698175906
transform 1 0 8288 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_142
timestamp 1698175906
transform 1 0 8624 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_144
timestamp 1698175906
transform 1 0 8736 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_153
timestamp 1698175906
transform 1 0 9240 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_155
timestamp 1698175906
transform 1 0 9352 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_165
timestamp 1698175906
transform 1 0 9912 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_173
timestamp 1698175906
transform 1 0 10360 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_194
timestamp 1698175906
transform 1 0 11536 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_204
timestamp 1698175906
transform 1 0 12096 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_208
timestamp 1698175906
transform 1 0 12320 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_212
timestamp 1698175906
transform 1 0 12544 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_220
timestamp 1698175906
transform 1 0 12992 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_224
timestamp 1698175906
transform 1 0 13216 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_226
timestamp 1698175906
transform 1 0 13328 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_256
timestamp 1698175906
transform 1 0 15008 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_260
timestamp 1698175906
transform 1 0 15232 0 -1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_276
timestamp 1698175906
transform 1 0 16128 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_282
timestamp 1698175906
transform 1 0 16464 0 -1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_346
timestamp 1698175906
transform 1 0 20048 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_348
timestamp 1698175906
transform 1 0 20160 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_28
timestamp 1698175906
transform 1 0 2240 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_32
timestamp 1698175906
transform 1 0 2464 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698175906
transform 1 0 2576 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_37
timestamp 1698175906
transform 1 0 2744 0 1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_101
timestamp 1698175906
transform 1 0 6328 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_115
timestamp 1698175906
transform 1 0 7112 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_119
timestamp 1698175906
transform 1 0 7336 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_160
timestamp 1698175906
transform 1 0 9632 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_164
timestamp 1698175906
transform 1 0 9856 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_172
timestamp 1698175906
transform 1 0 10304 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_174
timestamp 1698175906
transform 1 0 10416 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_177
timestamp 1698175906
transform 1 0 10584 0 1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_193
timestamp 1698175906
transform 1 0 11480 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_205
timestamp 1698175906
transform 1 0 12152 0 1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_221
timestamp 1698175906
transform 1 0 13048 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_229
timestamp 1698175906
transform 1 0 13496 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_231
timestamp 1698175906
transform 1 0 13608 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_243
timestamp 1698175906
transform 1 0 14280 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_256
timestamp 1698175906
transform 1 0 15008 0 1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_288
timestamp 1698175906
transform 1 0 16800 0 1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_304
timestamp 1698175906
transform 1 0 17696 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_312
timestamp 1698175906
transform 1 0 18144 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_314
timestamp 1698175906
transform 1 0 18256 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_317
timestamp 1698175906
transform 1 0 18424 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_321
timestamp 1698175906
transform 1 0 18648 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_28
timestamp 1698175906
transform 1 0 2240 0 -1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_60
timestamp 1698175906
transform 1 0 4032 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_68
timestamp 1698175906
transform 1 0 4480 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_72
timestamp 1698175906
transform 1 0 4704 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_80
timestamp 1698175906
transform 1 0 5152 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_84
timestamp 1698175906
transform 1 0 5376 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_86
timestamp 1698175906
transform 1 0 5488 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_124
timestamp 1698175906
transform 1 0 7616 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_161
timestamp 1698175906
transform 1 0 9688 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_169
timestamp 1698175906
transform 1 0 10136 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_193
timestamp 1698175906
transform 1 0 11480 0 -1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_209
timestamp 1698175906
transform 1 0 12376 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_212
timestamp 1698175906
transform 1 0 12544 0 -1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_228
timestamp 1698175906
transform 1 0 13440 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_232
timestamp 1698175906
transform 1 0 13664 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_234
timestamp 1698175906
transform 1 0 13776 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_243
timestamp 1698175906
transform 1 0 14280 0 -1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_275
timestamp 1698175906
transform 1 0 16072 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_279
timestamp 1698175906
transform 1 0 16296 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_282
timestamp 1698175906
transform 1 0 16464 0 -1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_314
timestamp 1698175906
transform 1 0 18256 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_322
timestamp 1698175906
transform 1 0 18704 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_2
timestamp 1698175906
transform 1 0 784 0 1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698175906
transform 1 0 2576 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_37
timestamp 1698175906
transform 1 0 2744 0 1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_101
timestamp 1698175906
transform 1 0 6328 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_107
timestamp 1698175906
transform 1 0 6664 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_115
timestamp 1698175906
transform 1 0 7112 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_118
timestamp 1698175906
transform 1 0 7280 0 1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_134
timestamp 1698175906
transform 1 0 8176 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_142
timestamp 1698175906
transform 1 0 8624 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_156
timestamp 1698175906
transform 1 0 9408 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_160
timestamp 1698175906
transform 1 0 9632 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_162
timestamp 1698175906
transform 1 0 9744 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_168
timestamp 1698175906
transform 1 0 10080 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_172
timestamp 1698175906
transform 1 0 10304 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_174
timestamp 1698175906
transform 1 0 10416 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_177
timestamp 1698175906
transform 1 0 10584 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_190
timestamp 1698175906
transform 1 0 11312 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_220
timestamp 1698175906
transform 1 0 12992 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_224
timestamp 1698175906
transform 1 0 13216 0 1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_240
timestamp 1698175906
transform 1 0 14112 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_244
timestamp 1698175906
transform 1 0 14336 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_247
timestamp 1698175906
transform 1 0 14504 0 1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_311
timestamp 1698175906
transform 1 0 18088 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_317
timestamp 1698175906
transform 1 0 18424 0 1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_2
timestamp 1698175906
transform 1 0 784 0 -1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_66
timestamp 1698175906
transform 1 0 4368 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_72
timestamp 1698175906
transform 1 0 4704 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_80
timestamp 1698175906
transform 1 0 5152 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_84
timestamp 1698175906
transform 1 0 5376 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_114
timestamp 1698175906
transform 1 0 7056 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_118
timestamp 1698175906
transform 1 0 7280 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_126
timestamp 1698175906
transform 1 0 7728 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_136
timestamp 1698175906
transform 1 0 8288 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_156
timestamp 1698175906
transform 1 0 9408 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_158
timestamp 1698175906
transform 1 0 9520 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_169
timestamp 1698175906
transform 1 0 10136 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_187
timestamp 1698175906
transform 1 0 11144 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_189
timestamp 1698175906
transform 1 0 11256 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_204
timestamp 1698175906
transform 1 0 12096 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_208
timestamp 1698175906
transform 1 0 12320 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_212
timestamp 1698175906
transform 1 0 12544 0 -1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_228
timestamp 1698175906
transform 1 0 13440 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_263
timestamp 1698175906
transform 1 0 15400 0 -1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_279
timestamp 1698175906
transform 1 0 16296 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_282
timestamp 1698175906
transform 1 0 16464 0 -1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_346
timestamp 1698175906
transform 1 0 20048 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_348
timestamp 1698175906
transform 1 0 20160 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_2
timestamp 1698175906
transform 1 0 784 0 1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698175906
transform 1 0 2576 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_37
timestamp 1698175906
transform 1 0 2744 0 1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_101
timestamp 1698175906
transform 1 0 6328 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_119
timestamp 1698175906
transform 1 0 7336 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_123
timestamp 1698175906
transform 1 0 7560 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_132
timestamp 1698175906
transform 1 0 8064 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_149
timestamp 1698175906
transform 1 0 9016 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_162
timestamp 1698175906
transform 1 0 9744 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_209
timestamp 1698175906
transform 1 0 12376 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_213
timestamp 1698175906
transform 1 0 12600 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_215
timestamp 1698175906
transform 1 0 12712 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_235
timestamp 1698175906
transform 1 0 13832 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_260
timestamp 1698175906
transform 1 0 15232 0 1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_292
timestamp 1698175906
transform 1 0 17024 0 1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_308
timestamp 1698175906
transform 1 0 17920 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_312
timestamp 1698175906
transform 1 0 18144 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_314
timestamp 1698175906
transform 1 0 18256 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_317
timestamp 1698175906
transform 1 0 18424 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_321
timestamp 1698175906
transform 1 0 18648 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_2
timestamp 1698175906
transform 1 0 784 0 -1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_66
timestamp 1698175906
transform 1 0 4368 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_72
timestamp 1698175906
transform 1 0 4704 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_80
timestamp 1698175906
transform 1 0 5152 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_84
timestamp 1698175906
transform 1 0 5376 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_86
timestamp 1698175906
transform 1 0 5488 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_136
timestamp 1698175906
transform 1 0 8288 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_142
timestamp 1698175906
transform 1 0 8624 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_212
timestamp 1698175906
transform 1 0 12544 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_214
timestamp 1698175906
transform 1 0 12656 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_230
timestamp 1698175906
transform 1 0 13552 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_266
timestamp 1698175906
transform 1 0 15568 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_274
timestamp 1698175906
transform 1 0 16016 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_278
timestamp 1698175906
transform 1 0 16240 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_282
timestamp 1698175906
transform 1 0 16464 0 -1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_314
timestamp 1698175906
transform 1 0 18256 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_322
timestamp 1698175906
transform 1 0 18704 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_2
timestamp 1698175906
transform 1 0 784 0 1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698175906
transform 1 0 2576 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_37
timestamp 1698175906
transform 1 0 2744 0 1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_101
timestamp 1698175906
transform 1 0 6328 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_107
timestamp 1698175906
transform 1 0 6664 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_117
timestamp 1698175906
transform 1 0 7224 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_121
timestamp 1698175906
transform 1 0 7448 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_190
timestamp 1698175906
transform 1 0 11312 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_247
timestamp 1698175906
transform 1 0 14504 0 1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_311
timestamp 1698175906
transform 1 0 18088 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_317
timestamp 1698175906
transform 1 0 18424 0 1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_2
timestamp 1698175906
transform 1 0 784 0 -1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_66
timestamp 1698175906
transform 1 0 4368 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_72
timestamp 1698175906
transform 1 0 4704 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_80
timestamp 1698175906
transform 1 0 5152 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_84
timestamp 1698175906
transform 1 0 5376 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_115
timestamp 1698175906
transform 1 0 7112 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_119
timestamp 1698175906
transform 1 0 7336 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_127
timestamp 1698175906
transform 1 0 7784 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_131
timestamp 1698175906
transform 1 0 8008 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_133
timestamp 1698175906
transform 1 0 8120 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_142
timestamp 1698175906
transform 1 0 8624 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_164
timestamp 1698175906
transform 1 0 9856 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_212
timestamp 1698175906
transform 1 0 12544 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_214
timestamp 1698175906
transform 1 0 12656 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_232
timestamp 1698175906
transform 1 0 13664 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_236
timestamp 1698175906
transform 1 0 13888 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_240
timestamp 1698175906
transform 1 0 14112 0 -1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_272
timestamp 1698175906
transform 1 0 15904 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_282
timestamp 1698175906
transform 1 0 16464 0 -1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_346
timestamp 1698175906
transform 1 0 20048 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_348
timestamp 1698175906
transform 1 0 20160 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_2
timestamp 1698175906
transform 1 0 784 0 1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698175906
transform 1 0 2576 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_37
timestamp 1698175906
transform 1 0 2744 0 1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_101
timestamp 1698175906
transform 1 0 6328 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_107
timestamp 1698175906
transform 1 0 6664 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_117
timestamp 1698175906
transform 1 0 7224 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_119
timestamp 1698175906
transform 1 0 7336 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_126
timestamp 1698175906
transform 1 0 7728 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_161
timestamp 1698175906
transform 1 0 9688 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_165
timestamp 1698175906
transform 1 0 9912 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_200
timestamp 1698175906
transform 1 0 11872 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_244
timestamp 1698175906
transform 1 0 14336 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_247
timestamp 1698175906
transform 1 0 14504 0 1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_311
timestamp 1698175906
transform 1 0 18088 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_317
timestamp 1698175906
transform 1 0 18424 0 1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_28
timestamp 1698175906
transform 1 0 2240 0 -1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_60
timestamp 1698175906
transform 1 0 4032 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_68
timestamp 1698175906
transform 1 0 4480 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_72
timestamp 1698175906
transform 1 0 4704 0 -1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_88
timestamp 1698175906
transform 1 0 5600 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_92
timestamp 1698175906
transform 1 0 5824 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_94
timestamp 1698175906
transform 1 0 5936 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_132
timestamp 1698175906
transform 1 0 8064 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_142
timestamp 1698175906
transform 1 0 8624 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_150
timestamp 1698175906
transform 1 0 9072 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_152
timestamp 1698175906
transform 1 0 9184 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_204
timestamp 1698175906
transform 1 0 12096 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_208
timestamp 1698175906
transform 1 0 12320 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_212
timestamp 1698175906
transform 1 0 12544 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_216
timestamp 1698175906
transform 1 0 12768 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_265
timestamp 1698175906
transform 1 0 15512 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_273
timestamp 1698175906
transform 1 0 15960 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_277
timestamp 1698175906
transform 1 0 16184 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_279
timestamp 1698175906
transform 1 0 16296 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_282
timestamp 1698175906
transform 1 0 16464 0 -1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_314
timestamp 1698175906
transform 1 0 18256 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_322
timestamp 1698175906
transform 1 0 18704 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_28
timestamp 1698175906
transform 1 0 2240 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_32
timestamp 1698175906
transform 1 0 2464 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698175906
transform 1 0 2576 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_37
timestamp 1698175906
transform 1 0 2744 0 1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_101
timestamp 1698175906
transform 1 0 6328 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_107
timestamp 1698175906
transform 1 0 6664 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_117
timestamp 1698175906
transform 1 0 7224 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_121
timestamp 1698175906
transform 1 0 7448 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_123
timestamp 1698175906
transform 1 0 7560 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_126
timestamp 1698175906
transform 1 0 7728 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_134
timestamp 1698175906
transform 1 0 8176 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_138
timestamp 1698175906
transform 1 0 8400 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_146
timestamp 1698175906
transform 1 0 8848 0 1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_162
timestamp 1698175906
transform 1 0 9744 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_170
timestamp 1698175906
transform 1 0 10192 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_174
timestamp 1698175906
transform 1 0 10416 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_177
timestamp 1698175906
transform 1 0 10584 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_191
timestamp 1698175906
transform 1 0 11368 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_195
timestamp 1698175906
transform 1 0 11592 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_197
timestamp 1698175906
transform 1 0 11704 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_212
timestamp 1698175906
transform 1 0 12544 0 1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_230
timestamp 1698175906
transform 1 0 13552 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_242
timestamp 1698175906
transform 1 0 14224 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_244
timestamp 1698175906
transform 1 0 14336 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_247
timestamp 1698175906
transform 1 0 14504 0 1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_311
timestamp 1698175906
transform 1 0 18088 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_317
timestamp 1698175906
transform 1 0 18424 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_321
timestamp 1698175906
transform 1 0 18648 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_2
timestamp 1698175906
transform 1 0 784 0 -1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_66
timestamp 1698175906
transform 1 0 4368 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_72
timestamp 1698175906
transform 1 0 4704 0 -1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_104
timestamp 1698175906
transform 1 0 6496 0 -1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_120
timestamp 1698175906
transform 1 0 7392 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_129
timestamp 1698175906
transform 1 0 7896 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_137
timestamp 1698175906
transform 1 0 8344 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_139
timestamp 1698175906
transform 1 0 8456 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_142
timestamp 1698175906
transform 1 0 8624 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_146
timestamp 1698175906
transform 1 0 8848 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_156
timestamp 1698175906
transform 1 0 9408 0 -1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_172
timestamp 1698175906
transform 1 0 10304 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_176
timestamp 1698175906
transform 1 0 10528 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_184
timestamp 1698175906
transform 1 0 10976 0 -1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_200
timestamp 1698175906
transform 1 0 11872 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_208
timestamp 1698175906
transform 1 0 12320 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_212
timestamp 1698175906
transform 1 0 12544 0 -1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_228
timestamp 1698175906
transform 1 0 13440 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_263
timestamp 1698175906
transform 1 0 15400 0 -1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_279
timestamp 1698175906
transform 1 0 16296 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_282
timestamp 1698175906
transform 1 0 16464 0 -1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_314
timestamp 1698175906
transform 1 0 18256 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_322
timestamp 1698175906
transform 1 0 18704 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_2
timestamp 1698175906
transform 1 0 784 0 1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698175906
transform 1 0 2576 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_37
timestamp 1698175906
transform 1 0 2744 0 1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_69
timestamp 1698175906
transform 1 0 4536 0 1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_85
timestamp 1698175906
transform 1 0 5432 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_93
timestamp 1698175906
transform 1 0 5880 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_97
timestamp 1698175906
transform 1 0 6104 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_104
timestamp 1698175906
transform 1 0 6496 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_107
timestamp 1698175906
transform 1 0 6664 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_115
timestamp 1698175906
transform 1 0 7112 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_129
timestamp 1698175906
transform 1 0 7896 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_133
timestamp 1698175906
transform 1 0 8120 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_163
timestamp 1698175906
transform 1 0 9800 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_167
timestamp 1698175906
transform 1 0 10024 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_169
timestamp 1698175906
transform 1 0 10136 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_189
timestamp 1698175906
transform 1 0 11256 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_197
timestamp 1698175906
transform 1 0 11704 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_201
timestamp 1698175906
transform 1 0 11928 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_210
timestamp 1698175906
transform 1 0 12432 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_218
timestamp 1698175906
transform 1 0 12880 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_222
timestamp 1698175906
transform 1 0 13104 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_228
timestamp 1698175906
transform 1 0 13440 0 1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_244
timestamp 1698175906
transform 1 0 14336 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_247
timestamp 1698175906
transform 1 0 14504 0 1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_311
timestamp 1698175906
transform 1 0 18088 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_317
timestamp 1698175906
transform 1 0 18424 0 1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_28
timestamp 1698175906
transform 1 0 2240 0 -1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_60
timestamp 1698175906
transform 1 0 4032 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_68
timestamp 1698175906
transform 1 0 4480 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_72
timestamp 1698175906
transform 1 0 4704 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_80
timestamp 1698175906
transform 1 0 5152 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_84
timestamp 1698175906
transform 1 0 5376 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_115
timestamp 1698175906
transform 1 0 7112 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_119
timestamp 1698175906
transform 1 0 7336 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_123
timestamp 1698175906
transform 1 0 7560 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_154
timestamp 1698175906
transform 1 0 9296 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_241
timestamp 1698175906
transform 1 0 14168 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_245
timestamp 1698175906
transform 1 0 14392 0 -1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_277
timestamp 1698175906
transform 1 0 16184 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_279
timestamp 1698175906
transform 1 0 16296 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_282
timestamp 1698175906
transform 1 0 16464 0 -1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_346
timestamp 1698175906
transform 1 0 20048 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_348
timestamp 1698175906
transform 1 0 20160 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_2
timestamp 1698175906
transform 1 0 784 0 1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698175906
transform 1 0 2576 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_37
timestamp 1698175906
transform 1 0 2744 0 1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_101
timestamp 1698175906
transform 1 0 6328 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_107
timestamp 1698175906
transform 1 0 6664 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_111
timestamp 1698175906
transform 1 0 6888 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_113
timestamp 1698175906
transform 1 0 7000 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_118
timestamp 1698175906
transform 1 0 7280 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_156
timestamp 1698175906
transform 1 0 9408 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_160
timestamp 1698175906
transform 1 0 9632 0 1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_168
timestamp 1698175906
transform 1 0 10080 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_225
timestamp 1698175906
transform 1 0 13272 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_229
timestamp 1698175906
transform 1 0 13496 0 1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_247
timestamp 1698175906
transform 1 0 14504 0 1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_311
timestamp 1698175906
transform 1 0 18088 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_317
timestamp 1698175906
transform 1 0 18424 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_321
timestamp 1698175906
transform 1 0 18648 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_2
timestamp 1698175906
transform 1 0 784 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_66
timestamp 1698175906
transform 1 0 4368 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_72
timestamp 1698175906
transform 1 0 4704 0 -1 14112
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_88
timestamp 1698175906
transform 1 0 5600 0 -1 14112
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_96
timestamp 1698175906
transform 1 0 6048 0 -1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_126
timestamp 1698175906
transform 1 0 7728 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_130
timestamp 1698175906
transform 1 0 7952 0 -1 14112
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_138
timestamp 1698175906
transform 1 0 8400 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_142
timestamp 1698175906
transform 1 0 8624 0 -1 14112
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_158
timestamp 1698175906
transform 1 0 9520 0 -1 14112
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_166
timestamp 1698175906
transform 1 0 9968 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_168
timestamp 1698175906
transform 1 0 10080 0 -1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_198
timestamp 1698175906
transform 1 0 11760 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_202
timestamp 1698175906
transform 1 0 11984 0 -1 14112
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_216
timestamp 1698175906
transform 1 0 12768 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_224
timestamp 1698175906
transform 1 0 13216 0 -1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_256
timestamp 1698175906
transform 1 0 15008 0 -1 14112
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_272
timestamp 1698175906
transform 1 0 15904 0 -1 14112
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_282
timestamp 1698175906
transform 1 0 16464 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_346
timestamp 1698175906
transform 1 0 20048 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_348
timestamp 1698175906
transform 1 0 20160 0 -1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_2
timestamp 1698175906
transform 1 0 784 0 1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698175906
transform 1 0 2576 0 1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_37
timestamp 1698175906
transform 1 0 2744 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_101
timestamp 1698175906
transform 1 0 6328 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_107
timestamp 1698175906
transform 1 0 6664 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_171
timestamp 1698175906
transform 1 0 10248 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_177
timestamp 1698175906
transform 1 0 10584 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_185
timestamp 1698175906
transform 1 0 11032 0 1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_217
timestamp 1698175906
transform 1 0 12824 0 1 14112
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_233
timestamp 1698175906
transform 1 0 13720 0 1 14112
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_241
timestamp 1698175906
transform 1 0 14168 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_247
timestamp 1698175906
transform 1 0 14504 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_311
timestamp 1698175906
transform 1 0 18088 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_317
timestamp 1698175906
transform 1 0 18424 0 1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_2
timestamp 1698175906
transform 1 0 784 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_66
timestamp 1698175906
transform 1 0 4368 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_72
timestamp 1698175906
transform 1 0 4704 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_136
timestamp 1698175906
transform 1 0 8288 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_142
timestamp 1698175906
transform 1 0 8624 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_206
timestamp 1698175906
transform 1 0 12208 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_212
timestamp 1698175906
transform 1 0 12544 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_276
timestamp 1698175906
transform 1 0 16128 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_282
timestamp 1698175906
transform 1 0 16464 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_346
timestamp 1698175906
transform 1 0 20048 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_348
timestamp 1698175906
transform 1 0 20160 0 -1 14896
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698175906
transform 1 0 784 0 1 14896
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698175906
transform 1 0 2576 0 1 14896
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_37
timestamp 1698175906
transform 1 0 2744 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_101
timestamp 1698175906
transform 1 0 6328 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_107
timestamp 1698175906
transform 1 0 6664 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_171
timestamp 1698175906
transform 1 0 10248 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_177
timestamp 1698175906
transform 1 0 10584 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_241
timestamp 1698175906
transform 1 0 14168 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_247
timestamp 1698175906
transform 1 0 14504 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_311
timestamp 1698175906
transform 1 0 18088 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_317
timestamp 1698175906
transform 1 0 18424 0 1 14896
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2
timestamp 1698175906
transform 1 0 784 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_66
timestamp 1698175906
transform 1 0 4368 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_72
timestamp 1698175906
transform 1 0 4704 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_136
timestamp 1698175906
transform 1 0 8288 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_142
timestamp 1698175906
transform 1 0 8624 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_206
timestamp 1698175906
transform 1 0 12208 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_212
timestamp 1698175906
transform 1 0 12544 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_276
timestamp 1698175906
transform 1 0 16128 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_282
timestamp 1698175906
transform 1 0 16464 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_346
timestamp 1698175906
transform 1 0 20048 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_348
timestamp 1698175906
transform 1 0 20160 0 -1 15680
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_2
timestamp 1698175906
transform 1 0 784 0 1 15680
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698175906
transform 1 0 2576 0 1 15680
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_37
timestamp 1698175906
transform 1 0 2744 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_101
timestamp 1698175906
transform 1 0 6328 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_107
timestamp 1698175906
transform 1 0 6664 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_171
timestamp 1698175906
transform 1 0 10248 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_177
timestamp 1698175906
transform 1 0 10584 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_241
timestamp 1698175906
transform 1 0 14168 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_247
timestamp 1698175906
transform 1 0 14504 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_311
timestamp 1698175906
transform 1 0 18088 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_317
timestamp 1698175906
transform 1 0 18424 0 1 15680
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2
timestamp 1698175906
transform 1 0 784 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_66
timestamp 1698175906
transform 1 0 4368 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_72
timestamp 1698175906
transform 1 0 4704 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_136
timestamp 1698175906
transform 1 0 8288 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_142
timestamp 1698175906
transform 1 0 8624 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_206
timestamp 1698175906
transform 1 0 12208 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_212
timestamp 1698175906
transform 1 0 12544 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_276
timestamp 1698175906
transform 1 0 16128 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_282
timestamp 1698175906
transform 1 0 16464 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_346
timestamp 1698175906
transform 1 0 20048 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_348
timestamp 1698175906
transform 1 0 20160 0 -1 16464
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698175906
transform 1 0 784 0 1 16464
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698175906
transform 1 0 2576 0 1 16464
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_37
timestamp 1698175906
transform 1 0 2744 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_101
timestamp 1698175906
transform 1 0 6328 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_107
timestamp 1698175906
transform 1 0 6664 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_171
timestamp 1698175906
transform 1 0 10248 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_177
timestamp 1698175906
transform 1 0 10584 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_241
timestamp 1698175906
transform 1 0 14168 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_247
timestamp 1698175906
transform 1 0 14504 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_311
timestamp 1698175906
transform 1 0 18088 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_317
timestamp 1698175906
transform 1 0 18424 0 1 16464
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_2
timestamp 1698175906
transform 1 0 784 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_66
timestamp 1698175906
transform 1 0 4368 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_72
timestamp 1698175906
transform 1 0 4704 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_136
timestamp 1698175906
transform 1 0 8288 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_142
timestamp 1698175906
transform 1 0 8624 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_206
timestamp 1698175906
transform 1 0 12208 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_212
timestamp 1698175906
transform 1 0 12544 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_276
timestamp 1698175906
transform 1 0 16128 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_282
timestamp 1698175906
transform 1 0 16464 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_346
timestamp 1698175906
transform 1 0 20048 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_348
timestamp 1698175906
transform 1 0 20160 0 -1 17248
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698175906
transform 1 0 784 0 1 17248
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698175906
transform 1 0 2576 0 1 17248
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_37
timestamp 1698175906
transform 1 0 2744 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_101
timestamp 1698175906
transform 1 0 6328 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_107
timestamp 1698175906
transform 1 0 6664 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_171
timestamp 1698175906
transform 1 0 10248 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_177
timestamp 1698175906
transform 1 0 10584 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_241
timestamp 1698175906
transform 1 0 14168 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_247
timestamp 1698175906
transform 1 0 14504 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_311
timestamp 1698175906
transform 1 0 18088 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_317
timestamp 1698175906
transform 1 0 18424 0 1 17248
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2
timestamp 1698175906
transform 1 0 784 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1698175906
transform 1 0 4368 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_72
timestamp 1698175906
transform 1 0 4704 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_136
timestamp 1698175906
transform 1 0 8288 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_142
timestamp 1698175906
transform 1 0 8624 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_206
timestamp 1698175906
transform 1 0 12208 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_212
timestamp 1698175906
transform 1 0 12544 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_276
timestamp 1698175906
transform 1 0 16128 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_282
timestamp 1698175906
transform 1 0 16464 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_346
timestamp 1698175906
transform 1 0 20048 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_348
timestamp 1698175906
transform 1 0 20160 0 -1 18032
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_2
timestamp 1698175906
transform 1 0 784 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698175906
transform 1 0 2576 0 1 18032
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_37
timestamp 1698175906
transform 1 0 2744 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_101
timestamp 1698175906
transform 1 0 6328 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_107
timestamp 1698175906
transform 1 0 6664 0 1 18032
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_123
timestamp 1698175906
transform 1 0 7560 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_153
timestamp 1698175906
transform 1 0 9240 0 1 18032
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_169
timestamp 1698175906
transform 1 0 10136 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_173
timestamp 1698175906
transform 1 0 10360 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_177
timestamp 1698175906
transform 1 0 10584 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_241
timestamp 1698175906
transform 1 0 14168 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_247
timestamp 1698175906
transform 1 0 14504 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_311
timestamp 1698175906
transform 1 0 18088 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_317
timestamp 1698175906
transform 1 0 18424 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_2
timestamp 1698175906
transform 1 0 784 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_66
timestamp 1698175906
transform 1 0 4368 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_72
timestamp 1698175906
transform 1 0 4704 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_136
timestamp 1698175906
transform 1 0 8288 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_142
timestamp 1698175906
transform 1 0 8624 0 -1 18816
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_150
timestamp 1698175906
transform 1 0 9072 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_154
timestamp 1698175906
transform 1 0 9296 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_156
timestamp 1698175906
transform 1 0 9408 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_183
timestamp 1698175906
transform 1 0 10920 0 -1 18816
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_199
timestamp 1698175906
transform 1 0 11816 0 -1 18816
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_207
timestamp 1698175906
transform 1 0 12264 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_209
timestamp 1698175906
transform 1 0 12376 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_212
timestamp 1698175906
transform 1 0 12544 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_216
timestamp 1698175906
transform 1 0 12768 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_243
timestamp 1698175906
transform 1 0 14280 0 -1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_275
timestamp 1698175906
transform 1 0 16072 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_279
timestamp 1698175906
transform 1 0 16296 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_282
timestamp 1698175906
transform 1 0 16464 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_346
timestamp 1698175906
transform 1 0 20048 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_348
timestamp 1698175906
transform 1 0 20160 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_2
timestamp 1698175906
transform 1 0 784 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_36
timestamp 1698175906
transform 1 0 2688 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_70
timestamp 1698175906
transform 1 0 4592 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_104
timestamp 1698175906
transform 1 0 6496 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_138
timestamp 1698175906
transform 1 0 8400 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_142
timestamp 1698175906
transform 1 0 8624 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_172
timestamp 1698175906
transform 1 0 10304 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_176
timestamp 1698175906
transform 1 0 10528 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_232
timestamp 1698175906
transform 1 0 13664 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_236
timestamp 1698175906
transform 1 0 13888 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_266
timestamp 1698175906
transform 1 0 15568 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_270
timestamp 1698175906
transform 1 0 15792 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_274
timestamp 1698175906
transform 1 0 16016 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_308
timestamp 1698175906
transform 1 0 17920 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_342
timestamp 1698175906
transform 1 0 19824 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_346
timestamp 1698175906
transform 1 0 20048 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_348
timestamp 1698175906
transform 1 0 20160 0 1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18760 0 -1 11760
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output2
timestamp 1698175906
transform -1 0 2240 0 1 11760
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output3
timestamp 1698175906
transform 1 0 8736 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output4
timestamp 1698175906
transform 1 0 18760 0 -1 12544
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output5
timestamp 1698175906
transform 1 0 18760 0 -1 10192
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output6
timestamp 1698175906
transform 1 0 14112 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output7
timestamp 1698175906
transform -1 0 2240 0 -1 13328
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output8
timestamp 1698175906
transform 1 0 18760 0 1 7840
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output9
timestamp 1698175906
transform 1 0 12824 0 -1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output10
timestamp 1698175906
transform 1 0 18760 0 1 9408
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output11
timestamp 1698175906
transform 1 0 8736 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output12
timestamp 1698175906
transform 1 0 7784 0 1 18032
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output13
timestamp 1698175906
transform 1 0 12208 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output14
timestamp 1698175906
transform 1 0 10640 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output15
timestamp 1698175906
transform 1 0 12544 0 -1 2352
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output16
timestamp 1698175906
transform -1 0 2240 0 -1 8624
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output17
timestamp 1698175906
transform -1 0 2240 0 1 7840
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output18
timestamp 1698175906
transform 1 0 8792 0 1 2352
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output19
timestamp 1698175906
transform 1 0 9800 0 -1 2352
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output20
timestamp 1698175906
transform 1 0 18760 0 1 11760
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output21
timestamp 1698175906
transform -1 0 2240 0 -1 11760
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output22
timestamp 1698175906
transform 1 0 10640 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output23
timestamp 1698175906
transform 1 0 18760 0 -1 8624
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output24
timestamp 1698175906
transform 1 0 12208 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output25
timestamp 1698175906
transform 1 0 18760 0 1 13328
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output26
timestamp 1698175906
transform 1 0 9464 0 -1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_45 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 672 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698175906
transform -1 0 20328 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_46
timestamp 1698175906
transform 1 0 672 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698175906
transform -1 0 20328 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_47
timestamp 1698175906
transform 1 0 672 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698175906
transform -1 0 20328 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_48
timestamp 1698175906
transform 1 0 672 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698175906
transform -1 0 20328 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_49
timestamp 1698175906
transform 1 0 672 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698175906
transform -1 0 20328 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_50
timestamp 1698175906
transform 1 0 672 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698175906
transform -1 0 20328 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_51
timestamp 1698175906
transform 1 0 672 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698175906
transform -1 0 20328 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_52
timestamp 1698175906
transform 1 0 672 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698175906
transform -1 0 20328 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_53
timestamp 1698175906
transform 1 0 672 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698175906
transform -1 0 20328 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_54
timestamp 1698175906
transform 1 0 672 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698175906
transform -1 0 20328 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_55
timestamp 1698175906
transform 1 0 672 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698175906
transform -1 0 20328 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_56
timestamp 1698175906
transform 1 0 672 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698175906
transform -1 0 20328 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_57
timestamp 1698175906
transform 1 0 672 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698175906
transform -1 0 20328 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_58
timestamp 1698175906
transform 1 0 672 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698175906
transform -1 0 20328 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_59
timestamp 1698175906
transform 1 0 672 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698175906
transform -1 0 20328 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_60
timestamp 1698175906
transform 1 0 672 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698175906
transform -1 0 20328 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_61
timestamp 1698175906
transform 1 0 672 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698175906
transform -1 0 20328 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_62
timestamp 1698175906
transform 1 0 672 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698175906
transform -1 0 20328 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_63
timestamp 1698175906
transform 1 0 672 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698175906
transform -1 0 20328 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_64
timestamp 1698175906
transform 1 0 672 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698175906
transform -1 0 20328 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_65
timestamp 1698175906
transform 1 0 672 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698175906
transform -1 0 20328 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_66
timestamp 1698175906
transform 1 0 672 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698175906
transform -1 0 20328 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_67
timestamp 1698175906
transform 1 0 672 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698175906
transform -1 0 20328 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_68
timestamp 1698175906
transform 1 0 672 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698175906
transform -1 0 20328 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_69
timestamp 1698175906
transform 1 0 672 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698175906
transform -1 0 20328 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_70
timestamp 1698175906
transform 1 0 672 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698175906
transform -1 0 20328 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_71
timestamp 1698175906
transform 1 0 672 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698175906
transform -1 0 20328 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_72
timestamp 1698175906
transform 1 0 672 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698175906
transform -1 0 20328 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_73
timestamp 1698175906
transform 1 0 672 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698175906
transform -1 0 20328 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_74
timestamp 1698175906
transform 1 0 672 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698175906
transform -1 0 20328 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_75
timestamp 1698175906
transform 1 0 672 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698175906
transform -1 0 20328 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_76
timestamp 1698175906
transform 1 0 672 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698175906
transform -1 0 20328 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_77
timestamp 1698175906
transform 1 0 672 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698175906
transform -1 0 20328 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_78
timestamp 1698175906
transform 1 0 672 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698175906
transform -1 0 20328 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_79
timestamp 1698175906
transform 1 0 672 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698175906
transform -1 0 20328 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_80
timestamp 1698175906
transform 1 0 672 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698175906
transform -1 0 20328 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_81
timestamp 1698175906
transform 1 0 672 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698175906
transform -1 0 20328 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_82
timestamp 1698175906
transform 1 0 672 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698175906
transform -1 0 20328 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_83
timestamp 1698175906
transform 1 0 672 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698175906
transform -1 0 20328 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_84
timestamp 1698175906
transform 1 0 672 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698175906
transform -1 0 20328 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_85
timestamp 1698175906
transform 1 0 672 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698175906
transform -1 0 20328 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_86
timestamp 1698175906
transform 1 0 672 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698175906
transform -1 0 20328 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_87
timestamp 1698175906
transform 1 0 672 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698175906
transform -1 0 20328 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_88
timestamp 1698175906
transform 1 0 672 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698175906
transform -1 0 20328 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_89
timestamp 1698175906
transform 1 0 672 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698175906
transform -1 0 20328 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_90 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 2576 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_91
timestamp 1698175906
transform 1 0 4480 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_92
timestamp 1698175906
transform 1 0 6384 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_93
timestamp 1698175906
transform 1 0 8288 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_94
timestamp 1698175906
transform 1 0 10192 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_95
timestamp 1698175906
transform 1 0 12096 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_96
timestamp 1698175906
transform 1 0 14000 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_97
timestamp 1698175906
transform 1 0 15904 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_98
timestamp 1698175906
transform 1 0 17808 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_99
timestamp 1698175906
transform 1 0 19712 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_100
timestamp 1698175906
transform 1 0 4592 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_101
timestamp 1698175906
transform 1 0 8512 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_102
timestamp 1698175906
transform 1 0 12432 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_103
timestamp 1698175906
transform 1 0 16352 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_104
timestamp 1698175906
transform 1 0 2632 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_105
timestamp 1698175906
transform 1 0 6552 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_106
timestamp 1698175906
transform 1 0 10472 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_107
timestamp 1698175906
transform 1 0 14392 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_108
timestamp 1698175906
transform 1 0 18312 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_109
timestamp 1698175906
transform 1 0 4592 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_110
timestamp 1698175906
transform 1 0 8512 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_111
timestamp 1698175906
transform 1 0 12432 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_112
timestamp 1698175906
transform 1 0 16352 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_113
timestamp 1698175906
transform 1 0 2632 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_114
timestamp 1698175906
transform 1 0 6552 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_115
timestamp 1698175906
transform 1 0 10472 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_116
timestamp 1698175906
transform 1 0 14392 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_117
timestamp 1698175906
transform 1 0 18312 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_118
timestamp 1698175906
transform 1 0 4592 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_119
timestamp 1698175906
transform 1 0 8512 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_120
timestamp 1698175906
transform 1 0 12432 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_121
timestamp 1698175906
transform 1 0 16352 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_122
timestamp 1698175906
transform 1 0 2632 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_123
timestamp 1698175906
transform 1 0 6552 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_124
timestamp 1698175906
transform 1 0 10472 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_125
timestamp 1698175906
transform 1 0 14392 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_126
timestamp 1698175906
transform 1 0 18312 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_127
timestamp 1698175906
transform 1 0 4592 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_128
timestamp 1698175906
transform 1 0 8512 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_129
timestamp 1698175906
transform 1 0 12432 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_130
timestamp 1698175906
transform 1 0 16352 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_131
timestamp 1698175906
transform 1 0 2632 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_132
timestamp 1698175906
transform 1 0 6552 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_133
timestamp 1698175906
transform 1 0 10472 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_134
timestamp 1698175906
transform 1 0 14392 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_135
timestamp 1698175906
transform 1 0 18312 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_136
timestamp 1698175906
transform 1 0 4592 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_137
timestamp 1698175906
transform 1 0 8512 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_138
timestamp 1698175906
transform 1 0 12432 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_139
timestamp 1698175906
transform 1 0 16352 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_140
timestamp 1698175906
transform 1 0 2632 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_141
timestamp 1698175906
transform 1 0 6552 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_142
timestamp 1698175906
transform 1 0 10472 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_143
timestamp 1698175906
transform 1 0 14392 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_144
timestamp 1698175906
transform 1 0 18312 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_145
timestamp 1698175906
transform 1 0 4592 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_146
timestamp 1698175906
transform 1 0 8512 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_147
timestamp 1698175906
transform 1 0 12432 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_148
timestamp 1698175906
transform 1 0 16352 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_149
timestamp 1698175906
transform 1 0 2632 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_150
timestamp 1698175906
transform 1 0 6552 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_151
timestamp 1698175906
transform 1 0 10472 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_152
timestamp 1698175906
transform 1 0 14392 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_153
timestamp 1698175906
transform 1 0 18312 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_154
timestamp 1698175906
transform 1 0 4592 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_155
timestamp 1698175906
transform 1 0 8512 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_156
timestamp 1698175906
transform 1 0 12432 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_157
timestamp 1698175906
transform 1 0 16352 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_158
timestamp 1698175906
transform 1 0 2632 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_159
timestamp 1698175906
transform 1 0 6552 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_160
timestamp 1698175906
transform 1 0 10472 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_161
timestamp 1698175906
transform 1 0 14392 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_162
timestamp 1698175906
transform 1 0 18312 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_163
timestamp 1698175906
transform 1 0 4592 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_164
timestamp 1698175906
transform 1 0 8512 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_165
timestamp 1698175906
transform 1 0 12432 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_166
timestamp 1698175906
transform 1 0 16352 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_167
timestamp 1698175906
transform 1 0 2632 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_168
timestamp 1698175906
transform 1 0 6552 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_169
timestamp 1698175906
transform 1 0 10472 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_170
timestamp 1698175906
transform 1 0 14392 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_171
timestamp 1698175906
transform 1 0 18312 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_172
timestamp 1698175906
transform 1 0 4592 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_173
timestamp 1698175906
transform 1 0 8512 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_174
timestamp 1698175906
transform 1 0 12432 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_175
timestamp 1698175906
transform 1 0 16352 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_176
timestamp 1698175906
transform 1 0 2632 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_177
timestamp 1698175906
transform 1 0 6552 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_178
timestamp 1698175906
transform 1 0 10472 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_179
timestamp 1698175906
transform 1 0 14392 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_180
timestamp 1698175906
transform 1 0 18312 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_181
timestamp 1698175906
transform 1 0 4592 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_182
timestamp 1698175906
transform 1 0 8512 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_183
timestamp 1698175906
transform 1 0 12432 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_184
timestamp 1698175906
transform 1 0 16352 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_185
timestamp 1698175906
transform 1 0 2632 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_186
timestamp 1698175906
transform 1 0 6552 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_187
timestamp 1698175906
transform 1 0 10472 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_188
timestamp 1698175906
transform 1 0 14392 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_189
timestamp 1698175906
transform 1 0 18312 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_190
timestamp 1698175906
transform 1 0 4592 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_191
timestamp 1698175906
transform 1 0 8512 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_192
timestamp 1698175906
transform 1 0 12432 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_193
timestamp 1698175906
transform 1 0 16352 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_194
timestamp 1698175906
transform 1 0 2632 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_195
timestamp 1698175906
transform 1 0 6552 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_196
timestamp 1698175906
transform 1 0 10472 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_197
timestamp 1698175906
transform 1 0 14392 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_198
timestamp 1698175906
transform 1 0 18312 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_199
timestamp 1698175906
transform 1 0 4592 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_200
timestamp 1698175906
transform 1 0 8512 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_201
timestamp 1698175906
transform 1 0 12432 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_202
timestamp 1698175906
transform 1 0 16352 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_203
timestamp 1698175906
transform 1 0 2632 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_204
timestamp 1698175906
transform 1 0 6552 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_205
timestamp 1698175906
transform 1 0 10472 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_206
timestamp 1698175906
transform 1 0 14392 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_207
timestamp 1698175906
transform 1 0 18312 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_208
timestamp 1698175906
transform 1 0 4592 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_209
timestamp 1698175906
transform 1 0 8512 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_210
timestamp 1698175906
transform 1 0 12432 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_211
timestamp 1698175906
transform 1 0 16352 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_212
timestamp 1698175906
transform 1 0 2632 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_213
timestamp 1698175906
transform 1 0 6552 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_214
timestamp 1698175906
transform 1 0 10472 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_215
timestamp 1698175906
transform 1 0 14392 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_216
timestamp 1698175906
transform 1 0 18312 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_217
timestamp 1698175906
transform 1 0 4592 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_218
timestamp 1698175906
transform 1 0 8512 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_219
timestamp 1698175906
transform 1 0 12432 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_220
timestamp 1698175906
transform 1 0 16352 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_221
timestamp 1698175906
transform 1 0 2632 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_222
timestamp 1698175906
transform 1 0 6552 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_223
timestamp 1698175906
transform 1 0 10472 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_224
timestamp 1698175906
transform 1 0 14392 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_225
timestamp 1698175906
transform 1 0 18312 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_226
timestamp 1698175906
transform 1 0 4592 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_227
timestamp 1698175906
transform 1 0 8512 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_228
timestamp 1698175906
transform 1 0 12432 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_229
timestamp 1698175906
transform 1 0 16352 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_230
timestamp 1698175906
transform 1 0 2632 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_231
timestamp 1698175906
transform 1 0 6552 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_232
timestamp 1698175906
transform 1 0 10472 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_233
timestamp 1698175906
transform 1 0 14392 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_234
timestamp 1698175906
transform 1 0 18312 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_235
timestamp 1698175906
transform 1 0 4592 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_236
timestamp 1698175906
transform 1 0 8512 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_237
timestamp 1698175906
transform 1 0 12432 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_238
timestamp 1698175906
transform 1 0 16352 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_239
timestamp 1698175906
transform 1 0 2632 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_240
timestamp 1698175906
transform 1 0 6552 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_241
timestamp 1698175906
transform 1 0 10472 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_242
timestamp 1698175906
transform 1 0 14392 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_243
timestamp 1698175906
transform 1 0 18312 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_244
timestamp 1698175906
transform 1 0 4592 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_245
timestamp 1698175906
transform 1 0 8512 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_246
timestamp 1698175906
transform 1 0 12432 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_247
timestamp 1698175906
transform 1 0 16352 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_248
timestamp 1698175906
transform 1 0 2632 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_249
timestamp 1698175906
transform 1 0 6552 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_250
timestamp 1698175906
transform 1 0 10472 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_251
timestamp 1698175906
transform 1 0 14392 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_252
timestamp 1698175906
transform 1 0 18312 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_253
timestamp 1698175906
transform 1 0 4592 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_254
timestamp 1698175906
transform 1 0 8512 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_255
timestamp 1698175906
transform 1 0 12432 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_256
timestamp 1698175906
transform 1 0 16352 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_257
timestamp 1698175906
transform 1 0 2632 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_258
timestamp 1698175906
transform 1 0 6552 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_259
timestamp 1698175906
transform 1 0 10472 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_260
timestamp 1698175906
transform 1 0 14392 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_261
timestamp 1698175906
transform 1 0 18312 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_262
timestamp 1698175906
transform 1 0 4592 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_263
timestamp 1698175906
transform 1 0 8512 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_264
timestamp 1698175906
transform 1 0 12432 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_265
timestamp 1698175906
transform 1 0 16352 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_266
timestamp 1698175906
transform 1 0 2632 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_267
timestamp 1698175906
transform 1 0 6552 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_268
timestamp 1698175906
transform 1 0 10472 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_269
timestamp 1698175906
transform 1 0 14392 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_270
timestamp 1698175906
transform 1 0 18312 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_271
timestamp 1698175906
transform 1 0 4592 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_272
timestamp 1698175906
transform 1 0 8512 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_273
timestamp 1698175906
transform 1 0 12432 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_274
timestamp 1698175906
transform 1 0 16352 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_275
timestamp 1698175906
transform 1 0 2632 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_276
timestamp 1698175906
transform 1 0 6552 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_277
timestamp 1698175906
transform 1 0 10472 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_278
timestamp 1698175906
transform 1 0 14392 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_279
timestamp 1698175906
transform 1 0 18312 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_280
timestamp 1698175906
transform 1 0 4592 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_281
timestamp 1698175906
transform 1 0 8512 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_282
timestamp 1698175906
transform 1 0 12432 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_283
timestamp 1698175906
transform 1 0 16352 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_284
timestamp 1698175906
transform 1 0 2632 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_285
timestamp 1698175906
transform 1 0 6552 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_286
timestamp 1698175906
transform 1 0 10472 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_287
timestamp 1698175906
transform 1 0 14392 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_288
timestamp 1698175906
transform 1 0 18312 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_289
timestamp 1698175906
transform 1 0 4592 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_290
timestamp 1698175906
transform 1 0 8512 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_291
timestamp 1698175906
transform 1 0 12432 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_292
timestamp 1698175906
transform 1 0 16352 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_293
timestamp 1698175906
transform 1 0 2576 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_294
timestamp 1698175906
transform 1 0 4480 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_295
timestamp 1698175906
transform 1 0 6384 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_296
timestamp 1698175906
transform 1 0 8288 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_297
timestamp 1698175906
transform 1 0 10192 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_298
timestamp 1698175906
transform 1 0 12096 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_299
timestamp 1698175906
transform 1 0 14000 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_300
timestamp 1698175906
transform 1 0 15904 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_301
timestamp 1698175906
transform 1 0 17808 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_302
timestamp 1698175906
transform 1 0 19712 0 1 18816
box -43 -43 155 435
<< labels >>
flabel metal3 s 0 13776 400 13832 0 FreeSans 224 0 0 0 clk
port 0 nsew signal input
flabel metal3 s 20600 11424 21000 11480 0 FreeSans 224 0 0 0 segm[0]
port 1 nsew signal tristate
flabel metal3 s 0 11760 400 11816 0 FreeSans 224 0 0 0 segm[10]
port 2 nsew signal tristate
flabel metal2 s 9072 0 9128 400 0 FreeSans 224 90 0 0 segm[11]
port 3 nsew signal tristate
flabel metal3 s 20600 12096 21000 12152 0 FreeSans 224 0 0 0 segm[12]
port 4 nsew signal tristate
flabel metal3 s 20600 9744 21000 9800 0 FreeSans 224 0 0 0 segm[13]
port 5 nsew signal tristate
flabel metal2 s 13104 20600 13160 21000 0 FreeSans 224 90 0 0 segm[1]
port 6 nsew signal tristate
flabel metal3 s 0 12768 400 12824 0 FreeSans 224 0 0 0 segm[2]
port 7 nsew signal tristate
flabel metal3 s 20600 7728 21000 7784 0 FreeSans 224 0 0 0 segm[3]
port 8 nsew signal tristate
flabel metal2 s 12768 20600 12824 21000 0 FreeSans 224 90 0 0 segm[4]
port 9 nsew signal tristate
flabel metal3 s 20600 9408 21000 9464 0 FreeSans 224 0 0 0 segm[5]
port 10 nsew signal tristate
flabel metal2 s 8736 20600 8792 21000 0 FreeSans 224 90 0 0 segm[6]
port 11 nsew signal tristate
flabel metal2 s 7728 20600 7784 21000 0 FreeSans 224 90 0 0 segm[7]
port 12 nsew signal tristate
flabel metal2 s 11424 20600 11480 21000 0 FreeSans 224 90 0 0 segm[8]
port 13 nsew signal tristate
flabel metal2 s 11088 20600 11144 21000 0 FreeSans 224 90 0 0 segm[9]
port 14 nsew signal tristate
flabel metal2 s 12096 0 12152 400 0 FreeSans 224 90 0 0 sel[0]
port 15 nsew signal tristate
flabel metal3 s 0 8064 400 8120 0 FreeSans 224 0 0 0 sel[10]
port 16 nsew signal tristate
flabel metal3 s 0 7728 400 7784 0 FreeSans 224 0 0 0 sel[11]
port 17 nsew signal tristate
flabel metal2 s 8736 0 8792 400 0 FreeSans 224 90 0 0 sel[1]
port 18 nsew signal tristate
flabel metal2 s 9744 0 9800 400 0 FreeSans 224 90 0 0 sel[2]
port 19 nsew signal tristate
flabel metal3 s 20600 11760 21000 11816 0 FreeSans 224 0 0 0 sel[3]
port 20 nsew signal tristate
flabel metal3 s 0 11424 400 11480 0 FreeSans 224 0 0 0 sel[4]
port 21 nsew signal tristate
flabel metal2 s 11088 0 11144 400 0 FreeSans 224 90 0 0 sel[5]
port 22 nsew signal tristate
flabel metal3 s 20600 8064 21000 8120 0 FreeSans 224 0 0 0 sel[6]
port 23 nsew signal tristate
flabel metal2 s 11424 0 11480 400 0 FreeSans 224 90 0 0 sel[7]
port 24 nsew signal tristate
flabel metal3 s 20600 13104 21000 13160 0 FreeSans 224 0 0 0 sel[8]
port 25 nsew signal tristate
flabel metal2 s 9408 20600 9464 21000 0 FreeSans 224 90 0 0 sel[9]
port 26 nsew signal tristate
flabel metal4 s 2224 1538 2384 19238 0 FreeSans 640 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 17584 1538 17744 19238 0 FreeSans 640 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 9904 1538 10064 19238 0 FreeSans 640 90 0 0 vss
port 28 nsew ground bidirectional
rlabel metal1 10500 19208 10500 19208 0 vdd
rlabel metal1 10500 18816 10500 18816 0 vss
rlabel metal2 12292 12936 12292 12936 0 _000_
rlabel metal2 13888 7700 13888 7700 0 _001_
rlabel metal2 13916 11368 13916 11368 0 _002_
rlabel metal2 10500 7616 10500 7616 0 _003_
rlabel metal2 9100 12572 9100 12572 0 _004_
rlabel metal2 10724 8064 10724 8064 0 _005_
rlabel metal2 11228 10836 11228 10836 0 _006_
rlabel metal2 12460 11536 12460 11536 0 _007_
rlabel metal2 12516 9016 12516 9016 0 _008_
rlabel metal2 7532 11368 7532 11368 0 _009_
rlabel metal2 8932 6636 8932 6636 0 _010_
rlabel metal2 7364 7280 7364 7280 0 _011_
rlabel metal2 11984 7308 11984 7308 0 _012_
rlabel metal2 11620 13440 11620 13440 0 _013_
rlabel metal2 10612 14000 10612 14000 0 _014_
rlabel metal2 10108 13356 10108 13356 0 _015_
rlabel metal2 13300 11984 13300 11984 0 _016_
rlabel metal2 14112 6916 14112 6916 0 _017_
rlabel metal2 14812 9800 14812 9800 0 _018_
rlabel metal2 14252 9324 14252 9324 0 _019_
rlabel metal2 11284 7028 11284 7028 0 _020_
rlabel metal2 6748 7672 6748 7672 0 _021_
rlabel metal2 6972 8232 6972 8232 0 _022_
rlabel metal2 6244 12880 6244 12880 0 _023_
rlabel metal2 8260 13020 8260 13020 0 _024_
rlabel metal2 7140 13748 7140 13748 0 _025_
rlabel metal2 6636 10892 6636 10892 0 _026_
rlabel metal2 7924 8148 7924 8148 0 _027_
rlabel metal2 10304 12628 10304 12628 0 _028_
rlabel metal2 9772 11704 9772 11704 0 _029_
rlabel metal2 9044 12992 9044 12992 0 _030_
rlabel metal2 11172 12964 11172 12964 0 _031_
rlabel metal2 11452 13552 11452 13552 0 _032_
rlabel metal2 8372 11060 8372 11060 0 _033_
rlabel metal2 8960 13244 8960 13244 0 _034_
rlabel metal2 9380 12880 9380 12880 0 _035_
rlabel metal2 6860 10178 6860 10178 0 _036_
rlabel metal2 10556 12152 10556 12152 0 _037_
rlabel metal2 12208 11900 12208 11900 0 _038_
rlabel metal2 11452 9240 11452 9240 0 _039_
rlabel metal2 8596 11284 8596 11284 0 _040_
rlabel metal3 8204 8428 8204 8428 0 _041_
rlabel metal2 9156 8456 9156 8456 0 _042_
rlabel metal2 7980 11228 7980 11228 0 _043_
rlabel metal2 7644 11312 7644 11312 0 _044_
rlabel metal2 9604 8036 9604 8036 0 _045_
rlabel metal2 8988 7056 8988 7056 0 _046_
rlabel metal2 9100 7252 9100 7252 0 _047_
rlabel metal2 8764 7420 8764 7420 0 _048_
rlabel metal2 11900 8568 11900 8568 0 _049_
rlabel metal2 11788 7868 11788 7868 0 _050_
rlabel metal2 11564 13664 11564 13664 0 _051_
rlabel metal2 11228 12656 11228 12656 0 _052_
rlabel metal2 11284 12320 11284 12320 0 _053_
rlabel metal2 10948 14280 10948 14280 0 _054_
rlabel metal2 10332 13132 10332 13132 0 _055_
rlabel metal2 10388 13552 10388 13552 0 _056_
rlabel metal2 13384 10668 13384 10668 0 _057_
rlabel metal2 13468 11732 13468 11732 0 _058_
rlabel metal3 14532 7980 14532 7980 0 _059_
rlabel metal2 15092 9688 15092 9688 0 _060_
rlabel metal2 13692 9884 13692 9884 0 _061_
rlabel metal2 14140 9688 14140 9688 0 _062_
rlabel metal2 11368 7364 11368 7364 0 _063_
rlabel metal3 7672 11060 7672 11060 0 _064_
rlabel metal2 7252 8092 7252 8092 0 _065_
rlabel metal2 6860 7644 6860 7644 0 _066_
rlabel metal2 7644 12600 7644 12600 0 _067_
rlabel metal2 8764 12824 8764 12824 0 _068_
rlabel metal3 8260 11228 8260 11228 0 _069_
rlabel metal3 7532 12460 7532 12460 0 _070_
rlabel metal3 6860 12684 6860 12684 0 _071_
rlabel metal3 8764 13132 8764 13132 0 _072_
rlabel metal3 7644 13188 7644 13188 0 _073_
rlabel metal2 6972 11256 6972 11256 0 _074_
rlabel metal2 6860 11592 6860 11592 0 _075_
rlabel metal2 8316 8624 8316 8624 0 _076_
rlabel metal2 9324 8232 9324 8232 0 _077_
rlabel metal3 8932 8092 8932 8092 0 _078_
rlabel metal2 11844 9352 11844 9352 0 _079_
rlabel metal2 11928 10836 11928 10836 0 _080_
rlabel metal2 13076 11228 13076 11228 0 _081_
rlabel metal2 10892 11788 10892 11788 0 _082_
rlabel metal2 11844 12040 11844 12040 0 _083_
rlabel metal2 10164 11228 10164 11228 0 _084_
rlabel metal2 14084 11760 14084 11760 0 _085_
rlabel metal3 12768 12740 12768 12740 0 _086_
rlabel metal2 9296 9996 9296 9996 0 _087_
rlabel metal2 10668 10458 10668 10458 0 _088_
rlabel metal2 8316 10430 8316 10430 0 _089_
rlabel metal3 10612 10808 10612 10808 0 _090_
rlabel metal2 11396 10780 11396 10780 0 _091_
rlabel metal3 12824 10780 12824 10780 0 _092_
rlabel metal2 10948 11088 10948 11088 0 _093_
rlabel metal2 10948 13104 10948 13104 0 _094_
rlabel metal2 11676 10892 11676 10892 0 _095_
rlabel metal3 8932 9156 8932 9156 0 _096_
rlabel metal2 8820 10920 8820 10920 0 _097_
rlabel metal2 13076 9856 13076 9856 0 _098_
rlabel metal2 14308 9492 14308 9492 0 _099_
rlabel metal2 14532 8092 14532 8092 0 _100_
rlabel metal3 10948 7644 10948 7644 0 _101_
rlabel metal2 11648 11508 11648 11508 0 _102_
rlabel metal2 11004 9436 11004 9436 0 _103_
rlabel metal2 11060 11424 11060 11424 0 _104_
rlabel metal2 13860 8400 13860 8400 0 _105_
rlabel metal3 12180 9604 12180 9604 0 _106_
rlabel metal2 13636 9660 13636 9660 0 _107_
rlabel metal3 14028 9604 14028 9604 0 _108_
rlabel metal2 10108 11340 10108 11340 0 _109_
rlabel metal2 11004 11452 11004 11452 0 _110_
rlabel metal2 11732 11200 11732 11200 0 _111_
rlabel metal2 14224 11284 14224 11284 0 _112_
rlabel metal2 13664 11116 13664 11116 0 _113_
rlabel metal2 11116 8652 11116 8652 0 _114_
rlabel metal2 11116 8932 11116 8932 0 _115_
rlabel metal2 10332 8120 10332 8120 0 _116_
rlabel metal2 10780 7392 10780 7392 0 _117_
rlabel metal3 1239 13804 1239 13804 0 clk
rlabel metal3 11732 10108 11732 10108 0 clknet_0_clk
rlabel metal2 10220 6664 10220 6664 0 clknet_1_0__leaf_clk
rlabel metal3 11116 13916 11116 13916 0 clknet_1_1__leaf_clk
rlabel metal2 7112 9604 7112 9604 0 dut34.count\[0\]
rlabel metal2 7056 9940 7056 9940 0 dut34.count\[1\]
rlabel metal3 10528 11060 10528 11060 0 dut34.count\[2\]
rlabel metal3 10920 10444 10920 10444 0 dut34.count\[3\]
rlabel metal2 15092 11312 15092 11312 0 net1
rlabel metal2 15484 9716 15484 9716 0 net10
rlabel metal2 8708 13356 8708 13356 0 net11
rlabel metal2 7700 13496 7700 13496 0 net12
rlabel metal3 11984 13860 11984 13860 0 net13
rlabel metal2 10836 13748 10836 13748 0 net14
rlabel metal2 12628 3178 12628 3178 0 net15
rlabel metal2 2156 8288 2156 8288 0 net16
rlabel metal2 5628 8092 5628 8092 0 net17
rlabel metal2 8428 6328 8428 6328 0 net18
rlabel metal2 9856 2156 9856 2156 0 net19
rlabel metal2 5572 11340 5572 11340 0 net2
rlabel metal3 15694 11620 15694 11620 0 net20
rlabel metal2 6076 11536 6076 11536 0 net21
rlabel metal2 10836 6972 10836 6972 0 net22
rlabel metal2 14952 7588 14952 7588 0 net23
rlabel metal2 12292 2982 12292 2982 0 net24
rlabel metal2 14084 13104 14084 13104 0 net25
rlabel metal2 9716 13160 9716 13160 0 net26
rlabel metal2 8820 2982 8820 2982 0 net3
rlabel metal2 15316 12124 15316 12124 0 net4
rlabel metal2 15316 9576 15316 9576 0 net5
rlabel metal3 13720 14028 13720 14028 0 net6
rlabel metal2 2156 13104 2156 13104 0 net7
rlabel metal2 15176 6804 15176 6804 0 net8
rlabel metal2 12684 14000 12684 14000 0 net9
rlabel metal3 20321 11452 20321 11452 0 segm[0]
rlabel metal3 679 11788 679 11788 0 segm[10]
rlabel metal2 9100 1099 9100 1099 0 segm[11]
rlabel metal2 20020 12180 20020 12180 0 segm[12]
rlabel metal2 20020 9828 20020 9828 0 segm[13]
rlabel metal2 13132 19873 13132 19873 0 segm[1]
rlabel metal3 679 12796 679 12796 0 segm[2]
rlabel metal2 20020 7924 20020 7924 0 segm[3]
rlabel metal2 12796 19957 12796 19957 0 segm[4]
rlabel metal2 20020 9548 20020 9548 0 segm[5]
rlabel metal2 8764 19873 8764 19873 0 segm[6]
rlabel metal2 7756 19481 7756 19481 0 segm[7]
rlabel metal2 11452 19873 11452 19873 0 segm[8]
rlabel metal2 11116 19873 11116 19873 0 segm[9]
rlabel metal2 12124 1211 12124 1211 0 sel[0]
rlabel metal3 679 8092 679 8092 0 sel[10]
rlabel metal3 707 7756 707 7756 0 sel[11]
rlabel metal2 8764 1491 8764 1491 0 sel[1]
rlabel metal2 9772 1211 9772 1211 0 sel[2]
rlabel metal2 20020 11900 20020 11900 0 sel[3]
rlabel metal3 679 11452 679 11452 0 sel[4]
rlabel metal2 11116 1015 11116 1015 0 sel[5]
rlabel metal2 19964 8232 19964 8232 0 sel[6]
rlabel metal2 11452 1099 11452 1099 0 sel[7]
rlabel metal2 20020 13356 20020 13356 0 sel[8]
rlabel metal3 9744 18732 9744 18732 0 sel[9]
<< properties >>
string FIXED_BBOX 0 0 21000 21000
<< end >>
