magic
tech gf180mcuD
magscale 1 5
timestamp 1699642381
<< metal1 >>
rect 672 19221 20328 19238
rect 672 19195 2239 19221
rect 2265 19195 2291 19221
rect 2317 19195 2343 19221
rect 2369 19195 17599 19221
rect 17625 19195 17651 19221
rect 17677 19195 17703 19221
rect 17729 19195 20328 19221
rect 672 19178 20328 19195
rect 9311 19137 9337 19143
rect 9311 19105 9337 19111
rect 10879 19137 10905 19143
rect 10879 19105 10905 19111
rect 12783 19137 12809 19143
rect 12783 19105 12809 19111
rect 8801 18999 8807 19025
rect 8833 18999 8839 19025
rect 10369 18999 10375 19025
rect 10401 18999 10407 19025
rect 12273 18999 12279 19025
rect 12305 18999 12311 19025
rect 672 18829 20328 18846
rect 672 18803 9919 18829
rect 9945 18803 9971 18829
rect 9997 18803 10023 18829
rect 10049 18803 20328 18829
rect 672 18786 20328 18803
rect 10039 18745 10065 18751
rect 10039 18713 10065 18719
rect 13119 18745 13145 18751
rect 13119 18713 13145 18719
rect 9529 18607 9535 18633
rect 9561 18607 9567 18633
rect 12609 18607 12615 18633
rect 12641 18607 12647 18633
rect 672 18437 20328 18454
rect 672 18411 2239 18437
rect 2265 18411 2291 18437
rect 2317 18411 2343 18437
rect 2369 18411 17599 18437
rect 17625 18411 17651 18437
rect 17677 18411 17703 18437
rect 17729 18411 20328 18437
rect 672 18394 20328 18411
rect 672 18045 20328 18062
rect 672 18019 9919 18045
rect 9945 18019 9971 18045
rect 9997 18019 10023 18045
rect 10049 18019 20328 18045
rect 672 18002 20328 18019
rect 672 17653 20328 17670
rect 672 17627 2239 17653
rect 2265 17627 2291 17653
rect 2317 17627 2343 17653
rect 2369 17627 17599 17653
rect 17625 17627 17651 17653
rect 17677 17627 17703 17653
rect 17729 17627 20328 17653
rect 672 17610 20328 17627
rect 672 17261 20328 17278
rect 672 17235 9919 17261
rect 9945 17235 9971 17261
rect 9997 17235 10023 17261
rect 10049 17235 20328 17261
rect 672 17218 20328 17235
rect 672 16869 20328 16886
rect 672 16843 2239 16869
rect 2265 16843 2291 16869
rect 2317 16843 2343 16869
rect 2369 16843 17599 16869
rect 17625 16843 17651 16869
rect 17677 16843 17703 16869
rect 17729 16843 20328 16869
rect 672 16826 20328 16843
rect 672 16477 20328 16494
rect 672 16451 9919 16477
rect 9945 16451 9971 16477
rect 9997 16451 10023 16477
rect 10049 16451 20328 16477
rect 672 16434 20328 16451
rect 672 16085 20328 16102
rect 672 16059 2239 16085
rect 2265 16059 2291 16085
rect 2317 16059 2343 16085
rect 2369 16059 17599 16085
rect 17625 16059 17651 16085
rect 17677 16059 17703 16085
rect 17729 16059 20328 16085
rect 672 16042 20328 16059
rect 672 15693 20328 15710
rect 672 15667 9919 15693
rect 9945 15667 9971 15693
rect 9997 15667 10023 15693
rect 10049 15667 20328 15693
rect 672 15650 20328 15667
rect 672 15301 20328 15318
rect 672 15275 2239 15301
rect 2265 15275 2291 15301
rect 2317 15275 2343 15301
rect 2369 15275 17599 15301
rect 17625 15275 17651 15301
rect 17677 15275 17703 15301
rect 17729 15275 20328 15301
rect 672 15258 20328 15275
rect 672 14909 20328 14926
rect 672 14883 9919 14909
rect 9945 14883 9971 14909
rect 9997 14883 10023 14909
rect 10049 14883 20328 14909
rect 672 14866 20328 14883
rect 672 14517 20328 14534
rect 672 14491 2239 14517
rect 2265 14491 2291 14517
rect 2317 14491 2343 14517
rect 2369 14491 17599 14517
rect 17625 14491 17651 14517
rect 17677 14491 17703 14517
rect 17729 14491 20328 14517
rect 672 14474 20328 14491
rect 10151 14265 10177 14271
rect 10151 14233 10177 14239
rect 10207 14265 10233 14271
rect 10207 14233 10233 14239
rect 10879 14265 10905 14271
rect 10879 14233 10905 14239
rect 10935 14265 10961 14271
rect 10935 14233 10961 14239
rect 10039 14209 10065 14215
rect 10039 14177 10065 14183
rect 11047 14209 11073 14215
rect 11047 14177 11073 14183
rect 672 14125 20328 14142
rect 672 14099 9919 14125
rect 9945 14099 9971 14125
rect 9997 14099 10023 14125
rect 10049 14099 20328 14125
rect 672 14082 20328 14099
rect 8801 13903 8807 13929
rect 8833 13903 8839 13929
rect 10425 13903 10431 13929
rect 10457 13903 10463 13929
rect 8471 13873 8497 13879
rect 12111 13873 12137 13879
rect 9137 13847 9143 13873
rect 9169 13847 9175 13873
rect 10201 13847 10207 13873
rect 10233 13847 10239 13873
rect 10761 13847 10767 13873
rect 10793 13847 10799 13873
rect 11825 13847 11831 13873
rect 11857 13847 11863 13873
rect 8471 13841 8497 13847
rect 12111 13841 12137 13847
rect 672 13733 20328 13750
rect 672 13707 2239 13733
rect 2265 13707 2291 13733
rect 2317 13707 2343 13733
rect 2369 13707 17599 13733
rect 17625 13707 17651 13733
rect 17677 13707 17703 13733
rect 17729 13707 20328 13733
rect 672 13690 20328 13707
rect 9927 13593 9953 13599
rect 20007 13593 20033 13599
rect 9473 13567 9479 13593
rect 9505 13567 9511 13593
rect 12329 13567 12335 13593
rect 12361 13567 12367 13593
rect 14289 13567 14295 13593
rect 14321 13567 14327 13593
rect 9927 13561 9953 13567
rect 20007 13561 20033 13567
rect 9815 13537 9841 13543
rect 8073 13511 8079 13537
rect 8105 13511 8111 13537
rect 9815 13505 9841 13511
rect 10039 13537 10065 13543
rect 10039 13505 10065 13511
rect 10095 13537 10121 13543
rect 12559 13537 12585 13543
rect 10929 13511 10935 13537
rect 10961 13511 10967 13537
rect 12889 13511 12895 13537
rect 12921 13511 12927 13537
rect 18825 13511 18831 13537
rect 18857 13511 18863 13537
rect 10095 13505 10121 13511
rect 12559 13505 12585 13511
rect 9703 13481 9729 13487
rect 8409 13455 8415 13481
rect 8441 13455 8447 13481
rect 11265 13455 11271 13481
rect 11297 13455 11303 13481
rect 13225 13455 13231 13481
rect 13257 13455 13263 13481
rect 9703 13449 9729 13455
rect 14631 13425 14657 13431
rect 14631 13393 14657 13399
rect 672 13341 20328 13358
rect 672 13315 9919 13341
rect 9945 13315 9971 13341
rect 9997 13315 10023 13341
rect 10049 13315 20328 13341
rect 672 13298 20328 13315
rect 9703 13257 9729 13263
rect 9703 13225 9729 13231
rect 9815 13257 9841 13263
rect 9815 13225 9841 13231
rect 10711 13257 10737 13263
rect 10711 13225 10737 13231
rect 11271 13257 11297 13263
rect 11271 13225 11297 13231
rect 11887 13257 11913 13263
rect 11887 13225 11913 13231
rect 14575 13257 14601 13263
rect 14575 13225 14601 13231
rect 10767 13201 10793 13207
rect 10767 13169 10793 13175
rect 10879 13201 10905 13207
rect 10879 13169 10905 13175
rect 11047 13201 11073 13207
rect 11047 13169 11073 13175
rect 9367 13145 9393 13151
rect 9367 13113 9393 13119
rect 9479 13145 9505 13151
rect 9479 13113 9505 13119
rect 9591 13145 9617 13151
rect 9591 13113 9617 13119
rect 9871 13145 9897 13151
rect 9871 13113 9897 13119
rect 10599 13145 10625 13151
rect 10599 13113 10625 13119
rect 11159 13145 11185 13151
rect 11159 13113 11185 13119
rect 11383 13145 11409 13151
rect 11383 13113 11409 13119
rect 11775 13145 11801 13151
rect 11775 13113 11801 13119
rect 11943 13145 11969 13151
rect 14463 13145 14489 13151
rect 12945 13119 12951 13145
rect 12977 13119 12983 13145
rect 11943 13113 11969 13119
rect 14463 13113 14489 13119
rect 14631 13145 14657 13151
rect 18937 13119 18943 13145
rect 18969 13119 18975 13145
rect 14631 13113 14657 13119
rect 9535 13089 9561 13095
rect 14855 13089 14881 13095
rect 13281 13063 13287 13089
rect 13313 13063 13319 13089
rect 14345 13063 14351 13089
rect 14377 13063 14383 13089
rect 19945 13063 19951 13089
rect 19977 13063 19983 13089
rect 9535 13057 9561 13063
rect 14855 13057 14881 13063
rect 672 12949 20328 12966
rect 672 12923 2239 12949
rect 2265 12923 2291 12949
rect 2317 12923 2343 12949
rect 2369 12923 17599 12949
rect 17625 12923 17651 12949
rect 17677 12923 17703 12949
rect 17729 12923 20328 12949
rect 672 12906 20328 12923
rect 9591 12865 9617 12871
rect 9591 12833 9617 12839
rect 13231 12865 13257 12871
rect 13231 12833 13257 12839
rect 13399 12865 13425 12871
rect 13399 12833 13425 12839
rect 14631 12865 14657 12871
rect 14631 12833 14657 12839
rect 20007 12809 20033 12815
rect 8633 12783 8639 12809
rect 8665 12783 8671 12809
rect 20007 12777 20033 12783
rect 10823 12753 10849 12759
rect 7177 12727 7183 12753
rect 7209 12727 7215 12753
rect 9249 12727 9255 12753
rect 9281 12727 9287 12753
rect 10823 12721 10849 12727
rect 13287 12753 13313 12759
rect 13287 12721 13313 12727
rect 13735 12753 13761 12759
rect 13735 12721 13761 12727
rect 14071 12753 14097 12759
rect 14071 12721 14097 12727
rect 14575 12753 14601 12759
rect 18825 12727 18831 12753
rect 18857 12727 18863 12753
rect 14575 12721 14601 12727
rect 9367 12697 9393 12703
rect 7569 12671 7575 12697
rect 7601 12671 7607 12697
rect 9367 12665 9393 12671
rect 9871 12697 9897 12703
rect 9871 12665 9897 12671
rect 10655 12697 10681 12703
rect 10655 12665 10681 12671
rect 13567 12697 13593 12703
rect 13567 12665 13593 12671
rect 8863 12641 8889 12647
rect 8863 12609 8889 12615
rect 9647 12641 9673 12647
rect 9647 12609 9673 12615
rect 9759 12641 9785 12647
rect 9759 12609 9785 12615
rect 10711 12641 10737 12647
rect 10711 12609 10737 12615
rect 13231 12641 13257 12647
rect 13231 12609 13257 12615
rect 13455 12641 13481 12647
rect 13455 12609 13481 12615
rect 13903 12641 13929 12647
rect 13903 12609 13929 12615
rect 14015 12641 14041 12647
rect 14015 12609 14041 12615
rect 14631 12641 14657 12647
rect 14631 12609 14657 12615
rect 672 12557 20328 12574
rect 672 12531 9919 12557
rect 9945 12531 9971 12557
rect 9997 12531 10023 12557
rect 10049 12531 20328 12557
rect 672 12514 20328 12531
rect 10431 12473 10457 12479
rect 9137 12447 9143 12473
rect 9169 12447 9175 12473
rect 10431 12441 10457 12447
rect 10599 12473 10625 12479
rect 11433 12447 11439 12473
rect 11465 12447 11471 12473
rect 10599 12441 10625 12447
rect 10543 12417 10569 12423
rect 15079 12417 15105 12423
rect 9081 12391 9087 12417
rect 9113 12391 9119 12417
rect 10705 12391 10711 12417
rect 10737 12391 10743 12417
rect 15241 12391 15247 12417
rect 15273 12391 15279 12417
rect 10543 12385 10569 12391
rect 15079 12385 15105 12391
rect 8751 12361 8777 12367
rect 2137 12335 2143 12361
rect 2169 12335 2175 12361
rect 8297 12335 8303 12361
rect 8329 12335 8335 12361
rect 8751 12329 8777 12335
rect 8919 12361 8945 12367
rect 8919 12329 8945 12335
rect 9423 12361 9449 12367
rect 10879 12361 10905 12367
rect 10313 12335 10319 12361
rect 10345 12335 10351 12361
rect 9423 12329 9449 12335
rect 10879 12329 10905 12335
rect 11271 12361 11297 12367
rect 13449 12335 13455 12361
rect 13481 12335 13487 12361
rect 18825 12335 18831 12361
rect 18857 12335 18863 12361
rect 11271 12329 11297 12335
rect 9311 12305 9337 12311
rect 6897 12279 6903 12305
rect 6929 12279 6935 12305
rect 7961 12279 7967 12305
rect 7993 12279 7999 12305
rect 9311 12273 9337 12279
rect 13287 12305 13313 12311
rect 13841 12279 13847 12305
rect 13873 12279 13879 12305
rect 14905 12279 14911 12305
rect 14937 12279 14943 12305
rect 13287 12273 13313 12279
rect 967 12249 993 12255
rect 967 12217 993 12223
rect 9199 12249 9225 12255
rect 9199 12217 9225 12223
rect 20007 12249 20033 12255
rect 20007 12217 20033 12223
rect 672 12165 20328 12182
rect 672 12139 2239 12165
rect 2265 12139 2291 12165
rect 2317 12139 2343 12165
rect 2369 12139 17599 12165
rect 17625 12139 17651 12165
rect 17677 12139 17703 12165
rect 17729 12139 20328 12165
rect 672 12122 20328 12139
rect 8247 12081 8273 12087
rect 8247 12049 8273 12055
rect 8415 12081 8441 12087
rect 8415 12049 8441 12055
rect 13847 12081 13873 12087
rect 13847 12049 13873 12055
rect 967 12025 993 12031
rect 9871 12025 9897 12031
rect 7961 11999 7967 12025
rect 7993 11999 7999 12025
rect 967 11993 993 11999
rect 9871 11993 9897 11999
rect 8695 11969 8721 11975
rect 2137 11943 2143 11969
rect 2169 11943 2175 11969
rect 7905 11943 7911 11969
rect 7937 11943 7943 11969
rect 8695 11937 8721 11943
rect 8919 11969 8945 11975
rect 8919 11937 8945 11943
rect 8975 11969 9001 11975
rect 8975 11937 9001 11943
rect 9087 11969 9113 11975
rect 9087 11937 9113 11943
rect 10039 11969 10065 11975
rect 12161 11943 12167 11969
rect 12193 11943 12199 11969
rect 13897 11943 13903 11969
rect 13929 11943 13935 11969
rect 10039 11937 10065 11943
rect 6791 11913 6817 11919
rect 6791 11881 6817 11887
rect 8079 11913 8105 11919
rect 8079 11881 8105 11887
rect 9199 11913 9225 11919
rect 9199 11881 9225 11887
rect 9927 11913 9953 11919
rect 9927 11881 9953 11887
rect 10263 11913 10289 11919
rect 10263 11881 10289 11887
rect 11999 11913 12025 11919
rect 11999 11881 12025 11887
rect 6735 11857 6761 11863
rect 6735 11825 6761 11831
rect 8303 11857 8329 11863
rect 10151 11857 10177 11863
rect 8913 11831 8919 11857
rect 8945 11831 8951 11857
rect 8303 11825 8329 11831
rect 10151 11825 10177 11831
rect 12055 11857 12081 11863
rect 12055 11825 12081 11831
rect 13679 11857 13705 11863
rect 13679 11825 13705 11831
rect 13791 11857 13817 11863
rect 13791 11825 13817 11831
rect 672 11773 20328 11790
rect 672 11747 9919 11773
rect 9945 11747 9971 11773
rect 9997 11747 10023 11773
rect 10049 11747 20328 11773
rect 672 11730 20328 11747
rect 7575 11689 7601 11695
rect 7575 11657 7601 11663
rect 7687 11689 7713 11695
rect 7687 11657 7713 11663
rect 10263 11689 10289 11695
rect 10263 11657 10289 11663
rect 10543 11689 10569 11695
rect 10543 11657 10569 11663
rect 7631 11633 7657 11639
rect 6729 11607 6735 11633
rect 6761 11607 6767 11633
rect 7631 11601 7657 11607
rect 9591 11633 9617 11639
rect 9591 11601 9617 11607
rect 10207 11633 10233 11639
rect 10207 11601 10233 11607
rect 10431 11633 10457 11639
rect 10431 11601 10457 11607
rect 7519 11577 7545 11583
rect 9927 11577 9953 11583
rect 10375 11577 10401 11583
rect 7121 11551 7127 11577
rect 7153 11551 7159 11577
rect 7401 11551 7407 11577
rect 7433 11551 7439 11577
rect 9137 11551 9143 11577
rect 9169 11551 9175 11577
rect 10089 11551 10095 11577
rect 10121 11551 10127 11577
rect 10929 11551 10935 11577
rect 10961 11551 10967 11577
rect 18825 11551 18831 11577
rect 18857 11551 18863 11577
rect 7519 11545 7545 11551
rect 9927 11545 9953 11551
rect 10375 11545 10401 11551
rect 7967 11521 7993 11527
rect 5665 11495 5671 11521
rect 5697 11495 5703 11521
rect 7967 11489 7993 11495
rect 9367 11521 9393 11527
rect 12671 11521 12697 11527
rect 9529 11495 9535 11521
rect 9561 11495 9567 11521
rect 11265 11495 11271 11521
rect 11297 11495 11303 11521
rect 12329 11495 12335 11521
rect 12361 11495 12367 11521
rect 9367 11489 9393 11495
rect 12671 11489 12697 11495
rect 9703 11465 9729 11471
rect 9703 11433 9729 11439
rect 20007 11465 20033 11471
rect 20007 11433 20033 11439
rect 672 11381 20328 11398
rect 672 11355 2239 11381
rect 2265 11355 2291 11381
rect 2317 11355 2343 11381
rect 2369 11355 17599 11381
rect 17625 11355 17651 11381
rect 17677 11355 17703 11381
rect 17729 11355 20328 11381
rect 672 11338 20328 11355
rect 11663 11297 11689 11303
rect 9081 11271 9087 11297
rect 9113 11271 9119 11297
rect 11663 11265 11689 11271
rect 10039 11241 10065 11247
rect 9193 11215 9199 11241
rect 9225 11215 9231 11241
rect 10039 11209 10065 11215
rect 20007 11241 20033 11247
rect 20007 11209 20033 11215
rect 9815 11185 9841 11191
rect 9305 11159 9311 11185
rect 9337 11159 9343 11185
rect 9473 11159 9479 11185
rect 9505 11159 9511 11185
rect 9815 11153 9841 11159
rect 9927 11185 9953 11191
rect 9927 11153 9953 11159
rect 10095 11185 10121 11191
rect 10095 11153 10121 11159
rect 10207 11185 10233 11191
rect 11887 11185 11913 11191
rect 11545 11159 11551 11185
rect 11577 11159 11583 11185
rect 10207 11153 10233 11159
rect 11887 11153 11913 11159
rect 13959 11185 13985 11191
rect 14519 11185 14545 11191
rect 14121 11159 14127 11185
rect 14153 11159 14159 11185
rect 18825 11159 18831 11185
rect 18857 11159 18863 11185
rect 13959 11153 13985 11159
rect 14519 11153 14545 11159
rect 10655 11129 10681 11135
rect 13847 11129 13873 11135
rect 10375 11101 10401 11107
rect 7239 11073 7265 11079
rect 7239 11041 7265 11047
rect 10319 11073 10345 11079
rect 11769 11103 11775 11129
rect 11801 11103 11807 11129
rect 13113 11103 13119 11129
rect 13145 11103 13151 11129
rect 10655 11097 10681 11103
rect 13847 11097 13873 11103
rect 14687 11129 14713 11135
rect 14687 11097 14713 11103
rect 10375 11069 10401 11075
rect 11495 11073 11521 11079
rect 10817 11047 10823 11073
rect 10849 11047 10855 11073
rect 10319 11041 10345 11047
rect 11495 11041 11521 11047
rect 12951 11073 12977 11079
rect 12951 11041 12977 11047
rect 13903 11073 13929 11079
rect 13903 11041 13929 11047
rect 14631 11073 14657 11079
rect 14631 11041 14657 11047
rect 672 10989 20328 11006
rect 672 10963 9919 10989
rect 9945 10963 9971 10989
rect 9997 10963 10023 10989
rect 10049 10963 20328 10989
rect 672 10946 20328 10963
rect 8359 10905 8385 10911
rect 9143 10905 9169 10911
rect 7457 10879 7463 10905
rect 7489 10879 7495 10905
rect 8913 10879 8919 10905
rect 8945 10879 8951 10905
rect 8359 10873 8385 10879
rect 9143 10873 9169 10879
rect 10991 10905 11017 10911
rect 12727 10905 12753 10911
rect 11209 10879 11215 10905
rect 11241 10879 11247 10905
rect 10991 10873 11017 10879
rect 12727 10873 12753 10879
rect 8415 10849 8441 10855
rect 10879 10849 10905 10855
rect 8129 10823 8135 10849
rect 8161 10823 8167 10849
rect 10313 10823 10319 10849
rect 10345 10823 10351 10849
rect 10425 10823 10431 10849
rect 10457 10823 10463 10849
rect 14009 10823 14015 10849
rect 14041 10823 14047 10849
rect 8415 10817 8441 10823
rect 10879 10817 10905 10823
rect 7295 10793 7321 10799
rect 9087 10793 9113 10799
rect 12615 10793 12641 10799
rect 6449 10767 6455 10793
rect 6481 10767 6487 10793
rect 8017 10767 8023 10793
rect 8049 10767 8055 10793
rect 8801 10767 8807 10793
rect 8833 10767 8839 10793
rect 9641 10767 9647 10793
rect 9673 10767 9679 10793
rect 10033 10767 10039 10793
rect 10065 10767 10071 10793
rect 10201 10767 10207 10793
rect 10233 10767 10239 10793
rect 11321 10767 11327 10793
rect 11353 10767 11359 10793
rect 11657 10767 11663 10793
rect 11689 10767 11695 10793
rect 7295 10761 7321 10767
rect 9087 10761 9113 10767
rect 12615 10761 12641 10767
rect 12951 10793 12977 10799
rect 13617 10767 13623 10793
rect 13649 10767 13655 10793
rect 18937 10767 18943 10793
rect 18969 10767 18975 10793
rect 12951 10761 12977 10767
rect 6679 10737 6705 10743
rect 6505 10711 6511 10737
rect 6537 10711 6543 10737
rect 6679 10705 6705 10711
rect 6903 10737 6929 10743
rect 10767 10737 10793 10743
rect 12055 10737 12081 10743
rect 9697 10711 9703 10737
rect 9729 10711 9735 10737
rect 9921 10711 9927 10737
rect 9953 10711 9959 10737
rect 11041 10711 11047 10737
rect 11073 10711 11079 10737
rect 11825 10711 11831 10737
rect 11857 10711 11863 10737
rect 6903 10705 6929 10711
rect 10767 10705 10793 10711
rect 12055 10705 12081 10711
rect 12671 10737 12697 10743
rect 12671 10705 12697 10711
rect 13455 10737 13481 10743
rect 15073 10711 15079 10737
rect 15105 10711 15111 10737
rect 19945 10711 19951 10737
rect 19977 10711 19983 10737
rect 13455 10705 13481 10711
rect 8359 10681 8385 10687
rect 8359 10649 8385 10655
rect 12111 10681 12137 10687
rect 12111 10649 12137 10655
rect 672 10597 20328 10614
rect 672 10571 2239 10597
rect 2265 10571 2291 10597
rect 2317 10571 2343 10597
rect 2369 10571 17599 10597
rect 17625 10571 17651 10597
rect 17677 10571 17703 10597
rect 17729 10571 20328 10597
rect 672 10554 20328 10571
rect 15079 10513 15105 10519
rect 15079 10481 15105 10487
rect 10879 10457 10905 10463
rect 20007 10457 20033 10463
rect 6449 10431 6455 10457
rect 6481 10431 6487 10457
rect 7737 10431 7743 10457
rect 7769 10431 7775 10457
rect 13449 10431 13455 10457
rect 13481 10431 13487 10457
rect 10879 10425 10905 10431
rect 20007 10425 20033 10431
rect 6791 10401 6817 10407
rect 14575 10401 14601 10407
rect 5049 10375 5055 10401
rect 5081 10375 5087 10401
rect 10033 10375 10039 10401
rect 10065 10375 10071 10401
rect 11265 10375 11271 10401
rect 11297 10375 11303 10401
rect 6791 10369 6817 10375
rect 14575 10369 14601 10375
rect 14911 10401 14937 10407
rect 14911 10369 14937 10375
rect 15023 10401 15049 10407
rect 18825 10375 18831 10401
rect 18857 10375 18863 10401
rect 15023 10369 15049 10375
rect 10711 10345 10737 10351
rect 5385 10319 5391 10345
rect 5417 10319 5423 10345
rect 7289 10319 7295 10345
rect 7321 10319 7327 10345
rect 10711 10313 10737 10319
rect 10935 10345 10961 10351
rect 10935 10313 10961 10319
rect 6959 10289 6985 10295
rect 6959 10257 6985 10263
rect 7463 10289 7489 10295
rect 7463 10257 7489 10263
rect 10823 10289 10849 10295
rect 10823 10257 10849 10263
rect 14631 10289 14657 10295
rect 14631 10257 14657 10263
rect 14687 10289 14713 10295
rect 14687 10257 14713 10263
rect 15079 10289 15105 10295
rect 15079 10257 15105 10263
rect 672 10205 20328 10222
rect 672 10179 9919 10205
rect 9945 10179 9971 10205
rect 9997 10179 10023 10205
rect 10049 10179 20328 10205
rect 672 10162 20328 10179
rect 7351 10121 7377 10127
rect 7351 10089 7377 10095
rect 8471 10121 8497 10127
rect 8471 10089 8497 10095
rect 9255 10121 9281 10127
rect 12945 10095 12951 10121
rect 12977 10095 12983 10121
rect 9255 10089 9281 10095
rect 6785 10039 6791 10065
rect 6817 10039 6823 10065
rect 11265 10039 11271 10065
rect 11297 10039 11303 10065
rect 14009 10039 14015 10065
rect 14041 10039 14047 10065
rect 8303 10009 8329 10015
rect 5049 9983 5055 10009
rect 5081 9983 5087 10009
rect 5385 9983 5391 10009
rect 5417 9983 5423 10009
rect 6673 9983 6679 10009
rect 6705 9983 6711 10009
rect 7065 9983 7071 10009
rect 7097 9983 7103 10009
rect 8073 9983 8079 10009
rect 8105 9983 8111 10009
rect 8303 9977 8329 9983
rect 8807 10009 8833 10015
rect 12671 10009 12697 10015
rect 9417 9983 9423 10009
rect 9449 9983 9455 10009
rect 8807 9977 8833 9983
rect 12671 9977 12697 9983
rect 12727 10009 12753 10015
rect 12727 9977 12753 9983
rect 12839 10009 12865 10015
rect 12839 9977 12865 9983
rect 12951 10009 12977 10015
rect 13617 9983 13623 10009
rect 13649 9983 13655 10009
rect 12951 9977 12977 9983
rect 8975 9953 9001 9959
rect 6449 9927 6455 9953
rect 6481 9927 6487 9953
rect 7177 9927 7183 9953
rect 7209 9927 7215 9953
rect 7569 9927 7575 9953
rect 7601 9927 7607 9953
rect 8241 9927 8247 9953
rect 8273 9927 8279 9953
rect 8975 9921 9001 9927
rect 13455 9953 13481 9959
rect 15073 9927 15079 9953
rect 15105 9927 15111 9953
rect 13455 9921 13481 9927
rect 672 9813 20328 9830
rect 672 9787 2239 9813
rect 2265 9787 2291 9813
rect 2317 9787 2343 9813
rect 2369 9787 17599 9813
rect 17625 9787 17651 9813
rect 17677 9787 17703 9813
rect 17729 9787 20328 9813
rect 672 9770 20328 9787
rect 8415 9673 8441 9679
rect 9529 9647 9535 9673
rect 9561 9647 9567 9673
rect 12217 9647 12223 9673
rect 12249 9647 12255 9673
rect 13281 9647 13287 9673
rect 13313 9647 13319 9673
rect 8415 9641 8441 9647
rect 8135 9617 8161 9623
rect 11663 9617 11689 9623
rect 7289 9591 7295 9617
rect 7321 9591 7327 9617
rect 7401 9591 7407 9617
rect 7433 9591 7439 9617
rect 8913 9591 8919 9617
rect 8945 9591 8951 9617
rect 10369 9591 10375 9617
rect 10401 9591 10407 9617
rect 11825 9591 11831 9617
rect 11857 9591 11863 9617
rect 8135 9585 8161 9591
rect 11663 9585 11689 9591
rect 11439 9561 11465 9567
rect 9193 9535 9199 9561
rect 9225 9535 9231 9561
rect 9585 9535 9591 9561
rect 9617 9535 9623 9561
rect 10929 9535 10935 9561
rect 10961 9535 10967 9561
rect 11439 9529 11465 9535
rect 14239 9561 14265 9567
rect 14239 9529 14265 9535
rect 6791 9505 6817 9511
rect 6791 9473 6817 9479
rect 7519 9505 7545 9511
rect 7519 9473 7545 9479
rect 7575 9505 7601 9511
rect 7575 9473 7601 9479
rect 11103 9505 11129 9511
rect 11103 9473 11129 9479
rect 11551 9505 11577 9511
rect 11551 9473 11577 9479
rect 11607 9505 11633 9511
rect 11607 9473 11633 9479
rect 13511 9505 13537 9511
rect 13511 9473 13537 9479
rect 14071 9505 14097 9511
rect 14071 9473 14097 9479
rect 14183 9505 14209 9511
rect 14183 9473 14209 9479
rect 672 9421 20328 9438
rect 672 9395 9919 9421
rect 9945 9395 9971 9421
rect 9997 9395 10023 9421
rect 10049 9395 20328 9421
rect 672 9378 20328 9395
rect 8751 9337 8777 9343
rect 8751 9305 8777 9311
rect 11719 9281 11745 9287
rect 8913 9255 8919 9281
rect 8945 9255 8951 9281
rect 10537 9255 10543 9281
rect 10569 9255 10575 9281
rect 10985 9255 10991 9281
rect 11017 9255 11023 9281
rect 11719 9249 11745 9255
rect 11831 9281 11857 9287
rect 11831 9249 11857 9255
rect 11943 9281 11969 9287
rect 11943 9249 11969 9255
rect 7127 9225 7153 9231
rect 7127 9193 7153 9199
rect 7239 9225 7265 9231
rect 7239 9193 7265 9199
rect 7463 9225 7489 9231
rect 8415 9225 8441 9231
rect 11999 9225 12025 9231
rect 7681 9199 7687 9225
rect 7713 9199 7719 9225
rect 8969 9199 8975 9225
rect 9001 9199 9007 9225
rect 9305 9199 9311 9225
rect 9337 9199 9343 9225
rect 9529 9199 9535 9225
rect 9561 9199 9567 9225
rect 9809 9199 9815 9225
rect 9841 9199 9847 9225
rect 11097 9199 11103 9225
rect 11129 9199 11135 9225
rect 13393 9199 13399 9225
rect 13425 9199 13431 9225
rect 18825 9199 18831 9225
rect 18857 9199 18863 9225
rect 7463 9193 7489 9199
rect 8415 9193 8441 9199
rect 11999 9193 12025 9199
rect 8695 9169 8721 9175
rect 8185 9143 8191 9169
rect 8217 9143 8223 9169
rect 8695 9137 8721 9143
rect 11887 9169 11913 9175
rect 11887 9137 11913 9143
rect 13231 9169 13257 9175
rect 13785 9143 13791 9169
rect 13817 9143 13823 9169
rect 14849 9143 14855 9169
rect 14881 9143 14887 9169
rect 13231 9137 13257 9143
rect 7407 9113 7433 9119
rect 6953 9087 6959 9113
rect 6985 9087 6991 9113
rect 7407 9081 7433 9087
rect 7575 9113 7601 9119
rect 7575 9081 7601 9087
rect 9703 9113 9729 9119
rect 9703 9081 9729 9087
rect 11383 9113 11409 9119
rect 11383 9081 11409 9087
rect 20007 9113 20033 9119
rect 20007 9081 20033 9087
rect 672 9029 20328 9046
rect 672 9003 2239 9029
rect 2265 9003 2291 9029
rect 2317 9003 2343 9029
rect 2369 9003 17599 9029
rect 17625 9003 17651 9029
rect 17677 9003 17703 9029
rect 17729 9003 20328 9029
rect 672 8986 20328 9003
rect 7183 8945 7209 8951
rect 7183 8913 7209 8919
rect 8527 8945 8553 8951
rect 8527 8913 8553 8919
rect 8975 8945 9001 8951
rect 8975 8913 9001 8919
rect 967 8889 993 8895
rect 9759 8889 9785 8895
rect 13511 8889 13537 8895
rect 4993 8863 4999 8889
rect 5025 8863 5031 8889
rect 11881 8863 11887 8889
rect 11913 8863 11919 8889
rect 12945 8863 12951 8889
rect 12977 8863 12983 8889
rect 967 8857 993 8863
rect 9759 8857 9785 8863
rect 13511 8857 13537 8863
rect 20007 8889 20033 8895
rect 20007 8857 20033 8863
rect 7295 8833 7321 8839
rect 2137 8807 2143 8833
rect 2169 8807 2175 8833
rect 6393 8807 6399 8833
rect 6425 8807 6431 8833
rect 7065 8807 7071 8833
rect 7097 8807 7103 8833
rect 7295 8801 7321 8807
rect 7407 8833 7433 8839
rect 9927 8833 9953 8839
rect 8689 8807 8695 8833
rect 8721 8807 8727 8833
rect 8857 8807 8863 8833
rect 8889 8807 8895 8833
rect 9249 8807 9255 8833
rect 9281 8807 9287 8833
rect 9473 8807 9479 8833
rect 9505 8807 9511 8833
rect 7407 8801 7433 8807
rect 9927 8801 9953 8807
rect 10151 8833 10177 8839
rect 10151 8801 10177 8807
rect 10599 8833 10625 8839
rect 10599 8801 10625 8807
rect 10823 8833 10849 8839
rect 10823 8801 10849 8807
rect 10935 8833 10961 8839
rect 10935 8801 10961 8807
rect 11103 8833 11129 8839
rect 13343 8833 13369 8839
rect 11545 8807 11551 8833
rect 11577 8807 11583 8833
rect 11103 8801 11129 8807
rect 13343 8801 13369 8807
rect 13455 8833 13481 8839
rect 13455 8801 13481 8807
rect 13623 8833 13649 8839
rect 13623 8801 13649 8807
rect 13735 8833 13761 8839
rect 13735 8801 13761 8807
rect 13903 8833 13929 8839
rect 13903 8801 13929 8807
rect 14071 8833 14097 8839
rect 14071 8801 14097 8807
rect 14295 8833 14321 8839
rect 18825 8807 18831 8833
rect 18857 8807 18863 8833
rect 14295 8801 14321 8807
rect 8583 8777 8609 8783
rect 10319 8777 10345 8783
rect 14127 8777 14153 8783
rect 6057 8751 6063 8777
rect 6089 8751 6095 8777
rect 8913 8751 8919 8777
rect 8945 8751 8951 8777
rect 11265 8751 11271 8777
rect 11297 8751 11303 8777
rect 8583 8745 8609 8751
rect 10319 8745 10345 8751
rect 14127 8745 14153 8751
rect 14239 8777 14265 8783
rect 14239 8745 14265 8751
rect 6791 8721 6817 8727
rect 6791 8689 6817 8695
rect 7127 8721 7153 8727
rect 7127 8689 7153 8695
rect 10375 8721 10401 8727
rect 10375 8689 10401 8695
rect 10767 8721 10793 8727
rect 10767 8689 10793 8695
rect 13903 8721 13929 8727
rect 13903 8689 13929 8695
rect 672 8637 20328 8654
rect 672 8611 9919 8637
rect 9945 8611 9971 8637
rect 9997 8611 10023 8637
rect 10049 8611 20328 8637
rect 672 8594 20328 8611
rect 5895 8553 5921 8559
rect 5895 8521 5921 8527
rect 6959 8553 6985 8559
rect 6959 8521 6985 8527
rect 7015 8553 7041 8559
rect 7015 8521 7041 8527
rect 7855 8553 7881 8559
rect 7855 8521 7881 8527
rect 8751 8553 8777 8559
rect 8751 8521 8777 8527
rect 9759 8553 9785 8559
rect 9759 8521 9785 8527
rect 10375 8553 10401 8559
rect 10375 8521 10401 8527
rect 10543 8553 10569 8559
rect 10705 8527 10711 8553
rect 10737 8527 10743 8553
rect 10873 8527 10879 8553
rect 10905 8527 10911 8553
rect 10543 8521 10569 8527
rect 7911 8497 7937 8503
rect 7569 8471 7575 8497
rect 7601 8471 7607 8497
rect 7911 8465 7937 8471
rect 8695 8497 8721 8503
rect 8695 8465 8721 8471
rect 11383 8497 11409 8503
rect 11545 8471 11551 8497
rect 11577 8471 11583 8497
rect 13841 8471 13847 8497
rect 13873 8471 13879 8497
rect 11383 8465 11409 8471
rect 7071 8441 7097 8447
rect 2137 8415 2143 8441
rect 2169 8415 2175 8441
rect 5777 8415 5783 8441
rect 5809 8415 5815 8441
rect 7071 8409 7097 8415
rect 7295 8441 7321 8447
rect 7743 8441 7769 8447
rect 9591 8441 9617 8447
rect 7457 8415 7463 8441
rect 7489 8415 7495 8441
rect 9193 8415 9199 8441
rect 9225 8415 9231 8441
rect 7295 8409 7321 8415
rect 7743 8409 7769 8415
rect 9591 8409 9617 8415
rect 10095 8441 10121 8447
rect 13063 8441 13089 8447
rect 10985 8415 10991 8441
rect 11017 8415 11023 8441
rect 10095 8409 10121 8415
rect 13063 8409 13089 8415
rect 13287 8441 13313 8447
rect 13449 8415 13455 8441
rect 13481 8415 13487 8441
rect 18937 8415 18943 8441
rect 18969 8415 18975 8441
rect 13287 8409 13313 8415
rect 9535 8385 9561 8391
rect 20007 8385 20033 8391
rect 9025 8359 9031 8385
rect 9057 8359 9063 8385
rect 14905 8359 14911 8385
rect 14937 8359 14943 8385
rect 9535 8353 9561 8359
rect 20007 8353 20033 8359
rect 967 8329 993 8335
rect 967 8297 993 8303
rect 8751 8329 8777 8335
rect 8751 8297 8777 8303
rect 672 8245 20328 8262
rect 672 8219 2239 8245
rect 2265 8219 2291 8245
rect 2317 8219 2343 8245
rect 2369 8219 17599 8245
rect 17625 8219 17651 8245
rect 17677 8219 17703 8245
rect 17729 8219 20328 8245
rect 672 8202 20328 8219
rect 6791 8161 6817 8167
rect 6791 8129 6817 8135
rect 9983 8105 10009 8111
rect 9983 8073 10009 8079
rect 6959 8049 6985 8055
rect 6959 8017 6985 8023
rect 7239 8049 7265 8055
rect 7239 8017 7265 8023
rect 7743 8049 7769 8055
rect 10599 8049 10625 8055
rect 12503 8049 12529 8055
rect 10201 8023 10207 8049
rect 10233 8023 10239 8049
rect 10761 8023 10767 8049
rect 10793 8023 10799 8049
rect 7743 8017 7769 8023
rect 10599 8017 10625 8023
rect 12503 8017 12529 8023
rect 7183 7993 7209 7999
rect 6847 7965 6873 7971
rect 6791 7937 6817 7943
rect 7183 7961 7209 7967
rect 7687 7993 7713 7999
rect 7687 7961 7713 7967
rect 6847 7933 6873 7939
rect 7071 7937 7097 7943
rect 6791 7905 6817 7911
rect 7071 7905 7097 7911
rect 7575 7937 7601 7943
rect 7575 7905 7601 7911
rect 10879 7937 10905 7943
rect 10879 7905 10905 7911
rect 10935 7937 10961 7943
rect 10935 7905 10961 7911
rect 12335 7937 12361 7943
rect 12335 7905 12361 7911
rect 12447 7937 12473 7943
rect 12447 7905 12473 7911
rect 672 7853 20328 7870
rect 672 7827 9919 7853
rect 9945 7827 9971 7853
rect 9997 7827 10023 7853
rect 10049 7827 20328 7853
rect 672 7810 20328 7827
rect 8751 7713 8777 7719
rect 6393 7687 6399 7713
rect 6425 7687 6431 7713
rect 7345 7687 7351 7713
rect 7377 7687 7383 7713
rect 8751 7681 8777 7687
rect 8807 7713 8833 7719
rect 8807 7681 8833 7687
rect 12111 7713 12137 7719
rect 12111 7681 12137 7687
rect 8639 7657 8665 7663
rect 6785 7631 6791 7657
rect 6817 7631 6823 7657
rect 7009 7631 7015 7657
rect 7041 7631 7047 7657
rect 8639 7625 8665 7631
rect 10095 7657 10121 7663
rect 10655 7657 10681 7663
rect 10313 7631 10319 7657
rect 10345 7631 10351 7657
rect 10095 7625 10121 7631
rect 10655 7625 10681 7631
rect 10711 7657 10737 7663
rect 10711 7625 10737 7631
rect 10823 7657 10849 7663
rect 11887 7657 11913 7663
rect 10929 7631 10935 7657
rect 10961 7631 10967 7657
rect 10823 7625 10849 7631
rect 11887 7625 11913 7631
rect 11999 7657 12025 7663
rect 11999 7625 12025 7631
rect 12167 7657 12193 7663
rect 12167 7625 12193 7631
rect 9031 7601 9057 7607
rect 5329 7575 5335 7601
rect 5361 7575 5367 7601
rect 8409 7575 8415 7601
rect 8441 7575 8447 7601
rect 9031 7569 9057 7575
rect 10207 7601 10233 7607
rect 10873 7575 10879 7601
rect 10905 7575 10911 7601
rect 10207 7569 10233 7575
rect 10039 7545 10065 7551
rect 10039 7513 10065 7519
rect 672 7461 20328 7478
rect 672 7435 2239 7461
rect 2265 7435 2291 7461
rect 2317 7435 2343 7461
rect 2369 7435 17599 7461
rect 17625 7435 17651 7461
rect 17677 7435 17703 7461
rect 17729 7435 20328 7461
rect 672 7418 20328 7435
rect 9871 7377 9897 7383
rect 9871 7345 9897 7351
rect 6903 7321 6929 7327
rect 9815 7321 9841 7327
rect 8577 7295 8583 7321
rect 8609 7295 8615 7321
rect 9641 7295 9647 7321
rect 9673 7295 9679 7321
rect 6903 7289 6929 7295
rect 9815 7289 9841 7295
rect 10095 7321 10121 7327
rect 12049 7295 12055 7321
rect 12081 7295 12087 7321
rect 13113 7295 13119 7321
rect 13145 7295 13151 7321
rect 10095 7289 10121 7295
rect 8241 7239 8247 7265
rect 8273 7239 8279 7265
rect 11657 7239 11663 7265
rect 11689 7239 11695 7265
rect 10711 7209 10737 7215
rect 10711 7177 10737 7183
rect 10767 7209 10793 7215
rect 10767 7177 10793 7183
rect 10599 7153 10625 7159
rect 10599 7121 10625 7127
rect 13343 7153 13369 7159
rect 13343 7121 13369 7127
rect 672 7069 20328 7086
rect 672 7043 9919 7069
rect 9945 7043 9971 7069
rect 9997 7043 10023 7069
rect 10049 7043 20328 7069
rect 672 7026 20328 7043
rect 12223 6985 12249 6991
rect 12223 6953 12249 6959
rect 12895 6985 12921 6991
rect 12895 6953 12921 6959
rect 8359 6929 8385 6935
rect 8359 6897 8385 6903
rect 8415 6929 8441 6935
rect 12615 6929 12641 6935
rect 10089 6903 10095 6929
rect 10121 6903 10127 6929
rect 8415 6897 8441 6903
rect 12615 6897 12641 6903
rect 12671 6929 12697 6935
rect 13057 6903 13063 6929
rect 13089 6903 13095 6929
rect 12671 6897 12697 6903
rect 8247 6873 8273 6879
rect 11999 6873 12025 6879
rect 9753 6847 9759 6873
rect 9785 6847 9791 6873
rect 8247 6841 8273 6847
rect 11999 6841 12025 6847
rect 12279 6873 12305 6879
rect 12279 6841 12305 6847
rect 12783 6873 12809 6879
rect 12783 6841 12809 6847
rect 11383 6817 11409 6823
rect 11153 6791 11159 6817
rect 11185 6791 11191 6817
rect 11383 6785 11409 6791
rect 12223 6761 12249 6767
rect 12223 6729 12249 6735
rect 672 6677 20328 6694
rect 672 6651 2239 6677
rect 2265 6651 2291 6677
rect 2317 6651 2343 6677
rect 2369 6651 17599 6677
rect 17625 6651 17651 6677
rect 17677 6651 17703 6677
rect 17729 6651 20328 6677
rect 672 6634 20328 6651
rect 8919 6593 8945 6599
rect 8919 6561 8945 6567
rect 10767 6593 10793 6599
rect 10767 6561 10793 6567
rect 9199 6537 9225 6543
rect 7625 6511 7631 6537
rect 7657 6511 7663 6537
rect 8689 6511 8695 6537
rect 8721 6511 8727 6537
rect 9199 6505 9225 6511
rect 11047 6537 11073 6543
rect 13511 6537 13537 6543
rect 12217 6511 12223 6537
rect 12249 6511 12255 6537
rect 13281 6511 13287 6537
rect 13313 6511 13319 6537
rect 11047 6505 11073 6511
rect 13511 6505 13537 6511
rect 8975 6481 9001 6487
rect 7289 6455 7295 6481
rect 7321 6455 7327 6481
rect 8975 6449 9001 6455
rect 10823 6481 10849 6487
rect 11825 6455 11831 6481
rect 11857 6455 11863 6481
rect 10823 6449 10849 6455
rect 8919 6369 8945 6375
rect 8919 6337 8945 6343
rect 10767 6369 10793 6375
rect 10767 6337 10793 6343
rect 672 6285 20328 6302
rect 672 6259 9919 6285
rect 9945 6259 9971 6285
rect 9997 6259 10023 6285
rect 10049 6259 20328 6285
rect 672 6242 20328 6259
rect 8863 6201 8889 6207
rect 8863 6169 8889 6175
rect 11439 6201 11465 6207
rect 11439 6169 11465 6175
rect 10145 6119 10151 6145
rect 10177 6119 10183 6145
rect 9753 6063 9759 6089
rect 9785 6063 9791 6089
rect 11209 6007 11215 6033
rect 11241 6007 11247 6033
rect 672 5893 20328 5910
rect 672 5867 2239 5893
rect 2265 5867 2291 5893
rect 2317 5867 2343 5893
rect 2369 5867 17599 5893
rect 17625 5867 17651 5893
rect 17677 5867 17703 5893
rect 17729 5867 20328 5893
rect 672 5850 20328 5867
rect 672 5501 20328 5518
rect 672 5475 9919 5501
rect 9945 5475 9971 5501
rect 9997 5475 10023 5501
rect 10049 5475 20328 5501
rect 672 5458 20328 5475
rect 672 5109 20328 5126
rect 672 5083 2239 5109
rect 2265 5083 2291 5109
rect 2317 5083 2343 5109
rect 2369 5083 17599 5109
rect 17625 5083 17651 5109
rect 17677 5083 17703 5109
rect 17729 5083 20328 5109
rect 672 5066 20328 5083
rect 672 4717 20328 4734
rect 672 4691 9919 4717
rect 9945 4691 9971 4717
rect 9997 4691 10023 4717
rect 10049 4691 20328 4717
rect 672 4674 20328 4691
rect 672 4325 20328 4342
rect 672 4299 2239 4325
rect 2265 4299 2291 4325
rect 2317 4299 2343 4325
rect 2369 4299 17599 4325
rect 17625 4299 17651 4325
rect 17677 4299 17703 4325
rect 17729 4299 20328 4325
rect 672 4282 20328 4299
rect 672 3933 20328 3950
rect 672 3907 9919 3933
rect 9945 3907 9971 3933
rect 9997 3907 10023 3933
rect 10049 3907 20328 3933
rect 672 3890 20328 3907
rect 672 3541 20328 3558
rect 672 3515 2239 3541
rect 2265 3515 2291 3541
rect 2317 3515 2343 3541
rect 2369 3515 17599 3541
rect 17625 3515 17651 3541
rect 17677 3515 17703 3541
rect 17729 3515 20328 3541
rect 672 3498 20328 3515
rect 672 3149 20328 3166
rect 672 3123 9919 3149
rect 9945 3123 9971 3149
rect 9997 3123 10023 3149
rect 10049 3123 20328 3149
rect 672 3106 20328 3123
rect 672 2757 20328 2774
rect 672 2731 2239 2757
rect 2265 2731 2291 2757
rect 2317 2731 2343 2757
rect 2369 2731 17599 2757
rect 17625 2731 17651 2757
rect 17677 2731 17703 2757
rect 17729 2731 20328 2757
rect 672 2714 20328 2731
rect 672 2365 20328 2382
rect 672 2339 9919 2365
rect 9945 2339 9971 2365
rect 9997 2339 10023 2365
rect 10049 2339 20328 2365
rect 672 2322 20328 2339
rect 10929 2143 10935 2169
rect 10961 2143 10967 2169
rect 12889 2143 12895 2169
rect 12921 2143 12927 2169
rect 11383 2057 11409 2063
rect 11383 2025 11409 2031
rect 13399 2057 13425 2063
rect 13399 2025 13425 2031
rect 672 1973 20328 1990
rect 672 1947 2239 1973
rect 2265 1947 2291 1973
rect 2317 1947 2343 1973
rect 2369 1947 17599 1973
rect 17625 1947 17651 1973
rect 17677 1947 17703 1973
rect 17729 1947 20328 1973
rect 672 1930 20328 1947
rect 13063 1833 13089 1839
rect 13063 1801 13089 1807
rect 14687 1833 14713 1839
rect 14687 1801 14713 1807
rect 8521 1751 8527 1777
rect 8553 1751 8559 1777
rect 10705 1751 10711 1777
rect 10737 1751 10743 1777
rect 12609 1751 12615 1777
rect 12641 1751 12647 1777
rect 14289 1751 14295 1777
rect 14321 1751 14327 1777
rect 9031 1665 9057 1671
rect 9031 1633 9057 1639
rect 11215 1665 11241 1671
rect 11215 1633 11241 1639
rect 672 1581 20328 1598
rect 672 1555 9919 1581
rect 9945 1555 9971 1581
rect 9997 1555 10023 1581
rect 10049 1555 20328 1581
rect 672 1538 20328 1555
<< via1 >>
rect 2239 19195 2265 19221
rect 2291 19195 2317 19221
rect 2343 19195 2369 19221
rect 17599 19195 17625 19221
rect 17651 19195 17677 19221
rect 17703 19195 17729 19221
rect 9311 19111 9337 19137
rect 10879 19111 10905 19137
rect 12783 19111 12809 19137
rect 8807 18999 8833 19025
rect 10375 18999 10401 19025
rect 12279 18999 12305 19025
rect 9919 18803 9945 18829
rect 9971 18803 9997 18829
rect 10023 18803 10049 18829
rect 10039 18719 10065 18745
rect 13119 18719 13145 18745
rect 9535 18607 9561 18633
rect 12615 18607 12641 18633
rect 2239 18411 2265 18437
rect 2291 18411 2317 18437
rect 2343 18411 2369 18437
rect 17599 18411 17625 18437
rect 17651 18411 17677 18437
rect 17703 18411 17729 18437
rect 9919 18019 9945 18045
rect 9971 18019 9997 18045
rect 10023 18019 10049 18045
rect 2239 17627 2265 17653
rect 2291 17627 2317 17653
rect 2343 17627 2369 17653
rect 17599 17627 17625 17653
rect 17651 17627 17677 17653
rect 17703 17627 17729 17653
rect 9919 17235 9945 17261
rect 9971 17235 9997 17261
rect 10023 17235 10049 17261
rect 2239 16843 2265 16869
rect 2291 16843 2317 16869
rect 2343 16843 2369 16869
rect 17599 16843 17625 16869
rect 17651 16843 17677 16869
rect 17703 16843 17729 16869
rect 9919 16451 9945 16477
rect 9971 16451 9997 16477
rect 10023 16451 10049 16477
rect 2239 16059 2265 16085
rect 2291 16059 2317 16085
rect 2343 16059 2369 16085
rect 17599 16059 17625 16085
rect 17651 16059 17677 16085
rect 17703 16059 17729 16085
rect 9919 15667 9945 15693
rect 9971 15667 9997 15693
rect 10023 15667 10049 15693
rect 2239 15275 2265 15301
rect 2291 15275 2317 15301
rect 2343 15275 2369 15301
rect 17599 15275 17625 15301
rect 17651 15275 17677 15301
rect 17703 15275 17729 15301
rect 9919 14883 9945 14909
rect 9971 14883 9997 14909
rect 10023 14883 10049 14909
rect 2239 14491 2265 14517
rect 2291 14491 2317 14517
rect 2343 14491 2369 14517
rect 17599 14491 17625 14517
rect 17651 14491 17677 14517
rect 17703 14491 17729 14517
rect 10151 14239 10177 14265
rect 10207 14239 10233 14265
rect 10879 14239 10905 14265
rect 10935 14239 10961 14265
rect 10039 14183 10065 14209
rect 11047 14183 11073 14209
rect 9919 14099 9945 14125
rect 9971 14099 9997 14125
rect 10023 14099 10049 14125
rect 8807 13903 8833 13929
rect 10431 13903 10457 13929
rect 8471 13847 8497 13873
rect 9143 13847 9169 13873
rect 10207 13847 10233 13873
rect 10767 13847 10793 13873
rect 11831 13847 11857 13873
rect 12111 13847 12137 13873
rect 2239 13707 2265 13733
rect 2291 13707 2317 13733
rect 2343 13707 2369 13733
rect 17599 13707 17625 13733
rect 17651 13707 17677 13733
rect 17703 13707 17729 13733
rect 9479 13567 9505 13593
rect 9927 13567 9953 13593
rect 12335 13567 12361 13593
rect 14295 13567 14321 13593
rect 20007 13567 20033 13593
rect 8079 13511 8105 13537
rect 9815 13511 9841 13537
rect 10039 13511 10065 13537
rect 10095 13511 10121 13537
rect 10935 13511 10961 13537
rect 12559 13511 12585 13537
rect 12895 13511 12921 13537
rect 18831 13511 18857 13537
rect 8415 13455 8441 13481
rect 9703 13455 9729 13481
rect 11271 13455 11297 13481
rect 13231 13455 13257 13481
rect 14631 13399 14657 13425
rect 9919 13315 9945 13341
rect 9971 13315 9997 13341
rect 10023 13315 10049 13341
rect 9703 13231 9729 13257
rect 9815 13231 9841 13257
rect 10711 13231 10737 13257
rect 11271 13231 11297 13257
rect 11887 13231 11913 13257
rect 14575 13231 14601 13257
rect 10767 13175 10793 13201
rect 10879 13175 10905 13201
rect 11047 13175 11073 13201
rect 9367 13119 9393 13145
rect 9479 13119 9505 13145
rect 9591 13119 9617 13145
rect 9871 13119 9897 13145
rect 10599 13119 10625 13145
rect 11159 13119 11185 13145
rect 11383 13119 11409 13145
rect 11775 13119 11801 13145
rect 11943 13119 11969 13145
rect 12951 13119 12977 13145
rect 14463 13119 14489 13145
rect 14631 13119 14657 13145
rect 18943 13119 18969 13145
rect 9535 13063 9561 13089
rect 13287 13063 13313 13089
rect 14351 13063 14377 13089
rect 14855 13063 14881 13089
rect 19951 13063 19977 13089
rect 2239 12923 2265 12949
rect 2291 12923 2317 12949
rect 2343 12923 2369 12949
rect 17599 12923 17625 12949
rect 17651 12923 17677 12949
rect 17703 12923 17729 12949
rect 9591 12839 9617 12865
rect 13231 12839 13257 12865
rect 13399 12839 13425 12865
rect 14631 12839 14657 12865
rect 8639 12783 8665 12809
rect 20007 12783 20033 12809
rect 7183 12727 7209 12753
rect 9255 12727 9281 12753
rect 10823 12727 10849 12753
rect 13287 12727 13313 12753
rect 13735 12727 13761 12753
rect 14071 12727 14097 12753
rect 14575 12727 14601 12753
rect 18831 12727 18857 12753
rect 7575 12671 7601 12697
rect 9367 12671 9393 12697
rect 9871 12671 9897 12697
rect 10655 12671 10681 12697
rect 13567 12671 13593 12697
rect 8863 12615 8889 12641
rect 9647 12615 9673 12641
rect 9759 12615 9785 12641
rect 10711 12615 10737 12641
rect 13231 12615 13257 12641
rect 13455 12615 13481 12641
rect 13903 12615 13929 12641
rect 14015 12615 14041 12641
rect 14631 12615 14657 12641
rect 9919 12531 9945 12557
rect 9971 12531 9997 12557
rect 10023 12531 10049 12557
rect 9143 12447 9169 12473
rect 10431 12447 10457 12473
rect 10599 12447 10625 12473
rect 11439 12447 11465 12473
rect 9087 12391 9113 12417
rect 10543 12391 10569 12417
rect 10711 12391 10737 12417
rect 15079 12391 15105 12417
rect 15247 12391 15273 12417
rect 2143 12335 2169 12361
rect 8303 12335 8329 12361
rect 8751 12335 8777 12361
rect 8919 12335 8945 12361
rect 9423 12335 9449 12361
rect 10319 12335 10345 12361
rect 10879 12335 10905 12361
rect 11271 12335 11297 12361
rect 13455 12335 13481 12361
rect 18831 12335 18857 12361
rect 6903 12279 6929 12305
rect 7967 12279 7993 12305
rect 9311 12279 9337 12305
rect 13287 12279 13313 12305
rect 13847 12279 13873 12305
rect 14911 12279 14937 12305
rect 967 12223 993 12249
rect 9199 12223 9225 12249
rect 20007 12223 20033 12249
rect 2239 12139 2265 12165
rect 2291 12139 2317 12165
rect 2343 12139 2369 12165
rect 17599 12139 17625 12165
rect 17651 12139 17677 12165
rect 17703 12139 17729 12165
rect 8247 12055 8273 12081
rect 8415 12055 8441 12081
rect 13847 12055 13873 12081
rect 967 11999 993 12025
rect 7967 11999 7993 12025
rect 9871 11999 9897 12025
rect 2143 11943 2169 11969
rect 7911 11943 7937 11969
rect 8695 11943 8721 11969
rect 8919 11943 8945 11969
rect 8975 11943 9001 11969
rect 9087 11943 9113 11969
rect 10039 11943 10065 11969
rect 12167 11943 12193 11969
rect 13903 11943 13929 11969
rect 6791 11887 6817 11913
rect 8079 11887 8105 11913
rect 9199 11887 9225 11913
rect 9927 11887 9953 11913
rect 10263 11887 10289 11913
rect 11999 11887 12025 11913
rect 6735 11831 6761 11857
rect 8303 11831 8329 11857
rect 8919 11831 8945 11857
rect 10151 11831 10177 11857
rect 12055 11831 12081 11857
rect 13679 11831 13705 11857
rect 13791 11831 13817 11857
rect 9919 11747 9945 11773
rect 9971 11747 9997 11773
rect 10023 11747 10049 11773
rect 7575 11663 7601 11689
rect 7687 11663 7713 11689
rect 10263 11663 10289 11689
rect 10543 11663 10569 11689
rect 6735 11607 6761 11633
rect 7631 11607 7657 11633
rect 9591 11607 9617 11633
rect 10207 11607 10233 11633
rect 10431 11607 10457 11633
rect 7127 11551 7153 11577
rect 7407 11551 7433 11577
rect 7519 11551 7545 11577
rect 9143 11551 9169 11577
rect 9927 11551 9953 11577
rect 10095 11551 10121 11577
rect 10375 11551 10401 11577
rect 10935 11551 10961 11577
rect 18831 11551 18857 11577
rect 5671 11495 5697 11521
rect 7967 11495 7993 11521
rect 9367 11495 9393 11521
rect 9535 11495 9561 11521
rect 11271 11495 11297 11521
rect 12335 11495 12361 11521
rect 12671 11495 12697 11521
rect 9703 11439 9729 11465
rect 20007 11439 20033 11465
rect 2239 11355 2265 11381
rect 2291 11355 2317 11381
rect 2343 11355 2369 11381
rect 17599 11355 17625 11381
rect 17651 11355 17677 11381
rect 17703 11355 17729 11381
rect 9087 11271 9113 11297
rect 11663 11271 11689 11297
rect 9199 11215 9225 11241
rect 10039 11215 10065 11241
rect 20007 11215 20033 11241
rect 9311 11159 9337 11185
rect 9479 11159 9505 11185
rect 9815 11159 9841 11185
rect 9927 11159 9953 11185
rect 10095 11159 10121 11185
rect 10207 11159 10233 11185
rect 11551 11159 11577 11185
rect 11887 11159 11913 11185
rect 13959 11159 13985 11185
rect 14127 11159 14153 11185
rect 14519 11159 14545 11185
rect 18831 11159 18857 11185
rect 7239 11047 7265 11073
rect 10319 11047 10345 11073
rect 10375 11075 10401 11101
rect 10655 11103 10681 11129
rect 11775 11103 11801 11129
rect 13119 11103 13145 11129
rect 13847 11103 13873 11129
rect 14687 11103 14713 11129
rect 10823 11047 10849 11073
rect 11495 11047 11521 11073
rect 12951 11047 12977 11073
rect 13903 11047 13929 11073
rect 14631 11047 14657 11073
rect 9919 10963 9945 10989
rect 9971 10963 9997 10989
rect 10023 10963 10049 10989
rect 7463 10879 7489 10905
rect 8359 10879 8385 10905
rect 8919 10879 8945 10905
rect 9143 10879 9169 10905
rect 10991 10879 11017 10905
rect 11215 10879 11241 10905
rect 12727 10879 12753 10905
rect 8135 10823 8161 10849
rect 8415 10823 8441 10849
rect 10319 10823 10345 10849
rect 10431 10823 10457 10849
rect 10879 10823 10905 10849
rect 14015 10823 14041 10849
rect 6455 10767 6481 10793
rect 7295 10767 7321 10793
rect 8023 10767 8049 10793
rect 8807 10767 8833 10793
rect 9087 10767 9113 10793
rect 9647 10767 9673 10793
rect 10039 10767 10065 10793
rect 10207 10767 10233 10793
rect 11327 10767 11353 10793
rect 11663 10767 11689 10793
rect 12615 10767 12641 10793
rect 12951 10767 12977 10793
rect 13623 10767 13649 10793
rect 18943 10767 18969 10793
rect 6511 10711 6537 10737
rect 6679 10711 6705 10737
rect 6903 10711 6929 10737
rect 9703 10711 9729 10737
rect 9927 10711 9953 10737
rect 10767 10711 10793 10737
rect 11047 10711 11073 10737
rect 11831 10711 11857 10737
rect 12055 10711 12081 10737
rect 12671 10711 12697 10737
rect 13455 10711 13481 10737
rect 15079 10711 15105 10737
rect 19951 10711 19977 10737
rect 8359 10655 8385 10681
rect 12111 10655 12137 10681
rect 2239 10571 2265 10597
rect 2291 10571 2317 10597
rect 2343 10571 2369 10597
rect 17599 10571 17625 10597
rect 17651 10571 17677 10597
rect 17703 10571 17729 10597
rect 15079 10487 15105 10513
rect 6455 10431 6481 10457
rect 7743 10431 7769 10457
rect 10879 10431 10905 10457
rect 13455 10431 13481 10457
rect 20007 10431 20033 10457
rect 5055 10375 5081 10401
rect 6791 10375 6817 10401
rect 10039 10375 10065 10401
rect 11271 10375 11297 10401
rect 14575 10375 14601 10401
rect 14911 10375 14937 10401
rect 15023 10375 15049 10401
rect 18831 10375 18857 10401
rect 5391 10319 5417 10345
rect 7295 10319 7321 10345
rect 10711 10319 10737 10345
rect 10935 10319 10961 10345
rect 6959 10263 6985 10289
rect 7463 10263 7489 10289
rect 10823 10263 10849 10289
rect 14631 10263 14657 10289
rect 14687 10263 14713 10289
rect 15079 10263 15105 10289
rect 9919 10179 9945 10205
rect 9971 10179 9997 10205
rect 10023 10179 10049 10205
rect 7351 10095 7377 10121
rect 8471 10095 8497 10121
rect 9255 10095 9281 10121
rect 12951 10095 12977 10121
rect 6791 10039 6817 10065
rect 11271 10039 11297 10065
rect 14015 10039 14041 10065
rect 5055 9983 5081 10009
rect 5391 9983 5417 10009
rect 6679 9983 6705 10009
rect 7071 9983 7097 10009
rect 8079 9983 8105 10009
rect 8303 9983 8329 10009
rect 8807 9983 8833 10009
rect 9423 9983 9449 10009
rect 12671 9983 12697 10009
rect 12727 9983 12753 10009
rect 12839 9983 12865 10009
rect 12951 9983 12977 10009
rect 13623 9983 13649 10009
rect 6455 9927 6481 9953
rect 7183 9927 7209 9953
rect 7575 9927 7601 9953
rect 8247 9927 8273 9953
rect 8975 9927 9001 9953
rect 13455 9927 13481 9953
rect 15079 9927 15105 9953
rect 2239 9787 2265 9813
rect 2291 9787 2317 9813
rect 2343 9787 2369 9813
rect 17599 9787 17625 9813
rect 17651 9787 17677 9813
rect 17703 9787 17729 9813
rect 8415 9647 8441 9673
rect 9535 9647 9561 9673
rect 12223 9647 12249 9673
rect 13287 9647 13313 9673
rect 7295 9591 7321 9617
rect 7407 9591 7433 9617
rect 8135 9591 8161 9617
rect 8919 9591 8945 9617
rect 10375 9591 10401 9617
rect 11663 9591 11689 9617
rect 11831 9591 11857 9617
rect 9199 9535 9225 9561
rect 9591 9535 9617 9561
rect 10935 9535 10961 9561
rect 11439 9535 11465 9561
rect 14239 9535 14265 9561
rect 6791 9479 6817 9505
rect 7519 9479 7545 9505
rect 7575 9479 7601 9505
rect 11103 9479 11129 9505
rect 11551 9479 11577 9505
rect 11607 9479 11633 9505
rect 13511 9479 13537 9505
rect 14071 9479 14097 9505
rect 14183 9479 14209 9505
rect 9919 9395 9945 9421
rect 9971 9395 9997 9421
rect 10023 9395 10049 9421
rect 8751 9311 8777 9337
rect 8919 9255 8945 9281
rect 10543 9255 10569 9281
rect 10991 9255 11017 9281
rect 11719 9255 11745 9281
rect 11831 9255 11857 9281
rect 11943 9255 11969 9281
rect 7127 9199 7153 9225
rect 7239 9199 7265 9225
rect 7463 9199 7489 9225
rect 7687 9199 7713 9225
rect 8415 9199 8441 9225
rect 8975 9199 9001 9225
rect 9311 9199 9337 9225
rect 9535 9199 9561 9225
rect 9815 9199 9841 9225
rect 11103 9199 11129 9225
rect 11999 9199 12025 9225
rect 13399 9199 13425 9225
rect 18831 9199 18857 9225
rect 8191 9143 8217 9169
rect 8695 9143 8721 9169
rect 11887 9143 11913 9169
rect 13231 9143 13257 9169
rect 13791 9143 13817 9169
rect 14855 9143 14881 9169
rect 6959 9087 6985 9113
rect 7407 9087 7433 9113
rect 7575 9087 7601 9113
rect 9703 9087 9729 9113
rect 11383 9087 11409 9113
rect 20007 9087 20033 9113
rect 2239 9003 2265 9029
rect 2291 9003 2317 9029
rect 2343 9003 2369 9029
rect 17599 9003 17625 9029
rect 17651 9003 17677 9029
rect 17703 9003 17729 9029
rect 7183 8919 7209 8945
rect 8527 8919 8553 8945
rect 8975 8919 9001 8945
rect 967 8863 993 8889
rect 4999 8863 5025 8889
rect 9759 8863 9785 8889
rect 11887 8863 11913 8889
rect 12951 8863 12977 8889
rect 13511 8863 13537 8889
rect 20007 8863 20033 8889
rect 2143 8807 2169 8833
rect 6399 8807 6425 8833
rect 7071 8807 7097 8833
rect 7295 8807 7321 8833
rect 7407 8807 7433 8833
rect 8695 8807 8721 8833
rect 8863 8807 8889 8833
rect 9255 8807 9281 8833
rect 9479 8807 9505 8833
rect 9927 8807 9953 8833
rect 10151 8807 10177 8833
rect 10599 8807 10625 8833
rect 10823 8807 10849 8833
rect 10935 8807 10961 8833
rect 11103 8807 11129 8833
rect 11551 8807 11577 8833
rect 13343 8807 13369 8833
rect 13455 8807 13481 8833
rect 13623 8807 13649 8833
rect 13735 8807 13761 8833
rect 13903 8807 13929 8833
rect 14071 8807 14097 8833
rect 14295 8807 14321 8833
rect 18831 8807 18857 8833
rect 6063 8751 6089 8777
rect 8583 8751 8609 8777
rect 8919 8751 8945 8777
rect 10319 8751 10345 8777
rect 11271 8751 11297 8777
rect 14127 8751 14153 8777
rect 14239 8751 14265 8777
rect 6791 8695 6817 8721
rect 7127 8695 7153 8721
rect 10375 8695 10401 8721
rect 10767 8695 10793 8721
rect 13903 8695 13929 8721
rect 9919 8611 9945 8637
rect 9971 8611 9997 8637
rect 10023 8611 10049 8637
rect 5895 8527 5921 8553
rect 6959 8527 6985 8553
rect 7015 8527 7041 8553
rect 7855 8527 7881 8553
rect 8751 8527 8777 8553
rect 9759 8527 9785 8553
rect 10375 8527 10401 8553
rect 10543 8527 10569 8553
rect 10711 8527 10737 8553
rect 10879 8527 10905 8553
rect 7575 8471 7601 8497
rect 7911 8471 7937 8497
rect 8695 8471 8721 8497
rect 11383 8471 11409 8497
rect 11551 8471 11577 8497
rect 13847 8471 13873 8497
rect 2143 8415 2169 8441
rect 5783 8415 5809 8441
rect 7071 8415 7097 8441
rect 7295 8415 7321 8441
rect 7463 8415 7489 8441
rect 7743 8415 7769 8441
rect 9199 8415 9225 8441
rect 9591 8415 9617 8441
rect 10095 8415 10121 8441
rect 10991 8415 11017 8441
rect 13063 8415 13089 8441
rect 13287 8415 13313 8441
rect 13455 8415 13481 8441
rect 18943 8415 18969 8441
rect 9031 8359 9057 8385
rect 9535 8359 9561 8385
rect 14911 8359 14937 8385
rect 20007 8359 20033 8385
rect 967 8303 993 8329
rect 8751 8303 8777 8329
rect 2239 8219 2265 8245
rect 2291 8219 2317 8245
rect 2343 8219 2369 8245
rect 17599 8219 17625 8245
rect 17651 8219 17677 8245
rect 17703 8219 17729 8245
rect 6791 8135 6817 8161
rect 9983 8079 10009 8105
rect 6959 8023 6985 8049
rect 7239 8023 7265 8049
rect 7743 8023 7769 8049
rect 10207 8023 10233 8049
rect 10599 8023 10625 8049
rect 10767 8023 10793 8049
rect 12503 8023 12529 8049
rect 6791 7911 6817 7937
rect 6847 7939 6873 7965
rect 7183 7967 7209 7993
rect 7687 7967 7713 7993
rect 7071 7911 7097 7937
rect 7575 7911 7601 7937
rect 10879 7911 10905 7937
rect 10935 7911 10961 7937
rect 12335 7911 12361 7937
rect 12447 7911 12473 7937
rect 9919 7827 9945 7853
rect 9971 7827 9997 7853
rect 10023 7827 10049 7853
rect 6399 7687 6425 7713
rect 7351 7687 7377 7713
rect 8751 7687 8777 7713
rect 8807 7687 8833 7713
rect 12111 7687 12137 7713
rect 6791 7631 6817 7657
rect 7015 7631 7041 7657
rect 8639 7631 8665 7657
rect 10095 7631 10121 7657
rect 10319 7631 10345 7657
rect 10655 7631 10681 7657
rect 10711 7631 10737 7657
rect 10823 7631 10849 7657
rect 10935 7631 10961 7657
rect 11887 7631 11913 7657
rect 11999 7631 12025 7657
rect 12167 7631 12193 7657
rect 5335 7575 5361 7601
rect 8415 7575 8441 7601
rect 9031 7575 9057 7601
rect 10207 7575 10233 7601
rect 10879 7575 10905 7601
rect 10039 7519 10065 7545
rect 2239 7435 2265 7461
rect 2291 7435 2317 7461
rect 2343 7435 2369 7461
rect 17599 7435 17625 7461
rect 17651 7435 17677 7461
rect 17703 7435 17729 7461
rect 9871 7351 9897 7377
rect 6903 7295 6929 7321
rect 8583 7295 8609 7321
rect 9647 7295 9673 7321
rect 9815 7295 9841 7321
rect 10095 7295 10121 7321
rect 12055 7295 12081 7321
rect 13119 7295 13145 7321
rect 8247 7239 8273 7265
rect 11663 7239 11689 7265
rect 10711 7183 10737 7209
rect 10767 7183 10793 7209
rect 10599 7127 10625 7153
rect 13343 7127 13369 7153
rect 9919 7043 9945 7069
rect 9971 7043 9997 7069
rect 10023 7043 10049 7069
rect 12223 6959 12249 6985
rect 12895 6959 12921 6985
rect 8359 6903 8385 6929
rect 8415 6903 8441 6929
rect 10095 6903 10121 6929
rect 12615 6903 12641 6929
rect 12671 6903 12697 6929
rect 13063 6903 13089 6929
rect 8247 6847 8273 6873
rect 9759 6847 9785 6873
rect 11999 6847 12025 6873
rect 12279 6847 12305 6873
rect 12783 6847 12809 6873
rect 11159 6791 11185 6817
rect 11383 6791 11409 6817
rect 12223 6735 12249 6761
rect 2239 6651 2265 6677
rect 2291 6651 2317 6677
rect 2343 6651 2369 6677
rect 17599 6651 17625 6677
rect 17651 6651 17677 6677
rect 17703 6651 17729 6677
rect 8919 6567 8945 6593
rect 10767 6567 10793 6593
rect 7631 6511 7657 6537
rect 8695 6511 8721 6537
rect 9199 6511 9225 6537
rect 11047 6511 11073 6537
rect 12223 6511 12249 6537
rect 13287 6511 13313 6537
rect 13511 6511 13537 6537
rect 7295 6455 7321 6481
rect 8975 6455 9001 6481
rect 10823 6455 10849 6481
rect 11831 6455 11857 6481
rect 8919 6343 8945 6369
rect 10767 6343 10793 6369
rect 9919 6259 9945 6285
rect 9971 6259 9997 6285
rect 10023 6259 10049 6285
rect 8863 6175 8889 6201
rect 11439 6175 11465 6201
rect 10151 6119 10177 6145
rect 9759 6063 9785 6089
rect 11215 6007 11241 6033
rect 2239 5867 2265 5893
rect 2291 5867 2317 5893
rect 2343 5867 2369 5893
rect 17599 5867 17625 5893
rect 17651 5867 17677 5893
rect 17703 5867 17729 5893
rect 9919 5475 9945 5501
rect 9971 5475 9997 5501
rect 10023 5475 10049 5501
rect 2239 5083 2265 5109
rect 2291 5083 2317 5109
rect 2343 5083 2369 5109
rect 17599 5083 17625 5109
rect 17651 5083 17677 5109
rect 17703 5083 17729 5109
rect 9919 4691 9945 4717
rect 9971 4691 9997 4717
rect 10023 4691 10049 4717
rect 2239 4299 2265 4325
rect 2291 4299 2317 4325
rect 2343 4299 2369 4325
rect 17599 4299 17625 4325
rect 17651 4299 17677 4325
rect 17703 4299 17729 4325
rect 9919 3907 9945 3933
rect 9971 3907 9997 3933
rect 10023 3907 10049 3933
rect 2239 3515 2265 3541
rect 2291 3515 2317 3541
rect 2343 3515 2369 3541
rect 17599 3515 17625 3541
rect 17651 3515 17677 3541
rect 17703 3515 17729 3541
rect 9919 3123 9945 3149
rect 9971 3123 9997 3149
rect 10023 3123 10049 3149
rect 2239 2731 2265 2757
rect 2291 2731 2317 2757
rect 2343 2731 2369 2757
rect 17599 2731 17625 2757
rect 17651 2731 17677 2757
rect 17703 2731 17729 2757
rect 9919 2339 9945 2365
rect 9971 2339 9997 2365
rect 10023 2339 10049 2365
rect 10935 2143 10961 2169
rect 12895 2143 12921 2169
rect 11383 2031 11409 2057
rect 13399 2031 13425 2057
rect 2239 1947 2265 1973
rect 2291 1947 2317 1973
rect 2343 1947 2369 1973
rect 17599 1947 17625 1973
rect 17651 1947 17677 1973
rect 17703 1947 17729 1973
rect 13063 1807 13089 1833
rect 14687 1807 14713 1833
rect 8527 1751 8553 1777
rect 10711 1751 10737 1777
rect 12615 1751 12641 1777
rect 14295 1751 14321 1777
rect 9031 1639 9057 1665
rect 11215 1639 11241 1665
rect 9919 1555 9945 1581
rect 9971 1555 9997 1581
rect 10023 1555 10049 1581
<< metal2 >>
rect 8736 20600 8792 21000
rect 9408 20600 9464 21000
rect 10080 20600 10136 21000
rect 11760 20600 11816 21000
rect 12096 20600 12152 21000
rect 2238 19222 2370 19227
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2238 19189 2370 19194
rect 8750 19138 8778 20600
rect 8750 19105 8778 19110
rect 9310 19138 9338 19143
rect 9310 19091 9338 19110
rect 8806 19025 8834 19031
rect 8806 18999 8807 19025
rect 8833 18999 8834 19025
rect 2238 18438 2370 18443
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2238 18405 2370 18410
rect 2238 17654 2370 17659
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2238 17621 2370 17626
rect 2238 16870 2370 16875
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2238 16837 2370 16842
rect 2238 16086 2370 16091
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2238 16053 2370 16058
rect 8806 15974 8834 18999
rect 9422 18746 9450 20600
rect 10094 19138 10122 20600
rect 10094 19105 10122 19110
rect 10878 19138 10906 19143
rect 10878 19091 10906 19110
rect 11774 19138 11802 20600
rect 11774 19105 11802 19110
rect 10374 19025 10402 19031
rect 10374 18999 10375 19025
rect 10401 18999 10402 19025
rect 9918 18830 10050 18835
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 9918 18797 10050 18802
rect 9422 18713 9450 18718
rect 10038 18746 10066 18751
rect 10038 18699 10066 18718
rect 9534 18633 9562 18639
rect 9534 18607 9535 18633
rect 9561 18607 9562 18633
rect 9534 15974 9562 18607
rect 9918 18046 10050 18051
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 9918 18013 10050 18018
rect 9918 17262 10050 17267
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 9918 17229 10050 17234
rect 9918 16478 10050 16483
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 9918 16445 10050 16450
rect 10374 15974 10402 18999
rect 12110 18746 12138 20600
rect 17598 19222 17730 19227
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17598 19189 17730 19194
rect 12782 19138 12810 19143
rect 12782 19091 12810 19110
rect 12110 18713 12138 18718
rect 12278 19025 12306 19031
rect 12278 18999 12279 19025
rect 12305 18999 12306 19025
rect 12278 15974 12306 18999
rect 13118 18746 13146 18751
rect 13118 18699 13146 18718
rect 8638 15946 8834 15974
rect 9478 15946 9562 15974
rect 10150 15946 10402 15974
rect 11830 15946 12306 15974
rect 12614 18633 12642 18639
rect 12614 18607 12615 18633
rect 12641 18607 12642 18633
rect 2238 15302 2370 15307
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2238 15269 2370 15274
rect 2238 14518 2370 14523
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2238 14485 2370 14490
rect 8470 13873 8498 13879
rect 8470 13847 8471 13873
rect 8497 13847 8498 13873
rect 2086 13818 2114 13823
rect 966 12250 994 12255
rect 966 12203 994 12222
rect 966 12025 994 12031
rect 966 11999 967 12025
rect 993 11999 994 12025
rect 966 11802 994 11999
rect 966 11769 994 11774
rect 2086 9954 2114 13790
rect 2238 13734 2370 13739
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2238 13701 2370 13706
rect 8078 13537 8106 13543
rect 8078 13511 8079 13537
rect 8105 13511 8106 13537
rect 8078 13482 8106 13511
rect 8078 13449 8106 13454
rect 8414 13481 8442 13487
rect 8414 13455 8415 13481
rect 8441 13455 8442 13481
rect 8414 13090 8442 13455
rect 8470 13482 8498 13847
rect 8470 13449 8498 13454
rect 8414 13057 8442 13062
rect 2238 12950 2370 12955
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2238 12917 2370 12922
rect 8638 12810 8666 15946
rect 8806 13930 8834 13935
rect 8806 13929 8890 13930
rect 8806 13903 8807 13929
rect 8833 13903 8890 13929
rect 8806 13902 8890 13903
rect 8806 13897 8834 13902
rect 8862 13482 8890 13902
rect 9142 13874 9170 13879
rect 9142 13827 9170 13846
rect 9478 13650 9506 15946
rect 9918 15694 10050 15699
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 9918 15661 10050 15666
rect 9918 14910 10050 14915
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 9918 14877 10050 14882
rect 10150 14265 10178 15946
rect 10150 14239 10151 14265
rect 10177 14239 10178 14265
rect 10038 14210 10066 14215
rect 10038 14209 10122 14210
rect 10038 14183 10039 14209
rect 10065 14183 10122 14209
rect 10038 14182 10122 14183
rect 10038 14177 10066 14182
rect 9918 14126 10050 14131
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 9918 14093 10050 14098
rect 10094 14042 10122 14182
rect 10038 14014 10122 14042
rect 9926 13874 9954 13879
rect 9478 13622 9898 13650
rect 9478 13593 9506 13622
rect 9478 13567 9479 13593
rect 9505 13567 9506 13593
rect 9478 13561 9506 13567
rect 9814 13538 9842 13543
rect 9758 13537 9842 13538
rect 9758 13511 9815 13537
rect 9841 13511 9842 13537
rect 9758 13510 9842 13511
rect 8638 12809 8722 12810
rect 8638 12783 8639 12809
rect 8665 12783 8722 12809
rect 8638 12782 8722 12783
rect 8638 12777 8666 12782
rect 7182 12753 7210 12759
rect 7182 12727 7183 12753
rect 7209 12727 7210 12753
rect 2142 12362 2170 12367
rect 2142 12315 2170 12334
rect 6902 12362 6930 12367
rect 6902 12305 6930 12334
rect 6902 12279 6903 12305
rect 6929 12279 6930 12305
rect 6902 12273 6930 12279
rect 7182 12362 7210 12727
rect 7574 12698 7602 12703
rect 7574 12697 8274 12698
rect 7574 12671 7575 12697
rect 7601 12671 8274 12697
rect 7574 12670 8274 12671
rect 7574 12665 7602 12670
rect 2238 12166 2370 12171
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2238 12133 2370 12138
rect 2142 11969 2170 11975
rect 2142 11943 2143 11969
rect 2169 11943 2170 11969
rect 2142 11522 2170 11943
rect 6790 11913 6818 11919
rect 6790 11887 6791 11913
rect 6817 11887 6818 11913
rect 6734 11857 6762 11863
rect 6734 11831 6735 11857
rect 6761 11831 6762 11857
rect 6734 11633 6762 11831
rect 6790 11690 6818 11887
rect 6790 11657 6818 11662
rect 6734 11607 6735 11633
rect 6761 11607 6762 11633
rect 6734 11601 6762 11607
rect 2142 11489 2170 11494
rect 5670 11578 5698 11583
rect 5670 11521 5698 11550
rect 5670 11495 5671 11521
rect 5697 11495 5698 11521
rect 5670 11489 5698 11495
rect 7126 11578 7154 11583
rect 7182 11578 7210 12334
rect 7966 12305 7994 12311
rect 7966 12279 7967 12305
rect 7993 12279 7994 12305
rect 7966 12025 7994 12279
rect 8246 12081 8274 12670
rect 8414 12474 8442 12479
rect 8302 12362 8330 12367
rect 8302 12315 8330 12334
rect 8246 12055 8247 12081
rect 8273 12055 8274 12081
rect 8246 12049 8274 12055
rect 8414 12081 8442 12446
rect 8414 12055 8415 12081
rect 8441 12055 8442 12081
rect 8414 12049 8442 12055
rect 8638 12306 8666 12311
rect 7966 11999 7967 12025
rect 7993 11999 7994 12025
rect 7966 11993 7994 11999
rect 7910 11969 7938 11975
rect 7910 11943 7911 11969
rect 7937 11943 7938 11969
rect 7686 11746 7714 11751
rect 7574 11690 7602 11695
rect 7574 11643 7602 11662
rect 7686 11689 7714 11718
rect 7910 11746 7938 11943
rect 8638 11970 8666 12278
rect 8694 12250 8722 12782
rect 8862 12641 8890 13454
rect 9702 13482 9730 13487
rect 9702 13435 9730 13454
rect 9702 13258 9730 13263
rect 9534 13257 9730 13258
rect 9534 13231 9703 13257
rect 9729 13231 9730 13257
rect 9534 13230 9730 13231
rect 9534 13202 9562 13230
rect 9702 13225 9730 13230
rect 9478 13174 9562 13202
rect 9366 13146 9394 13151
rect 8862 12615 8863 12641
rect 8889 12615 8890 12641
rect 8750 12362 8778 12367
rect 8862 12362 8890 12615
rect 9254 12753 9282 12759
rect 9254 12727 9255 12753
rect 9281 12727 9282 12753
rect 9086 12586 9114 12591
rect 9086 12417 9114 12558
rect 9142 12474 9170 12479
rect 9142 12427 9170 12446
rect 9086 12391 9087 12417
rect 9113 12391 9114 12417
rect 9086 12385 9114 12391
rect 8778 12334 8890 12362
rect 8918 12361 8946 12367
rect 8918 12335 8919 12361
rect 8945 12335 8946 12361
rect 8750 12315 8778 12334
rect 8918 12250 8946 12335
rect 8694 12222 8946 12250
rect 9198 12249 9226 12255
rect 9198 12223 9199 12249
rect 9225 12223 9226 12249
rect 9198 12082 9226 12223
rect 9030 12054 9226 12082
rect 8694 11970 8722 11975
rect 8638 11969 8722 11970
rect 8638 11943 8695 11969
rect 8721 11943 8722 11969
rect 8638 11942 8722 11943
rect 8694 11937 8722 11942
rect 8918 11970 8946 11989
rect 8918 11937 8946 11942
rect 8974 11970 9002 11975
rect 9030 11970 9058 12054
rect 8974 11969 9058 11970
rect 8974 11943 8975 11969
rect 9001 11943 9058 11969
rect 8974 11942 9058 11943
rect 9086 11969 9114 11975
rect 9086 11943 9087 11969
rect 9113 11943 9114 11969
rect 8078 11913 8106 11919
rect 8078 11887 8079 11913
rect 8105 11887 8106 11913
rect 8078 11858 8106 11887
rect 8078 11825 8106 11830
rect 8302 11857 8330 11863
rect 8302 11831 8303 11857
rect 8329 11831 8330 11857
rect 7910 11713 7938 11718
rect 8302 11746 8330 11831
rect 8918 11858 8946 11863
rect 8918 11811 8946 11830
rect 7686 11663 7687 11689
rect 7713 11663 7714 11689
rect 7686 11657 7714 11663
rect 7630 11634 7658 11639
rect 7126 11577 7210 11578
rect 7126 11551 7127 11577
rect 7153 11551 7210 11577
rect 7126 11550 7210 11551
rect 7406 11578 7434 11583
rect 2238 11382 2370 11387
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2238 11349 2370 11354
rect 6454 10794 6482 10799
rect 2238 10598 2370 10603
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2238 10565 2370 10570
rect 6454 10457 6482 10766
rect 6454 10431 6455 10457
rect 6481 10431 6482 10457
rect 6454 10425 6482 10431
rect 6510 10737 6538 10743
rect 6510 10711 6511 10737
rect 6537 10711 6538 10737
rect 5054 10401 5082 10407
rect 5054 10375 5055 10401
rect 5081 10375 5082 10401
rect 5054 10122 5082 10375
rect 6510 10402 6538 10711
rect 5390 10346 5418 10351
rect 5390 10299 5418 10318
rect 6510 10094 6538 10374
rect 5054 10009 5082 10094
rect 6454 10066 6538 10094
rect 6678 10737 6706 10743
rect 6678 10711 6679 10737
rect 6705 10711 6706 10737
rect 5054 9983 5055 10009
rect 5081 9983 5082 10009
rect 5054 9977 5082 9983
rect 5390 10010 5418 10015
rect 5390 9963 5418 9982
rect 2086 9921 2114 9926
rect 6454 9953 6482 10066
rect 6678 10009 6706 10711
rect 6902 10738 6930 10743
rect 7126 10738 7154 11550
rect 7406 11531 7434 11550
rect 7518 11577 7546 11583
rect 7518 11551 7519 11577
rect 7545 11551 7546 11577
rect 7518 11354 7546 11551
rect 7518 11321 7546 11326
rect 7238 11073 7266 11079
rect 7238 11047 7239 11073
rect 7265 11047 7266 11073
rect 7238 10738 7266 11047
rect 7462 10906 7490 10911
rect 7630 10906 7658 11606
rect 7966 11521 7994 11527
rect 7966 11495 7967 11521
rect 7993 11495 7994 11521
rect 7966 11410 7994 11495
rect 7966 11377 7994 11382
rect 8302 11298 8330 11718
rect 8302 11265 8330 11270
rect 8358 11634 8386 11639
rect 7462 10905 7658 10906
rect 7462 10879 7463 10905
rect 7489 10879 7658 10905
rect 7462 10878 7658 10879
rect 7686 10906 7714 10911
rect 7462 10873 7490 10878
rect 7294 10794 7322 10799
rect 7322 10766 7378 10794
rect 7294 10747 7322 10766
rect 6902 10737 7266 10738
rect 6902 10711 6903 10737
rect 6929 10711 7266 10737
rect 6902 10710 7266 10711
rect 6790 10402 6818 10407
rect 6790 10355 6818 10374
rect 6902 10122 6930 10710
rect 7238 10458 7266 10710
rect 7238 10425 7266 10430
rect 7294 10346 7322 10351
rect 7294 10299 7322 10318
rect 6958 10289 6986 10295
rect 6958 10263 6959 10289
rect 6985 10263 6986 10289
rect 6958 10178 6986 10263
rect 6958 10145 6986 10150
rect 7350 10121 7378 10766
rect 7462 10290 7490 10295
rect 7350 10095 7351 10121
rect 7377 10095 7378 10121
rect 7350 10094 7378 10095
rect 6790 10066 6818 10071
rect 6678 9983 6679 10009
rect 6705 9983 6706 10009
rect 6678 9977 6706 9983
rect 6734 10065 6818 10066
rect 6734 10039 6791 10065
rect 6817 10039 6818 10065
rect 6734 10038 6818 10039
rect 6734 10010 6762 10038
rect 6790 10033 6818 10038
rect 6454 9927 6455 9953
rect 6481 9927 6482 9953
rect 6454 9921 6482 9927
rect 2238 9814 2370 9819
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2238 9781 2370 9786
rect 6734 9394 6762 9982
rect 6734 9361 6762 9366
rect 6790 9506 6818 9511
rect 6902 9506 6930 10094
rect 7070 10066 7378 10094
rect 7406 10289 7490 10290
rect 7406 10263 7463 10289
rect 7489 10263 7490 10289
rect 7406 10262 7490 10263
rect 7070 10009 7098 10066
rect 7070 9983 7071 10009
rect 7097 9983 7098 10009
rect 7070 9977 7098 9983
rect 7182 9954 7210 9959
rect 7406 9954 7434 10262
rect 7462 10257 7490 10262
rect 7182 9953 7434 9954
rect 7182 9927 7183 9953
rect 7209 9927 7434 9953
rect 7182 9926 7434 9927
rect 7182 9921 7210 9926
rect 7406 9730 7434 9926
rect 7350 9702 7434 9730
rect 7462 10122 7490 10127
rect 6790 9505 6930 9506
rect 6790 9479 6791 9505
rect 6817 9479 6930 9505
rect 6790 9478 6930 9479
rect 7294 9618 7322 9623
rect 2238 9030 2370 9035
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2238 8997 2370 9002
rect 966 8890 994 8895
rect 966 8843 994 8862
rect 4998 8889 5026 8895
rect 4998 8863 4999 8889
rect 5025 8863 5026 8889
rect 2142 8834 2170 8839
rect 2142 8787 2170 8806
rect 4998 8834 5026 8863
rect 2142 8441 2170 8447
rect 2142 8415 2143 8441
rect 2169 8415 2170 8441
rect 966 8329 994 8335
rect 966 8303 967 8329
rect 993 8303 994 8329
rect 966 8106 994 8303
rect 966 8073 994 8078
rect 2142 7602 2170 8415
rect 4998 8442 5026 8806
rect 6398 8834 6426 8839
rect 6398 8787 6426 8806
rect 6734 8834 6762 8839
rect 6062 8778 6090 8783
rect 5894 8777 6090 8778
rect 5894 8751 6063 8777
rect 6089 8751 6090 8777
rect 5894 8750 6090 8751
rect 4998 8409 5026 8414
rect 5782 8722 5810 8727
rect 5782 8441 5810 8694
rect 5894 8553 5922 8750
rect 6062 8745 6090 8750
rect 5894 8527 5895 8553
rect 5921 8527 5922 8553
rect 5894 8521 5922 8527
rect 6734 8722 6762 8806
rect 6790 8722 6818 9478
rect 7126 9394 7154 9399
rect 7126 9225 7154 9366
rect 7126 9199 7127 9225
rect 7153 9199 7154 9225
rect 7126 9193 7154 9199
rect 7238 9226 7266 9231
rect 7294 9226 7322 9590
rect 7350 9506 7378 9702
rect 7406 9618 7434 9623
rect 7462 9618 7490 10094
rect 7574 9954 7602 9959
rect 7406 9617 7490 9618
rect 7406 9591 7407 9617
rect 7433 9591 7490 9617
rect 7406 9590 7490 9591
rect 7518 9953 7602 9954
rect 7518 9927 7575 9953
rect 7601 9927 7602 9953
rect 7518 9926 7602 9927
rect 7406 9585 7434 9590
rect 7406 9506 7434 9511
rect 7518 9506 7546 9926
rect 7574 9921 7602 9926
rect 7350 9478 7406 9506
rect 7406 9473 7434 9478
rect 7462 9505 7546 9506
rect 7462 9479 7519 9505
rect 7545 9479 7546 9505
rect 7462 9478 7546 9479
rect 7238 9225 7322 9226
rect 7238 9199 7239 9225
rect 7265 9199 7322 9225
rect 7238 9198 7322 9199
rect 7462 9282 7490 9478
rect 7518 9473 7546 9478
rect 7574 9505 7602 9511
rect 7574 9479 7575 9505
rect 7601 9479 7602 9505
rect 7574 9394 7602 9479
rect 7462 9225 7490 9254
rect 7462 9199 7463 9225
rect 7489 9199 7490 9225
rect 7238 9193 7266 9198
rect 7462 9193 7490 9199
rect 7518 9366 7602 9394
rect 6958 9114 6986 9119
rect 7406 9114 7434 9119
rect 6958 9113 7098 9114
rect 6958 9087 6959 9113
rect 6985 9087 7098 9113
rect 6958 9086 7098 9087
rect 6958 9081 6986 9086
rect 7070 9002 7098 9086
rect 7294 9113 7434 9114
rect 7294 9087 7407 9113
rect 7433 9087 7434 9113
rect 7294 9086 7434 9087
rect 7070 8974 7210 9002
rect 6734 8721 6818 8722
rect 6734 8695 6791 8721
rect 6817 8695 6818 8721
rect 6734 8694 6818 8695
rect 5782 8415 5783 8441
rect 5809 8415 5810 8441
rect 5782 8409 5810 8415
rect 2238 8246 2370 8251
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2238 8213 2370 8218
rect 6398 7938 6426 7943
rect 2142 7569 2170 7574
rect 5334 7770 5362 7775
rect 5334 7602 5362 7742
rect 6398 7713 6426 7910
rect 6398 7687 6399 7713
rect 6425 7687 6426 7713
rect 6398 7681 6426 7687
rect 6734 7658 6762 8694
rect 6790 8689 6818 8694
rect 6958 8918 7154 8946
rect 6958 8553 6986 8918
rect 7070 8833 7098 8839
rect 7070 8807 7071 8833
rect 7097 8807 7098 8833
rect 6958 8527 6959 8553
rect 6985 8527 6986 8553
rect 6958 8521 6986 8527
rect 7014 8554 7042 8559
rect 7070 8554 7098 8807
rect 7126 8834 7154 8918
rect 7182 8945 7210 8974
rect 7294 8946 7322 9086
rect 7406 9081 7434 9086
rect 7182 8919 7183 8945
rect 7209 8919 7210 8945
rect 7182 8913 7210 8919
rect 7238 8918 7322 8946
rect 7238 8834 7266 8918
rect 7350 8890 7378 8895
rect 7126 8806 7266 8834
rect 7294 8862 7350 8890
rect 7294 8833 7322 8862
rect 7350 8857 7378 8862
rect 7294 8807 7295 8833
rect 7321 8807 7322 8833
rect 7294 8778 7322 8807
rect 7238 8750 7322 8778
rect 7406 8833 7434 8839
rect 7406 8807 7407 8833
rect 7433 8807 7434 8833
rect 7406 8778 7434 8807
rect 7126 8722 7154 8727
rect 7126 8675 7154 8694
rect 7014 8553 7098 8554
rect 7014 8527 7015 8553
rect 7041 8527 7098 8553
rect 7014 8526 7098 8527
rect 7014 8521 7042 8526
rect 7126 8498 7154 8503
rect 7070 8442 7098 8447
rect 7070 8395 7098 8414
rect 7126 8330 7154 8470
rect 7014 8302 7154 8330
rect 6790 8161 6818 8167
rect 6790 8135 6791 8161
rect 6817 8135 6818 8161
rect 6790 8106 6818 8135
rect 6790 8078 6986 8106
rect 6958 8049 6986 8078
rect 6958 8023 6959 8049
rect 6985 8023 6986 8049
rect 6958 8017 6986 8023
rect 6846 7965 6874 7971
rect 6790 7937 6818 7943
rect 6790 7911 6791 7937
rect 6817 7911 6818 7937
rect 6790 7770 6818 7911
rect 6846 7939 6847 7965
rect 6873 7939 6874 7965
rect 6846 7938 6874 7939
rect 7014 7938 7042 8302
rect 7238 8049 7266 8750
rect 7406 8745 7434 8750
rect 7294 8442 7322 8447
rect 7462 8442 7490 8447
rect 7518 8442 7546 9366
rect 7686 9226 7714 10878
rect 8358 10905 8386 11606
rect 8358 10879 8359 10905
rect 8385 10879 8386 10905
rect 8358 10873 8386 10879
rect 8806 11242 8834 11247
rect 8134 10850 8162 10855
rect 8134 10803 8162 10822
rect 8414 10850 8442 10855
rect 8414 10803 8442 10822
rect 8022 10794 8050 10799
rect 7742 10458 7770 10463
rect 7742 10411 7770 10430
rect 8022 10122 8050 10766
rect 8806 10793 8834 11214
rect 8918 10906 8946 10911
rect 8918 10859 8946 10878
rect 8806 10767 8807 10793
rect 8833 10767 8834 10793
rect 8806 10761 8834 10767
rect 8470 10738 8498 10743
rect 8358 10681 8386 10687
rect 8358 10655 8359 10681
rect 8385 10655 8386 10681
rect 8022 9618 8050 10094
rect 8078 10346 8106 10351
rect 8078 10009 8106 10318
rect 8078 9983 8079 10009
rect 8105 9983 8106 10009
rect 8078 9977 8106 9983
rect 8302 10009 8330 10015
rect 8302 9983 8303 10009
rect 8329 9983 8330 10009
rect 8246 9954 8274 9959
rect 8246 9907 8274 9926
rect 8302 9730 8330 9983
rect 8302 9697 8330 9702
rect 8134 9618 8162 9623
rect 8022 9617 8162 9618
rect 8022 9591 8135 9617
rect 8161 9591 8162 9617
rect 8022 9590 8162 9591
rect 8134 9585 8162 9590
rect 8190 9226 8218 9231
rect 7686 9225 7882 9226
rect 7686 9199 7687 9225
rect 7713 9199 7882 9225
rect 7686 9198 7882 9199
rect 7686 9193 7714 9198
rect 7574 9114 7602 9119
rect 7574 9067 7602 9086
rect 7854 8554 7882 9198
rect 7854 8507 7882 8526
rect 7910 9170 7938 9175
rect 7294 8441 7546 8442
rect 7294 8415 7295 8441
rect 7321 8415 7463 8441
rect 7489 8415 7546 8441
rect 7294 8414 7546 8415
rect 7574 8497 7602 8503
rect 7574 8471 7575 8497
rect 7601 8471 7602 8497
rect 7294 8409 7322 8414
rect 7462 8409 7490 8414
rect 7238 8023 7239 8049
rect 7265 8023 7266 8049
rect 7238 8017 7266 8023
rect 7574 8050 7602 8471
rect 7910 8497 7938 9142
rect 8190 9169 8218 9198
rect 8190 9143 8191 9169
rect 8217 9143 8218 9169
rect 8190 9137 8218 9143
rect 8358 9170 8386 10655
rect 8470 10121 8498 10710
rect 8974 10738 9002 11942
rect 9086 11690 9114 11943
rect 9198 11914 9226 11919
rect 9198 11867 9226 11886
rect 9198 11746 9226 11751
rect 9254 11746 9282 12727
rect 9366 12697 9394 13118
rect 9478 13145 9506 13174
rect 9478 13119 9479 13145
rect 9505 13119 9506 13145
rect 9478 13113 9506 13119
rect 9590 13145 9618 13151
rect 9590 13119 9591 13145
rect 9617 13119 9618 13145
rect 9534 13090 9562 13095
rect 9534 13043 9562 13062
rect 9590 12865 9618 13119
rect 9590 12839 9591 12865
rect 9617 12839 9618 12865
rect 9590 12833 9618 12839
rect 9758 12754 9786 13510
rect 9814 13505 9842 13510
rect 9870 13454 9898 13622
rect 9926 13593 9954 13846
rect 9926 13567 9927 13593
rect 9953 13567 9954 13593
rect 9926 13561 9954 13567
rect 10038 13537 10066 14014
rect 10150 13874 10178 14239
rect 10206 14266 10234 14271
rect 10878 14266 10906 14271
rect 10206 14265 10906 14266
rect 10206 14239 10207 14265
rect 10233 14239 10879 14265
rect 10905 14239 10906 14265
rect 10206 14238 10906 14239
rect 10206 14233 10234 14238
rect 10206 13874 10234 13879
rect 10150 13873 10234 13874
rect 10150 13847 10207 13873
rect 10233 13847 10234 13873
rect 10150 13846 10234 13847
rect 10206 13841 10234 13846
rect 10038 13511 10039 13537
rect 10065 13511 10066 13537
rect 10038 13505 10066 13511
rect 10094 13537 10122 13543
rect 10094 13511 10095 13537
rect 10121 13511 10122 13537
rect 9814 13426 9898 13454
rect 9814 13257 9842 13426
rect 9918 13342 10050 13347
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 9918 13309 10050 13314
rect 9814 13231 9815 13257
rect 9841 13231 9842 13257
rect 9814 13225 9842 13231
rect 9870 13146 9898 13151
rect 10094 13146 10122 13511
rect 9870 13145 9954 13146
rect 9870 13119 9871 13145
rect 9897 13119 9954 13145
rect 9870 13118 9954 13119
rect 9870 13113 9898 13118
rect 9926 13034 9954 13118
rect 10094 13113 10122 13118
rect 10262 13034 10290 14238
rect 10878 14233 10906 14238
rect 10934 14266 10962 14271
rect 10934 14219 10962 14238
rect 11830 14266 11858 15946
rect 12614 14266 12642 18607
rect 17598 18438 17730 18443
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17598 18405 17730 18410
rect 17598 17654 17730 17659
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17598 17621 17730 17626
rect 17598 16870 17730 16875
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17598 16837 17730 16842
rect 17598 16086 17730 16091
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17598 16053 17730 16058
rect 17598 15302 17730 15307
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17598 15269 17730 15274
rect 17598 14518 17730 14523
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17598 14485 17730 14490
rect 11046 14210 11074 14215
rect 10990 14209 11074 14210
rect 10990 14183 11047 14209
rect 11073 14183 11074 14209
rect 10990 14182 11074 14183
rect 10430 13929 10458 13935
rect 10430 13903 10431 13929
rect 10457 13903 10458 13929
rect 10430 13538 10458 13903
rect 10766 13874 10794 13879
rect 10430 13505 10458 13510
rect 10710 13873 10794 13874
rect 10710 13847 10767 13873
rect 10793 13847 10794 13873
rect 10710 13846 10794 13847
rect 10710 13257 10738 13846
rect 10766 13841 10794 13846
rect 10990 13706 11018 14182
rect 11046 14177 11074 14182
rect 11830 13873 11858 14238
rect 12334 14238 12642 14266
rect 11830 13847 11831 13873
rect 11857 13847 11858 13873
rect 11830 13841 11858 13847
rect 12110 13873 12138 13879
rect 12110 13847 12111 13873
rect 12137 13847 12138 13873
rect 10710 13231 10711 13257
rect 10737 13231 10738 13257
rect 10710 13225 10738 13231
rect 10766 13678 11018 13706
rect 10766 13201 10794 13678
rect 11886 13594 11914 13599
rect 10934 13538 10962 13543
rect 10934 13491 10962 13510
rect 11270 13481 11298 13487
rect 11270 13455 11271 13481
rect 11297 13455 11298 13481
rect 11270 13257 11298 13455
rect 11270 13231 11271 13257
rect 11297 13231 11298 13257
rect 11270 13225 11298 13231
rect 11886 13257 11914 13566
rect 12110 13538 12138 13847
rect 12334 13594 12362 14238
rect 17598 13734 17730 13739
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17598 13701 17730 13706
rect 12334 13547 12362 13566
rect 14294 13593 14322 13599
rect 14294 13567 14295 13593
rect 14321 13567 14322 13593
rect 12110 13505 12138 13510
rect 12558 13538 12586 13543
rect 12558 13491 12586 13510
rect 12894 13538 12922 13543
rect 14294 13538 14322 13567
rect 20006 13593 20034 13599
rect 20006 13567 20007 13593
rect 20033 13567 20034 13593
rect 14350 13538 14378 13543
rect 14294 13510 14350 13538
rect 12894 13454 12922 13510
rect 14350 13505 14378 13510
rect 14574 13538 14602 13543
rect 13230 13481 13258 13487
rect 13230 13455 13231 13481
rect 13257 13455 13258 13481
rect 12894 13426 12978 13454
rect 11886 13231 11887 13257
rect 11913 13231 11914 13257
rect 11886 13225 11914 13231
rect 10766 13175 10767 13201
rect 10793 13175 10794 13201
rect 10766 13169 10794 13175
rect 10878 13202 10906 13207
rect 11046 13202 11074 13207
rect 10906 13201 11074 13202
rect 10906 13175 11047 13201
rect 11073 13175 11074 13201
rect 10906 13174 11074 13175
rect 10878 13155 10906 13174
rect 11046 13169 11074 13174
rect 9926 13006 10290 13034
rect 9758 12726 9842 12754
rect 9366 12671 9367 12697
rect 9393 12671 9394 12697
rect 9366 12665 9394 12671
rect 9646 12641 9674 12647
rect 9646 12615 9647 12641
rect 9673 12615 9674 12641
rect 9646 12474 9674 12615
rect 9646 12441 9674 12446
rect 9702 12642 9730 12647
rect 9758 12642 9786 12647
rect 9730 12641 9786 12642
rect 9730 12615 9759 12641
rect 9785 12615 9786 12641
rect 9730 12614 9786 12615
rect 9422 12361 9450 12367
rect 9422 12335 9423 12361
rect 9449 12335 9450 12361
rect 9310 12305 9338 12311
rect 9310 12279 9311 12305
rect 9337 12279 9338 12305
rect 9310 11914 9338 12279
rect 9310 11881 9338 11886
rect 9226 11718 9282 11746
rect 9198 11713 9226 11718
rect 9086 11657 9114 11662
rect 9142 11578 9170 11583
rect 9142 11577 9338 11578
rect 9142 11551 9143 11577
rect 9169 11551 9338 11577
rect 9142 11550 9338 11551
rect 9086 11298 9114 11303
rect 9086 11251 9114 11270
rect 9142 10905 9170 11550
rect 9142 10879 9143 10905
rect 9169 10879 9170 10905
rect 9142 10873 9170 10879
rect 9198 11242 9226 11247
rect 9086 10794 9114 10799
rect 9086 10747 9114 10766
rect 8974 10705 9002 10710
rect 8470 10095 8471 10121
rect 8497 10095 8498 10121
rect 8470 10089 8498 10095
rect 8750 10122 8778 10127
rect 8526 9954 8554 9959
rect 8414 9730 8442 9735
rect 8414 9673 8442 9702
rect 8414 9647 8415 9673
rect 8441 9647 8442 9673
rect 8414 9641 8442 9647
rect 8358 9137 8386 9142
rect 8414 9225 8442 9231
rect 8414 9199 8415 9225
rect 8441 9199 8442 9225
rect 7910 8471 7911 8497
rect 7937 8471 7938 8497
rect 7910 8465 7938 8471
rect 8414 8498 8442 9199
rect 8526 8945 8554 9926
rect 8750 9337 8778 10094
rect 8806 10010 8834 10015
rect 8806 9963 8834 9982
rect 8974 9953 9002 9959
rect 8974 9927 8975 9953
rect 9001 9927 9002 9953
rect 8750 9311 8751 9337
rect 8777 9311 8778 9337
rect 8750 9305 8778 9311
rect 8918 9618 8946 9623
rect 8974 9618 9002 9927
rect 8918 9617 9002 9618
rect 8918 9591 8919 9617
rect 8945 9591 9002 9617
rect 8918 9590 9002 9591
rect 8862 9282 8890 9287
rect 8806 9254 8862 9282
rect 8526 8919 8527 8945
rect 8553 8919 8554 8945
rect 8526 8913 8554 8919
rect 8638 9170 8666 9175
rect 8582 8778 8610 8783
rect 8582 8731 8610 8750
rect 8638 8498 8666 9142
rect 8694 9169 8722 9175
rect 8694 9143 8695 9169
rect 8721 9143 8722 9169
rect 8694 8946 8722 9143
rect 8694 8913 8722 8918
rect 8694 8833 8722 8839
rect 8694 8807 8695 8833
rect 8721 8807 8722 8833
rect 8694 8722 8722 8807
rect 8806 8834 8834 9254
rect 8862 9249 8890 9254
rect 8918 9281 8946 9590
rect 9198 9561 9226 11214
rect 9310 11186 9338 11550
rect 9310 11139 9338 11158
rect 9366 11521 9394 11527
rect 9366 11495 9367 11521
rect 9393 11495 9394 11521
rect 9366 11466 9394 11495
rect 9254 10122 9282 10127
rect 9254 10075 9282 10094
rect 9310 9730 9338 9735
rect 9198 9535 9199 9561
rect 9225 9535 9226 9561
rect 9030 9394 9058 9399
rect 8918 9255 8919 9281
rect 8945 9255 8946 9281
rect 8862 8834 8890 8839
rect 8806 8833 8890 8834
rect 8806 8807 8863 8833
rect 8889 8807 8890 8833
rect 8806 8806 8890 8807
rect 8862 8801 8890 8806
rect 8918 8777 8946 9255
rect 8974 9282 9002 9287
rect 8974 9225 9002 9254
rect 8974 9199 8975 9225
rect 9001 9199 9002 9225
rect 8974 9193 9002 9199
rect 8918 8751 8919 8777
rect 8945 8751 8946 8777
rect 8918 8722 8946 8751
rect 8694 8694 8946 8722
rect 8974 8945 9002 8951
rect 8974 8919 8975 8945
rect 9001 8919 9002 8945
rect 8750 8554 8778 8559
rect 8750 8507 8778 8526
rect 8694 8498 8722 8503
rect 8974 8498 9002 8919
rect 8638 8497 8722 8498
rect 8638 8471 8695 8497
rect 8721 8471 8722 8497
rect 8638 8470 8722 8471
rect 7742 8441 7770 8447
rect 7742 8415 7743 8441
rect 7769 8415 7770 8441
rect 7574 8022 7658 8050
rect 7182 7994 7210 7999
rect 7630 7994 7658 8022
rect 7742 8049 7770 8415
rect 7742 8023 7743 8049
rect 7769 8023 7770 8049
rect 7742 8017 7770 8023
rect 7686 7994 7714 7999
rect 7630 7966 7686 7994
rect 7182 7947 7210 7966
rect 7686 7947 7714 7966
rect 6846 7910 7042 7938
rect 7070 7938 7098 7943
rect 7574 7938 7602 7943
rect 7070 7891 7098 7910
rect 7350 7937 7602 7938
rect 7350 7911 7575 7937
rect 7601 7911 7602 7937
rect 7350 7910 7602 7911
rect 6790 7737 6818 7742
rect 7350 7713 7378 7910
rect 7574 7905 7602 7910
rect 7350 7687 7351 7713
rect 7377 7687 7378 7713
rect 7350 7681 7378 7687
rect 6790 7658 6818 7663
rect 6734 7657 6818 7658
rect 6734 7631 6791 7657
rect 6817 7631 6818 7657
rect 6734 7630 6818 7631
rect 5334 7555 5362 7574
rect 2238 7462 2370 7467
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2238 7429 2370 7434
rect 6790 7322 6818 7630
rect 7014 7657 7042 7663
rect 7014 7631 7015 7657
rect 7041 7631 7042 7657
rect 6902 7322 6930 7327
rect 7014 7322 7042 7631
rect 8414 7601 8442 8470
rect 8694 8465 8722 8470
rect 8862 8470 9002 8498
rect 8750 8330 8778 8335
rect 8750 8329 8834 8330
rect 8750 8303 8751 8329
rect 8777 8303 8834 8329
rect 8750 8302 8834 8303
rect 8750 8297 8778 8302
rect 8750 7713 8778 7719
rect 8750 7687 8751 7713
rect 8777 7687 8778 7713
rect 8414 7575 8415 7601
rect 8441 7575 8442 7601
rect 8414 7569 8442 7575
rect 8638 7657 8666 7663
rect 8638 7631 8639 7657
rect 8665 7631 8666 7657
rect 8470 7546 8498 7551
rect 6790 7321 7014 7322
rect 6790 7295 6903 7321
rect 6929 7295 7014 7321
rect 6790 7294 7014 7295
rect 6902 7289 6930 7294
rect 7014 7289 7042 7294
rect 7294 7322 7322 7327
rect 2238 6678 2370 6683
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2238 6645 2370 6650
rect 7294 6481 7322 7294
rect 8246 7322 8274 7327
rect 8246 7265 8274 7294
rect 8246 7239 8247 7265
rect 8273 7239 8274 7265
rect 8246 7233 8274 7239
rect 8358 6929 8386 6935
rect 8358 6903 8359 6929
rect 8385 6903 8386 6929
rect 8246 6874 8274 6879
rect 7630 6873 8274 6874
rect 7630 6847 8247 6873
rect 8273 6847 8274 6873
rect 7630 6846 8274 6847
rect 7630 6537 7658 6846
rect 8246 6841 8274 6846
rect 8358 6594 8386 6903
rect 8414 6930 8442 6935
rect 8470 6930 8498 7518
rect 8582 7322 8610 7327
rect 8638 7322 8666 7631
rect 8750 7602 8778 7687
rect 8806 7713 8834 8302
rect 8806 7687 8807 7713
rect 8833 7687 8834 7713
rect 8806 7681 8834 7687
rect 8862 7602 8890 8470
rect 9030 8385 9058 9366
rect 9198 9226 9226 9535
rect 9198 8834 9226 9198
rect 9198 8801 9226 8806
rect 9254 9702 9310 9730
rect 9254 8833 9282 9702
rect 9310 9697 9338 9702
rect 9310 9226 9338 9231
rect 9366 9226 9394 11438
rect 9422 11354 9450 12335
rect 9534 11690 9562 11695
rect 9646 11690 9674 11695
rect 9534 11521 9562 11662
rect 9590 11662 9646 11690
rect 9590 11634 9618 11662
rect 9646 11657 9674 11662
rect 9590 11587 9618 11606
rect 9702 11578 9730 12614
rect 9758 12609 9786 12614
rect 9814 12026 9842 12726
rect 9870 12698 9898 12703
rect 9870 12651 9898 12670
rect 9926 12642 9954 13006
rect 9926 12609 9954 12614
rect 9918 12558 10050 12563
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 9918 12525 10050 12530
rect 10038 12474 10066 12479
rect 9870 12026 9898 12031
rect 9814 12025 9898 12026
rect 9814 11999 9871 12025
rect 9897 11999 9898 12025
rect 9814 11998 9898 11999
rect 9870 11993 9898 11998
rect 10038 11969 10066 12446
rect 10262 12418 10290 13006
rect 10598 13145 10626 13151
rect 10598 13119 10599 13145
rect 10625 13119 10626 13145
rect 10262 12385 10290 12390
rect 10318 12698 10346 12703
rect 10038 11943 10039 11969
rect 10065 11943 10066 11969
rect 10038 11937 10066 11943
rect 10094 12362 10122 12367
rect 10094 11970 10122 12334
rect 10318 12361 10346 12670
rect 10430 12474 10458 12479
rect 10458 12446 10514 12474
rect 10430 12427 10458 12446
rect 10318 12335 10319 12361
rect 10345 12335 10346 12361
rect 10318 12082 10346 12335
rect 9534 11495 9535 11521
rect 9561 11495 9562 11521
rect 9534 11489 9562 11495
rect 9646 11550 9730 11578
rect 9758 11914 9786 11919
rect 9646 11410 9674 11550
rect 9702 11466 9730 11471
rect 9702 11419 9730 11438
rect 9422 11321 9450 11326
rect 9534 11382 9674 11410
rect 9478 11242 9506 11247
rect 9478 11185 9506 11214
rect 9478 11159 9479 11185
rect 9505 11159 9506 11185
rect 9478 11153 9506 11159
rect 9422 10010 9450 10015
rect 9422 9963 9450 9982
rect 9534 9673 9562 11382
rect 9646 10793 9674 10799
rect 9646 10767 9647 10793
rect 9673 10767 9674 10793
rect 9646 9730 9674 10767
rect 9646 9697 9674 9702
rect 9702 10737 9730 10743
rect 9702 10711 9703 10737
rect 9729 10711 9730 10737
rect 9702 9954 9730 10711
rect 9534 9647 9535 9673
rect 9561 9647 9562 9673
rect 9534 9618 9562 9647
rect 9338 9198 9394 9226
rect 9478 9590 9562 9618
rect 9310 9179 9338 9198
rect 9478 9002 9506 9590
rect 9590 9561 9618 9567
rect 9590 9535 9591 9561
rect 9617 9535 9618 9561
rect 9534 9506 9562 9511
rect 9590 9506 9618 9535
rect 9562 9478 9618 9506
rect 9534 9473 9562 9478
rect 9534 9394 9562 9399
rect 9534 9225 9562 9366
rect 9702 9394 9730 9926
rect 9702 9361 9730 9366
rect 9534 9199 9535 9225
rect 9561 9199 9562 9225
rect 9534 9193 9562 9199
rect 9478 8969 9506 8974
rect 9702 9113 9730 9119
rect 9702 9087 9703 9113
rect 9729 9087 9730 9113
rect 9590 8946 9618 8951
rect 9254 8807 9255 8833
rect 9281 8807 9282 8833
rect 9254 8801 9282 8807
rect 9478 8834 9506 8839
rect 9478 8787 9506 8806
rect 9030 8359 9031 8385
rect 9057 8359 9058 8385
rect 9030 8353 9058 8359
rect 9198 8498 9226 8503
rect 9198 8441 9226 8470
rect 9198 8415 9199 8441
rect 9225 8415 9226 8441
rect 9198 8386 9226 8415
rect 9590 8441 9618 8918
rect 9590 8415 9591 8441
rect 9617 8415 9618 8441
rect 9198 8353 9226 8358
rect 9534 8386 9562 8391
rect 9534 8339 9562 8358
rect 9590 7938 9618 8415
rect 9702 8050 9730 9087
rect 9758 8890 9786 11886
rect 9926 11914 9954 11919
rect 9926 11867 9954 11886
rect 9918 11774 10050 11779
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 9918 11741 10050 11746
rect 10094 11690 10122 11942
rect 10206 12054 10346 12082
rect 10038 11662 10122 11690
rect 10150 11858 10178 11863
rect 10206 11858 10234 12054
rect 10150 11857 10234 11858
rect 10150 11831 10151 11857
rect 10177 11831 10234 11857
rect 10150 11830 10234 11831
rect 10262 11913 10290 11919
rect 10262 11887 10263 11913
rect 10289 11887 10290 11913
rect 9926 11578 9954 11583
rect 9870 11577 9954 11578
rect 9870 11551 9927 11577
rect 9953 11551 9954 11577
rect 9870 11550 9954 11551
rect 9814 11242 9842 11247
rect 9814 11185 9842 11214
rect 9814 11159 9815 11185
rect 9841 11159 9842 11185
rect 9814 11153 9842 11159
rect 9870 11074 9898 11550
rect 9926 11545 9954 11550
rect 9982 11242 10010 11247
rect 9926 11186 9954 11191
rect 9926 11139 9954 11158
rect 9982 11130 10010 11214
rect 10038 11241 10066 11662
rect 10094 11577 10122 11583
rect 10094 11551 10095 11577
rect 10121 11551 10122 11577
rect 10094 11298 10122 11551
rect 10094 11265 10122 11270
rect 10038 11215 10039 11241
rect 10065 11215 10066 11241
rect 10038 11209 10066 11215
rect 10094 11186 10122 11191
rect 10094 11139 10122 11158
rect 9982 11097 10010 11102
rect 9814 11046 9898 11074
rect 9814 9338 9842 11046
rect 10150 11018 10178 11830
rect 10262 11689 10290 11887
rect 10262 11663 10263 11689
rect 10289 11663 10290 11689
rect 10262 11657 10290 11663
rect 10486 11690 10514 12446
rect 10598 12473 10626 13119
rect 10822 13146 10850 13151
rect 10822 12753 10850 13118
rect 11158 13146 11186 13151
rect 11158 13099 11186 13118
rect 11382 13146 11410 13151
rect 11382 13099 11410 13118
rect 11774 13146 11802 13151
rect 11774 13099 11802 13118
rect 11942 13145 11970 13151
rect 11942 13119 11943 13145
rect 11969 13119 11970 13145
rect 10822 12727 10823 12753
rect 10849 12727 10850 12753
rect 10822 12721 10850 12727
rect 11438 12866 11466 12871
rect 10654 12698 10682 12703
rect 10654 12651 10682 12670
rect 10710 12641 10738 12647
rect 10710 12615 10711 12641
rect 10737 12615 10738 12641
rect 10710 12530 10738 12615
rect 10598 12447 10599 12473
rect 10625 12447 10626 12473
rect 10598 12441 10626 12447
rect 10654 12502 10738 12530
rect 10654 12474 10682 12502
rect 10654 12441 10682 12446
rect 11438 12473 11466 12838
rect 11942 12866 11970 13119
rect 11942 12833 11970 12838
rect 12950 13145 12978 13426
rect 12950 13119 12951 13145
rect 12977 13119 12978 13145
rect 11438 12447 11439 12473
rect 11465 12447 11466 12473
rect 11438 12441 11466 12447
rect 10542 12417 10570 12423
rect 10542 12391 10543 12417
rect 10569 12391 10570 12417
rect 10542 12194 10570 12391
rect 10710 12418 10738 12423
rect 10710 12371 10738 12390
rect 10878 12362 10906 12367
rect 10878 12315 10906 12334
rect 11270 12362 11298 12367
rect 11270 12315 11298 12334
rect 12950 12306 12978 13119
rect 13230 12865 13258 13455
rect 14574 13257 14602 13510
rect 18830 13538 18858 13543
rect 18830 13491 18858 13510
rect 14630 13426 14658 13431
rect 14630 13425 14714 13426
rect 14630 13399 14631 13425
rect 14657 13399 14714 13425
rect 14630 13398 14714 13399
rect 14630 13393 14658 13398
rect 14574 13231 14575 13257
rect 14601 13231 14602 13257
rect 14574 13225 14602 13231
rect 14462 13145 14490 13151
rect 14630 13146 14658 13151
rect 14462 13119 14463 13145
rect 14489 13119 14490 13145
rect 13286 13090 13314 13095
rect 13286 13089 13426 13090
rect 13286 13063 13287 13089
rect 13313 13063 13426 13089
rect 13286 13062 13426 13063
rect 13286 13057 13314 13062
rect 13230 12839 13231 12865
rect 13257 12839 13258 12865
rect 13230 12833 13258 12839
rect 13398 12865 13426 13062
rect 14350 13089 14378 13095
rect 14350 13063 14351 13089
rect 14377 13063 14378 13089
rect 13398 12839 13399 12865
rect 13425 12839 13426 12865
rect 13398 12833 13426 12839
rect 14070 12866 14098 12871
rect 13734 12810 13762 12815
rect 13286 12754 13314 12759
rect 13286 12707 13314 12726
rect 13734 12753 13762 12782
rect 13734 12727 13735 12753
rect 13761 12727 13762 12753
rect 13734 12721 13762 12727
rect 14070 12753 14098 12838
rect 14070 12727 14071 12753
rect 14097 12727 14098 12753
rect 14070 12721 14098 12727
rect 13566 12698 13594 12703
rect 13566 12651 13594 12670
rect 13230 12642 13258 12647
rect 13230 12595 13258 12614
rect 13454 12642 13482 12647
rect 13454 12595 13482 12614
rect 13678 12642 13706 12647
rect 13454 12361 13482 12367
rect 13454 12335 13455 12361
rect 13481 12335 13482 12361
rect 12950 12273 12978 12278
rect 13286 12306 13314 12311
rect 13398 12306 13426 12311
rect 13454 12306 13482 12335
rect 13286 12305 13398 12306
rect 13286 12279 13287 12305
rect 13313 12279 13398 12305
rect 13286 12278 13398 12279
rect 13426 12278 13482 12306
rect 10542 12166 10626 12194
rect 10598 11914 10626 12166
rect 12166 11969 12194 11975
rect 12166 11943 12167 11969
rect 12193 11943 12194 11969
rect 10542 11690 10570 11695
rect 10486 11689 10570 11690
rect 10486 11663 10543 11689
rect 10569 11663 10570 11689
rect 10486 11662 10570 11663
rect 10542 11657 10570 11662
rect 10206 11633 10234 11639
rect 10206 11607 10207 11633
rect 10233 11607 10234 11633
rect 10206 11298 10234 11607
rect 10430 11634 10458 11639
rect 10430 11633 10514 11634
rect 10430 11607 10431 11633
rect 10457 11607 10514 11633
rect 10430 11606 10514 11607
rect 10430 11601 10458 11606
rect 10374 11578 10402 11583
rect 10374 11531 10402 11550
rect 10430 11466 10458 11471
rect 10206 11265 10234 11270
rect 10262 11354 10290 11359
rect 10206 11186 10234 11191
rect 10262 11186 10290 11326
rect 10206 11185 10290 11186
rect 10206 11159 10207 11185
rect 10233 11159 10290 11185
rect 10206 11158 10290 11159
rect 10206 11153 10234 11158
rect 10430 11130 10458 11438
rect 10374 11102 10458 11130
rect 10374 11101 10402 11102
rect 9918 10990 10050 10995
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 9918 10957 10050 10962
rect 10094 10990 10178 11018
rect 10318 11073 10346 11079
rect 10318 11047 10319 11073
rect 10345 11047 10346 11073
rect 10374 11075 10375 11101
rect 10401 11075 10402 11101
rect 10374 11069 10402 11075
rect 10318 11018 10346 11047
rect 10318 10990 10402 11018
rect 10094 10906 10122 10990
rect 9926 10878 10122 10906
rect 10262 10906 10290 10911
rect 9926 10737 9954 10878
rect 10038 10794 10066 10799
rect 10206 10794 10234 10799
rect 10262 10794 10290 10878
rect 10038 10793 10122 10794
rect 10038 10767 10039 10793
rect 10065 10767 10122 10793
rect 10038 10766 10122 10767
rect 10038 10761 10066 10766
rect 9926 10711 9927 10737
rect 9953 10711 9954 10737
rect 9926 10705 9954 10711
rect 10038 10402 10066 10407
rect 10038 10355 10066 10374
rect 10094 10290 10122 10766
rect 10094 10257 10122 10262
rect 10206 10793 10290 10794
rect 10206 10767 10207 10793
rect 10233 10767 10290 10793
rect 10206 10766 10290 10767
rect 10318 10849 10346 10855
rect 10318 10823 10319 10849
rect 10345 10823 10346 10849
rect 10318 10794 10346 10823
rect 10374 10850 10402 10990
rect 10430 10850 10458 10855
rect 10374 10849 10458 10850
rect 10374 10823 10431 10849
rect 10457 10823 10458 10849
rect 10374 10822 10458 10823
rect 9918 10206 10050 10211
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 9918 10173 10050 10178
rect 10150 9674 10178 9679
rect 9918 9422 10050 9427
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 9918 9389 10050 9394
rect 9814 9305 9842 9310
rect 9870 9282 9898 9287
rect 9814 9226 9842 9231
rect 9814 9179 9842 9198
rect 9758 8843 9786 8862
rect 9870 8778 9898 9254
rect 9758 8750 9898 8778
rect 9926 8834 9954 8839
rect 9758 8553 9786 8750
rect 9926 8722 9954 8806
rect 9758 8527 9759 8553
rect 9785 8527 9786 8553
rect 9758 8521 9786 8527
rect 9814 8694 9954 8722
rect 10150 8833 10178 9646
rect 10206 9618 10234 10766
rect 10318 10761 10346 10766
rect 10430 10346 10458 10822
rect 10486 10794 10514 11606
rect 10486 10761 10514 10766
rect 10430 10313 10458 10318
rect 10206 9282 10234 9590
rect 10374 9730 10402 9735
rect 10374 9617 10402 9702
rect 10374 9591 10375 9617
rect 10401 9591 10402 9617
rect 10374 9585 10402 9591
rect 10206 9249 10234 9254
rect 10542 9506 10570 9511
rect 10542 9281 10570 9478
rect 10598 9450 10626 11886
rect 11998 11913 12026 11919
rect 11998 11887 11999 11913
rect 12025 11887 12026 11913
rect 11662 11858 11690 11863
rect 10934 11577 10962 11583
rect 10934 11551 10935 11577
rect 10961 11551 10962 11577
rect 10934 11522 10962 11551
rect 10822 11298 10850 11303
rect 10710 11186 10738 11191
rect 10738 11158 10794 11186
rect 10710 11153 10738 11158
rect 10654 11130 10682 11135
rect 10654 11083 10682 11102
rect 10766 10906 10794 11158
rect 10822 11074 10850 11270
rect 10822 11027 10850 11046
rect 10654 10878 10906 10906
rect 10654 9674 10682 10878
rect 10878 10849 10906 10878
rect 10878 10823 10879 10849
rect 10905 10823 10906 10849
rect 10878 10817 10906 10823
rect 10710 10794 10738 10799
rect 10934 10794 10962 11494
rect 11270 11521 11298 11527
rect 11270 11495 11271 11521
rect 11297 11495 11298 11521
rect 10990 11130 11018 11135
rect 10990 10906 11018 11102
rect 11270 11074 11298 11495
rect 11662 11297 11690 11830
rect 11662 11271 11663 11297
rect 11689 11271 11690 11297
rect 11662 11265 11690 11271
rect 11830 11410 11858 11415
rect 11550 11185 11578 11191
rect 11550 11159 11551 11185
rect 11577 11159 11578 11185
rect 11494 11074 11522 11079
rect 11270 11073 11522 11074
rect 11270 11047 11495 11073
rect 11521 11047 11522 11073
rect 11270 11046 11522 11047
rect 11494 11041 11522 11046
rect 11214 10906 11242 10911
rect 10990 10905 11242 10906
rect 10990 10879 10991 10905
rect 11017 10879 11215 10905
rect 11241 10879 11242 10905
rect 10990 10878 11242 10879
rect 10990 10873 11018 10878
rect 11214 10873 11242 10878
rect 11046 10794 11074 10799
rect 10934 10766 11018 10794
rect 10710 10345 10738 10766
rect 10710 10319 10711 10345
rect 10737 10319 10738 10345
rect 10710 10313 10738 10319
rect 10766 10737 10794 10743
rect 10766 10711 10767 10737
rect 10793 10711 10794 10737
rect 10654 9641 10682 9646
rect 10598 9422 10682 9450
rect 10542 9255 10543 9281
rect 10569 9255 10570 9281
rect 10542 9249 10570 9255
rect 10598 9338 10626 9343
rect 10150 8807 10151 8833
rect 10177 8807 10178 8833
rect 9814 8106 9842 8694
rect 9918 8638 10050 8643
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 9918 8605 10050 8610
rect 10094 8442 10122 8447
rect 10150 8442 10178 8807
rect 10598 8833 10626 9310
rect 10654 9170 10682 9422
rect 10766 9282 10794 10711
rect 10878 10458 10906 10463
rect 10878 10411 10906 10430
rect 10934 10345 10962 10351
rect 10934 10319 10935 10345
rect 10961 10319 10962 10345
rect 10822 10290 10850 10295
rect 10850 10262 10906 10290
rect 10822 10243 10850 10262
rect 10766 9249 10794 9254
rect 10822 10066 10850 10071
rect 10654 9137 10682 9142
rect 10822 8834 10850 10038
rect 10598 8807 10599 8833
rect 10625 8807 10626 8833
rect 10598 8801 10626 8807
rect 10710 8833 10850 8834
rect 10710 8807 10823 8833
rect 10849 8807 10850 8833
rect 10710 8806 10850 8807
rect 10206 8778 10234 8783
rect 10234 8750 10290 8778
rect 10206 8745 10234 8750
rect 10094 8441 10178 8442
rect 10094 8415 10095 8441
rect 10121 8415 10178 8441
rect 10094 8414 10178 8415
rect 10262 8498 10290 8750
rect 10094 8409 10122 8414
rect 10206 8330 10234 8335
rect 9982 8106 10010 8111
rect 9814 8105 10010 8106
rect 9814 8079 9983 8105
rect 10009 8079 10010 8105
rect 9814 8078 10010 8079
rect 9982 8073 10010 8078
rect 9702 8017 9730 8022
rect 10206 8049 10234 8302
rect 10206 8023 10207 8049
rect 10233 8023 10234 8049
rect 8750 7574 8890 7602
rect 8862 7546 8890 7574
rect 8862 7513 8890 7518
rect 9030 7601 9058 7607
rect 9030 7575 9031 7601
rect 9057 7575 9058 7601
rect 8582 7321 8666 7322
rect 8582 7295 8583 7321
rect 8609 7295 8666 7321
rect 8582 7294 8666 7295
rect 8862 7322 8890 7327
rect 8582 7289 8610 7294
rect 8414 6929 8498 6930
rect 8414 6903 8415 6929
rect 8441 6903 8498 6929
rect 8414 6902 8498 6903
rect 8414 6897 8442 6902
rect 8358 6561 8386 6566
rect 7630 6511 7631 6537
rect 7657 6511 7658 6537
rect 7630 6505 7658 6511
rect 8694 6537 8722 6543
rect 8694 6511 8695 6537
rect 8721 6511 8722 6537
rect 7294 6455 7295 6481
rect 7321 6455 7322 6481
rect 7294 6449 7322 6455
rect 8694 6090 8722 6511
rect 8862 6201 8890 7294
rect 9030 7322 9058 7575
rect 9590 7574 9618 7910
rect 10206 7938 10234 8023
rect 10206 7905 10234 7910
rect 9918 7854 10050 7859
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 10262 7826 10290 8470
rect 10318 8777 10346 8783
rect 10318 8751 10319 8777
rect 10345 8751 10346 8777
rect 10318 8442 10346 8751
rect 10374 8721 10402 8727
rect 10374 8695 10375 8721
rect 10401 8695 10402 8721
rect 10374 8554 10402 8695
rect 10542 8554 10570 8559
rect 10374 8553 10570 8554
rect 10374 8527 10375 8553
rect 10401 8527 10543 8553
rect 10569 8527 10570 8553
rect 10374 8526 10570 8527
rect 10374 8521 10402 8526
rect 10542 8521 10570 8526
rect 10710 8553 10738 8806
rect 10822 8801 10850 8806
rect 10878 9114 10906 10262
rect 10934 10066 10962 10319
rect 10934 10033 10962 10038
rect 10990 10010 11018 10766
rect 11046 10737 11074 10766
rect 11046 10711 11047 10737
rect 11073 10711 11074 10737
rect 11046 10705 11074 10711
rect 11326 10793 11354 10799
rect 11326 10767 11327 10793
rect 11353 10767 11354 10793
rect 11270 10402 11298 10407
rect 11270 10065 11298 10374
rect 11326 10122 11354 10767
rect 11326 10089 11354 10094
rect 11270 10039 11271 10065
rect 11297 10039 11298 10065
rect 11270 10033 11298 10039
rect 11550 10066 11578 11159
rect 11774 11130 11802 11135
rect 11774 11083 11802 11102
rect 11662 10794 11690 10799
rect 11662 10747 11690 10766
rect 11830 10738 11858 11382
rect 11886 11354 11914 11359
rect 11886 11186 11914 11326
rect 11886 11185 11970 11186
rect 11886 11159 11887 11185
rect 11913 11159 11970 11185
rect 11886 11158 11970 11159
rect 11886 11153 11914 11158
rect 11942 10962 11970 11158
rect 11998 11130 12026 11887
rect 12054 11858 12082 11863
rect 12054 11811 12082 11830
rect 12166 11522 12194 11943
rect 12334 11522 12362 11527
rect 12166 11521 12362 11522
rect 12166 11495 12335 11521
rect 12361 11495 12362 11521
rect 12166 11494 12362 11495
rect 12334 11466 12362 11494
rect 12670 11522 12698 11527
rect 12670 11475 12698 11494
rect 13286 11522 13314 12278
rect 13398 12259 13426 12278
rect 13286 11489 13314 11494
rect 13678 11857 13706 12614
rect 13902 12641 13930 12647
rect 13902 12615 13903 12641
rect 13929 12615 13930 12641
rect 13846 12305 13874 12311
rect 13846 12279 13847 12305
rect 13873 12279 13874 12305
rect 13846 12081 13874 12279
rect 13846 12055 13847 12081
rect 13873 12055 13874 12081
rect 13846 12049 13874 12055
rect 13902 11969 13930 12615
rect 14014 12641 14042 12647
rect 14014 12615 14015 12641
rect 14041 12615 14042 12641
rect 14014 12418 14042 12615
rect 14350 12642 14378 13063
rect 14462 12754 14490 13119
rect 14462 12721 14490 12726
rect 14574 13145 14658 13146
rect 14574 13119 14631 13145
rect 14657 13119 14658 13145
rect 14574 13118 14658 13119
rect 14574 12866 14602 13118
rect 14630 13113 14658 13118
rect 14686 13090 14714 13398
rect 18942 13145 18970 13151
rect 18942 13119 18943 13145
rect 18969 13119 18970 13145
rect 14854 13090 14882 13095
rect 14686 13089 14882 13090
rect 14686 13063 14855 13089
rect 14881 13063 14882 13089
rect 14686 13062 14882 13063
rect 14574 12753 14602 12838
rect 14630 12865 14658 12871
rect 14630 12839 14631 12865
rect 14657 12839 14658 12865
rect 14630 12810 14658 12839
rect 14630 12777 14658 12782
rect 14574 12727 14575 12753
rect 14601 12727 14602 12753
rect 14574 12721 14602 12727
rect 14350 12609 14378 12614
rect 14630 12642 14658 12647
rect 14630 12595 14658 12614
rect 14014 12385 14042 12390
rect 14630 12306 14658 12311
rect 14686 12306 14714 13062
rect 14854 13057 14882 13062
rect 17598 12950 17730 12955
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17598 12917 17730 12922
rect 18830 12753 18858 12759
rect 18830 12727 18831 12753
rect 18857 12727 18858 12753
rect 18830 12474 18858 12727
rect 18942 12642 18970 13119
rect 20006 13146 20034 13567
rect 20006 13113 20034 13118
rect 19950 13089 19978 13095
rect 19950 13063 19951 13089
rect 19977 13063 19978 13089
rect 19950 12810 19978 13063
rect 19950 12777 19978 12782
rect 20006 12809 20034 12815
rect 20006 12783 20007 12809
rect 20033 12783 20034 12809
rect 18942 12609 18970 12614
rect 18830 12441 18858 12446
rect 20006 12474 20034 12783
rect 20006 12441 20034 12446
rect 14658 12278 14714 12306
rect 14910 12418 14938 12423
rect 15078 12418 15106 12423
rect 14938 12417 15106 12418
rect 14938 12391 15079 12417
rect 15105 12391 15106 12417
rect 14938 12390 15106 12391
rect 14910 12305 14938 12390
rect 15078 12385 15106 12390
rect 15246 12418 15274 12423
rect 15246 12371 15274 12390
rect 18830 12362 18858 12367
rect 18830 12315 18858 12334
rect 14910 12279 14911 12305
rect 14937 12279 14938 12305
rect 14630 12273 14658 12278
rect 14910 12273 14938 12279
rect 20006 12249 20034 12255
rect 20006 12223 20007 12249
rect 20033 12223 20034 12249
rect 17598 12166 17730 12171
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17598 12133 17730 12138
rect 20006 12138 20034 12223
rect 20006 12105 20034 12110
rect 13902 11943 13903 11969
rect 13929 11943 13930 11969
rect 13902 11937 13930 11943
rect 13678 11831 13679 11857
rect 13705 11831 13706 11857
rect 12334 11433 12362 11438
rect 11998 11097 12026 11102
rect 12726 11130 12754 11135
rect 11942 10934 12026 10962
rect 11774 10737 11858 10738
rect 11774 10711 11831 10737
rect 11857 10711 11858 10737
rect 11774 10710 11858 10711
rect 11578 10038 11690 10066
rect 11550 10033 11578 10038
rect 11438 10010 11466 10015
rect 10990 9982 11074 10010
rect 10990 9674 11018 9679
rect 10934 9562 10962 9567
rect 10934 9515 10962 9534
rect 10990 9281 11018 9646
rect 11046 9394 11074 9982
rect 11438 9562 11466 9982
rect 11662 9617 11690 10038
rect 11662 9591 11663 9617
rect 11689 9591 11690 9617
rect 11662 9585 11690 9591
rect 11046 9361 11074 9366
rect 11102 9505 11130 9511
rect 11102 9479 11103 9505
rect 11129 9479 11130 9505
rect 10990 9255 10991 9281
rect 11017 9255 11018 9281
rect 10990 9249 11018 9255
rect 10878 8834 10906 9086
rect 11102 9225 11130 9479
rect 11102 9199 11103 9225
rect 11129 9199 11130 9225
rect 10934 8834 10962 8839
rect 10878 8833 10962 8834
rect 10878 8807 10935 8833
rect 10961 8807 10962 8833
rect 10878 8806 10962 8807
rect 10710 8527 10711 8553
rect 10737 8527 10738 8553
rect 10710 8521 10738 8527
rect 10766 8721 10794 8727
rect 10766 8695 10767 8721
rect 10793 8695 10794 8721
rect 10318 8409 10346 8414
rect 9918 7821 10050 7826
rect 10094 7798 10290 7826
rect 10598 8050 10626 8055
rect 10766 8050 10794 8695
rect 10878 8553 10906 8806
rect 10934 8801 10962 8806
rect 11102 8834 11130 9199
rect 11102 8787 11130 8806
rect 11270 9338 11298 9343
rect 10878 8527 10879 8553
rect 10905 8527 10906 8553
rect 10878 8521 10906 8527
rect 11270 8777 11298 9310
rect 11382 9114 11410 9119
rect 11382 9067 11410 9086
rect 11270 8751 11271 8777
rect 11297 8751 11298 8777
rect 11270 8554 11298 8751
rect 11270 8521 11298 8526
rect 11382 8498 11410 8503
rect 11382 8451 11410 8470
rect 10990 8441 11018 8447
rect 10990 8415 10991 8441
rect 11017 8415 11018 8441
rect 10990 8330 11018 8415
rect 10990 8297 11018 8302
rect 10094 7657 10122 7798
rect 10094 7631 10095 7657
rect 10121 7631 10122 7657
rect 10094 7625 10122 7631
rect 10318 7657 10346 7663
rect 10318 7631 10319 7657
rect 10345 7631 10346 7657
rect 9870 7602 9898 7607
rect 9590 7546 9674 7574
rect 9030 7289 9058 7294
rect 9646 7321 9674 7546
rect 9646 7295 9647 7321
rect 9673 7295 9674 7321
rect 9646 7289 9674 7295
rect 9814 7546 9842 7551
rect 9814 7321 9842 7518
rect 9870 7377 9898 7574
rect 10206 7602 10234 7621
rect 10206 7569 10234 7574
rect 10318 7602 10346 7631
rect 10318 7569 10346 7574
rect 9870 7351 9871 7377
rect 9897 7351 9898 7377
rect 9870 7345 9898 7351
rect 10038 7545 10066 7551
rect 10038 7519 10039 7545
rect 10065 7519 10066 7545
rect 9814 7295 9815 7321
rect 9841 7295 9842 7321
rect 9814 7289 9842 7295
rect 10038 7154 10066 7519
rect 10598 7546 10626 8022
rect 10710 8049 10794 8050
rect 10710 8023 10767 8049
rect 10793 8023 10794 8049
rect 10710 8022 10794 8023
rect 10710 7826 10738 8022
rect 10766 8017 10794 8022
rect 10990 8050 11018 8055
rect 10654 7798 10738 7826
rect 10878 7994 10906 7999
rect 10878 7937 10906 7966
rect 10878 7911 10879 7937
rect 10905 7911 10906 7937
rect 10654 7657 10682 7798
rect 10878 7770 10906 7911
rect 10934 7938 10962 7943
rect 10934 7891 10962 7910
rect 10766 7742 10906 7770
rect 10654 7631 10655 7657
rect 10681 7631 10682 7657
rect 10654 7625 10682 7631
rect 10710 7658 10738 7663
rect 10766 7658 10794 7742
rect 10710 7657 10794 7658
rect 10710 7631 10711 7657
rect 10737 7631 10794 7657
rect 10710 7630 10794 7631
rect 10822 7657 10850 7663
rect 10822 7631 10823 7657
rect 10849 7631 10850 7657
rect 10710 7625 10738 7630
rect 10598 7518 10738 7546
rect 10094 7322 10122 7327
rect 10094 7275 10122 7294
rect 10710 7209 10738 7518
rect 10710 7183 10711 7209
rect 10737 7183 10738 7209
rect 10710 7177 10738 7183
rect 10766 7209 10794 7215
rect 10766 7183 10767 7209
rect 10793 7183 10794 7209
rect 10598 7154 10626 7159
rect 10038 7126 10122 7154
rect 9918 7070 10050 7075
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 9918 7037 10050 7042
rect 10094 6929 10122 7126
rect 10094 6903 10095 6929
rect 10121 6903 10122 6929
rect 10094 6897 10122 6903
rect 10150 7153 10626 7154
rect 10150 7127 10599 7153
rect 10625 7127 10626 7153
rect 10150 7126 10626 7127
rect 9758 6873 9786 6879
rect 9758 6847 9759 6873
rect 9785 6847 9786 6873
rect 9758 6762 9786 6847
rect 8918 6594 8946 6599
rect 8918 6547 8946 6566
rect 9198 6538 9226 6543
rect 8974 6510 9198 6538
rect 8974 6481 9002 6510
rect 9198 6491 9226 6510
rect 8974 6455 8975 6481
rect 9001 6455 9002 6481
rect 8974 6449 9002 6455
rect 8862 6175 8863 6201
rect 8889 6175 8890 6201
rect 8862 6169 8890 6175
rect 8918 6369 8946 6375
rect 8918 6343 8919 6369
rect 8945 6343 8946 6369
rect 8918 6090 8946 6343
rect 8694 6062 8946 6090
rect 9758 6089 9786 6734
rect 9918 6286 10050 6291
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 9918 6253 10050 6258
rect 10150 6145 10178 7126
rect 10598 7121 10626 7126
rect 10150 6119 10151 6145
rect 10177 6119 10178 6145
rect 10150 6113 10178 6119
rect 10710 6818 10738 6823
rect 9758 6063 9759 6089
rect 9785 6063 9786 6089
rect 2238 5894 2370 5899
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2238 5861 2370 5866
rect 2238 5110 2370 5115
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2238 5077 2370 5082
rect 2238 4326 2370 4331
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2238 4293 2370 4298
rect 8694 4214 8722 6062
rect 9758 6057 9786 6063
rect 9918 5502 10050 5507
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 9918 5469 10050 5474
rect 9918 4718 10050 4723
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 9918 4685 10050 4690
rect 8526 4186 8722 4214
rect 2238 3542 2370 3547
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2238 3509 2370 3514
rect 2238 2758 2370 2763
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2238 2725 2370 2730
rect 2238 1974 2370 1979
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2238 1941 2370 1946
rect 8526 1777 8554 4186
rect 9918 3934 10050 3939
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 9918 3901 10050 3906
rect 9918 3150 10050 3155
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 9918 3117 10050 3122
rect 9918 2366 10050 2371
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 9918 2333 10050 2338
rect 8526 1751 8527 1777
rect 8553 1751 8554 1777
rect 8526 1745 8554 1751
rect 10710 1777 10738 6790
rect 10766 6593 10794 7183
rect 10822 6818 10850 7631
rect 10934 7658 10962 7663
rect 10990 7658 11018 8022
rect 11438 8050 11466 9534
rect 11550 9506 11578 9511
rect 11550 9459 11578 9478
rect 11606 9505 11634 9511
rect 11606 9479 11607 9505
rect 11633 9479 11634 9505
rect 11550 9394 11578 9399
rect 11550 8834 11578 9366
rect 11606 9282 11634 9479
rect 11718 9282 11746 9287
rect 11606 9281 11746 9282
rect 11606 9255 11719 9281
rect 11745 9255 11746 9281
rect 11606 9254 11746 9255
rect 11718 9249 11746 9254
rect 11550 8833 11634 8834
rect 11550 8807 11551 8833
rect 11577 8807 11634 8833
rect 11550 8806 11634 8807
rect 11550 8801 11578 8806
rect 11550 8497 11578 8503
rect 11550 8471 11551 8497
rect 11577 8471 11578 8497
rect 11550 8386 11578 8471
rect 11550 8353 11578 8358
rect 11438 8017 11466 8022
rect 10934 7657 11018 7658
rect 10934 7631 10935 7657
rect 10961 7631 11018 7657
rect 10934 7630 11018 7631
rect 10934 7625 10962 7630
rect 10878 7602 10906 7621
rect 10878 7569 10906 7574
rect 11606 7266 11634 8806
rect 11662 7266 11690 7271
rect 11606 7265 11690 7266
rect 11606 7239 11663 7265
rect 11689 7239 11690 7265
rect 11606 7238 11690 7239
rect 10822 6785 10850 6790
rect 11158 6818 11186 6823
rect 11158 6771 11186 6790
rect 11382 6817 11410 6823
rect 11382 6791 11383 6817
rect 11409 6791 11410 6817
rect 10766 6567 10767 6593
rect 10793 6567 10794 6593
rect 10766 6561 10794 6567
rect 11382 6762 11410 6791
rect 10822 6538 10850 6543
rect 10822 6481 10850 6510
rect 11046 6538 11074 6543
rect 11046 6491 11074 6510
rect 10822 6455 10823 6481
rect 10849 6455 10850 6481
rect 10822 6449 10850 6455
rect 11382 6482 11410 6734
rect 10766 6369 10794 6375
rect 10766 6343 10767 6369
rect 10793 6343 10794 6369
rect 10766 6034 10794 6343
rect 11382 6202 11410 6454
rect 11662 6482 11690 7238
rect 11774 7210 11802 10710
rect 11830 10705 11858 10710
rect 11886 9730 11914 9735
rect 11830 9617 11858 9623
rect 11830 9591 11831 9617
rect 11857 9591 11858 9617
rect 11830 9394 11858 9591
rect 11830 9361 11858 9366
rect 11830 9282 11858 9287
rect 11886 9282 11914 9702
rect 11858 9254 11914 9282
rect 11942 9281 11970 9287
rect 11942 9255 11943 9281
rect 11969 9255 11970 9281
rect 11830 9235 11858 9254
rect 11886 9169 11914 9175
rect 11886 9143 11887 9169
rect 11913 9143 11914 9169
rect 11830 9114 11858 9119
rect 11830 7574 11858 9086
rect 11886 8889 11914 9143
rect 11886 8863 11887 8889
rect 11913 8863 11914 8889
rect 11886 8857 11914 8863
rect 11942 8946 11970 9255
rect 11998 9225 12026 10934
rect 12726 10905 12754 11102
rect 13118 11130 13146 11135
rect 13118 11083 13146 11102
rect 13678 11130 13706 11831
rect 13678 11097 13706 11102
rect 13790 11857 13818 11863
rect 13790 11831 13791 11857
rect 13817 11831 13818 11857
rect 12950 11074 12978 11079
rect 12726 10879 12727 10905
rect 12753 10879 12754 10905
rect 12726 10873 12754 10879
rect 12782 11073 12978 11074
rect 12782 11047 12951 11073
rect 12977 11047 12978 11073
rect 12782 11046 12978 11047
rect 12614 10793 12642 10799
rect 12614 10767 12615 10793
rect 12641 10767 12642 10793
rect 12054 10738 12082 10743
rect 12054 10691 12082 10710
rect 12222 10738 12250 10743
rect 12110 10682 12138 10687
rect 12110 10635 12138 10654
rect 12222 9673 12250 10710
rect 12614 10682 12642 10767
rect 12670 10738 12698 10743
rect 12670 10691 12698 10710
rect 12614 10402 12642 10654
rect 12614 10369 12642 10374
rect 12670 10458 12698 10463
rect 12782 10458 12810 11046
rect 12950 11041 12978 11046
rect 12698 10430 12810 10458
rect 12950 10793 12978 10799
rect 12950 10767 12951 10793
rect 12977 10767 12978 10793
rect 12670 10009 12698 10430
rect 12950 10121 12978 10767
rect 13622 10793 13650 10799
rect 13622 10767 13623 10793
rect 13649 10767 13650 10793
rect 13454 10738 13482 10743
rect 13622 10738 13650 10767
rect 13454 10737 13650 10738
rect 13454 10711 13455 10737
rect 13481 10711 13650 10737
rect 13454 10710 13650 10711
rect 13454 10457 13482 10710
rect 13454 10431 13455 10457
rect 13481 10431 13482 10457
rect 13454 10425 13482 10431
rect 12950 10095 12951 10121
rect 12977 10095 12978 10121
rect 12950 10089 12978 10095
rect 12670 9983 12671 10009
rect 12697 9983 12698 10009
rect 12670 9977 12698 9983
rect 12726 10009 12754 10015
rect 12726 9983 12727 10009
rect 12753 9983 12754 10009
rect 12222 9647 12223 9673
rect 12249 9647 12250 9673
rect 12222 9641 12250 9647
rect 11998 9199 11999 9225
rect 12025 9199 12026 9225
rect 11998 9193 12026 9199
rect 12726 9114 12754 9983
rect 12838 10010 12866 10015
rect 12838 9963 12866 9982
rect 12950 10009 12978 10015
rect 12950 9983 12951 10009
rect 12977 9983 12978 10009
rect 12950 9674 12978 9983
rect 13622 10009 13650 10710
rect 13622 9983 13623 10009
rect 13649 9983 13650 10009
rect 13454 9954 13482 9959
rect 13622 9954 13650 9983
rect 13454 9953 13650 9954
rect 13454 9927 13455 9953
rect 13481 9927 13650 9953
rect 13454 9926 13650 9927
rect 12950 9641 12978 9646
rect 13286 9674 13314 9679
rect 13286 9627 13314 9646
rect 12726 9081 12754 9086
rect 12950 9506 12978 9511
rect 13454 9506 13482 9926
rect 13566 9730 13594 9735
rect 13790 9730 13818 11831
rect 13958 11690 13986 11695
rect 13958 11185 13986 11662
rect 18830 11578 18858 11583
rect 18830 11531 18858 11550
rect 20006 11466 20034 11471
rect 20006 11419 20034 11438
rect 17598 11382 17730 11387
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17598 11349 17730 11354
rect 20006 11241 20034 11247
rect 20006 11215 20007 11241
rect 20033 11215 20034 11241
rect 13958 11159 13959 11185
rect 13985 11159 13986 11185
rect 13958 11153 13986 11159
rect 14126 11186 14154 11191
rect 14126 11139 14154 11158
rect 14518 11186 14546 11191
rect 14518 11139 14546 11158
rect 18830 11186 18858 11191
rect 18830 11139 18858 11158
rect 13846 11130 13874 11135
rect 13846 11083 13874 11102
rect 14686 11129 14714 11135
rect 14686 11103 14687 11129
rect 14713 11103 14714 11129
rect 13902 11073 13930 11079
rect 13902 11047 13903 11073
rect 13929 11047 13930 11073
rect 13902 10850 13930 11047
rect 14630 11074 14658 11079
rect 14630 11027 14658 11046
rect 14014 10850 14042 10855
rect 13902 10849 14042 10850
rect 13902 10823 14015 10849
rect 14041 10823 14042 10849
rect 13902 10822 14042 10823
rect 14014 10817 14042 10822
rect 14686 10794 14714 11103
rect 20006 11130 20034 11215
rect 20006 11097 20034 11102
rect 14574 10402 14602 10407
rect 14574 10355 14602 10374
rect 14686 10402 14714 10766
rect 15078 11074 15106 11079
rect 15078 10737 15106 11046
rect 15078 10711 15079 10737
rect 15105 10711 15106 10737
rect 15078 10705 15106 10711
rect 18942 10793 18970 10799
rect 18942 10767 18943 10793
rect 18969 10767 18970 10793
rect 17598 10598 17730 10603
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17598 10565 17730 10570
rect 15078 10514 15106 10519
rect 14686 10369 14714 10374
rect 14910 10513 15106 10514
rect 14910 10487 15079 10513
rect 15105 10487 15106 10513
rect 14910 10486 15106 10487
rect 14910 10401 14938 10486
rect 15078 10481 15106 10486
rect 14910 10375 14911 10401
rect 14937 10375 14938 10401
rect 14910 10369 14938 10375
rect 15022 10402 15050 10407
rect 15022 10355 15050 10374
rect 18830 10401 18858 10407
rect 18830 10375 18831 10401
rect 18857 10375 18858 10401
rect 14014 10290 14042 10295
rect 14014 10065 14042 10262
rect 14630 10290 14658 10295
rect 14630 10243 14658 10262
rect 14686 10289 14714 10295
rect 14686 10263 14687 10289
rect 14713 10263 14714 10289
rect 14014 10039 14015 10065
rect 14041 10039 14042 10065
rect 14014 10033 14042 10039
rect 13594 9702 13650 9730
rect 13566 9697 13594 9702
rect 13510 9506 13538 9511
rect 13454 9505 13538 9506
rect 13454 9479 13511 9505
rect 13537 9479 13538 9505
rect 13454 9478 13538 9479
rect 11942 8386 11970 8918
rect 12950 8890 12978 9478
rect 13398 9226 13426 9231
rect 13510 9226 13538 9478
rect 13342 9225 13538 9226
rect 13342 9199 13399 9225
rect 13425 9199 13538 9225
rect 13342 9198 13538 9199
rect 12950 8843 12978 8862
rect 13230 9170 13258 9175
rect 13342 9170 13370 9198
rect 13398 9179 13426 9198
rect 13230 9169 13370 9170
rect 13230 9143 13231 9169
rect 13257 9143 13370 9169
rect 13230 9142 13370 9143
rect 13062 8442 13090 8447
rect 13230 8442 13258 9142
rect 13342 8946 13370 8951
rect 13342 8833 13370 8918
rect 13510 8890 13538 8895
rect 13510 8889 13594 8890
rect 13510 8863 13511 8889
rect 13537 8863 13594 8889
rect 13510 8862 13594 8863
rect 13510 8857 13538 8862
rect 13342 8807 13343 8833
rect 13369 8807 13370 8833
rect 13342 8801 13370 8807
rect 13454 8833 13482 8839
rect 13454 8807 13455 8833
rect 13481 8807 13482 8833
rect 13454 8778 13482 8807
rect 13510 8778 13538 8783
rect 13454 8750 13510 8778
rect 13510 8745 13538 8750
rect 13566 8722 13594 8862
rect 13622 8833 13650 9702
rect 13790 9697 13818 9702
rect 14238 9562 14266 9567
rect 14294 9562 14322 9567
rect 14238 9561 14294 9562
rect 14238 9535 14239 9561
rect 14265 9535 14294 9561
rect 14238 9534 14294 9535
rect 14238 9529 14266 9534
rect 14070 9505 14098 9511
rect 14070 9479 14071 9505
rect 14097 9479 14098 9505
rect 13790 9169 13818 9175
rect 13790 9143 13791 9169
rect 13817 9143 13818 9169
rect 13622 8807 13623 8833
rect 13649 8807 13650 8833
rect 13622 8801 13650 8807
rect 13734 8946 13762 8951
rect 13734 8833 13762 8918
rect 13734 8807 13735 8833
rect 13761 8807 13762 8833
rect 13734 8801 13762 8807
rect 13790 8722 13818 9143
rect 13846 9002 13874 9007
rect 13874 8974 13930 9002
rect 13846 8969 13874 8974
rect 13902 8833 13930 8974
rect 13902 8807 13903 8833
rect 13929 8807 13930 8833
rect 13902 8801 13930 8807
rect 14070 8833 14098 9479
rect 14182 9506 14210 9511
rect 14182 9459 14210 9478
rect 14294 9282 14322 9534
rect 14686 9562 14714 10263
rect 15078 10289 15106 10295
rect 15078 10263 15079 10289
rect 15105 10263 15106 10289
rect 15078 10122 15106 10263
rect 15078 9953 15106 10094
rect 18830 10122 18858 10375
rect 18830 10089 18858 10094
rect 15078 9927 15079 9953
rect 15105 9927 15106 9953
rect 15078 9921 15106 9927
rect 17598 9814 17730 9819
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17598 9781 17730 9786
rect 18942 9674 18970 10767
rect 19950 10737 19978 10743
rect 19950 10711 19951 10737
rect 19977 10711 19978 10737
rect 19950 10458 19978 10711
rect 19950 10425 19978 10430
rect 20006 10457 20034 10463
rect 20006 10431 20007 10457
rect 20033 10431 20034 10457
rect 20006 10122 20034 10431
rect 20006 10089 20034 10094
rect 18942 9641 18970 9646
rect 14686 9529 14714 9534
rect 14070 8807 14071 8833
rect 14097 8807 14098 8833
rect 14070 8801 14098 8807
rect 14238 9170 14266 9175
rect 14126 8778 14154 8783
rect 14126 8731 14154 8750
rect 14238 8777 14266 9142
rect 14294 8833 14322 9254
rect 14910 9506 14938 9511
rect 14854 9170 14882 9175
rect 14854 9123 14882 9142
rect 14294 8807 14295 8833
rect 14321 8807 14322 8833
rect 14294 8801 14322 8807
rect 14910 8834 14938 9478
rect 18830 9225 18858 9231
rect 18830 9199 18831 9225
rect 18857 9199 18858 9225
rect 17598 9030 17730 9035
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17598 8997 17730 9002
rect 18830 8946 18858 9199
rect 18830 8913 18858 8918
rect 18942 9170 18970 9175
rect 14238 8751 14239 8777
rect 14265 8751 14266 8777
rect 14238 8745 14266 8751
rect 13566 8694 13818 8722
rect 13902 8721 13930 8727
rect 13902 8695 13903 8721
rect 13929 8695 13930 8721
rect 13846 8498 13874 8503
rect 13902 8498 13930 8695
rect 13846 8497 13930 8498
rect 13846 8471 13847 8497
rect 13873 8471 13930 8497
rect 13846 8470 13930 8471
rect 13846 8465 13874 8470
rect 13286 8442 13314 8447
rect 13454 8442 13482 8447
rect 13062 8441 13482 8442
rect 13062 8415 13063 8441
rect 13089 8415 13287 8441
rect 13313 8415 13455 8441
rect 13481 8415 13482 8441
rect 13062 8414 13482 8415
rect 13062 8409 13090 8414
rect 11886 7938 11914 7943
rect 11886 7657 11914 7910
rect 11942 7714 11970 8358
rect 12502 8050 12530 8055
rect 12502 8003 12530 8022
rect 12334 7938 12362 7943
rect 11942 7681 11970 7686
rect 12110 7937 12362 7938
rect 12110 7911 12335 7937
rect 12361 7911 12362 7937
rect 12110 7910 12362 7911
rect 12110 7713 12138 7910
rect 12334 7905 12362 7910
rect 12446 7938 12474 7943
rect 12446 7891 12474 7910
rect 13118 7938 13146 7943
rect 12110 7687 12111 7713
rect 12137 7687 12138 7713
rect 12110 7681 12138 7687
rect 12166 7714 12194 7719
rect 11886 7631 11887 7657
rect 11913 7631 11914 7657
rect 11886 7625 11914 7631
rect 11998 7658 12026 7663
rect 11998 7657 12082 7658
rect 11998 7631 11999 7657
rect 12025 7631 12082 7657
rect 11998 7630 12082 7631
rect 11998 7625 12026 7630
rect 11830 7546 12026 7574
rect 11774 7182 11970 7210
rect 11942 6930 11970 7182
rect 11998 6986 12026 7546
rect 12054 7321 12082 7630
rect 12166 7657 12194 7686
rect 12166 7631 12167 7657
rect 12193 7631 12194 7657
rect 12166 7625 12194 7631
rect 12054 7295 12055 7321
rect 12081 7295 12082 7321
rect 12054 7289 12082 7295
rect 13118 7321 13146 7910
rect 13118 7295 13119 7321
rect 13145 7295 13146 7321
rect 12222 6986 12250 6991
rect 12894 6986 12922 6991
rect 11998 6985 12250 6986
rect 11998 6959 12223 6985
rect 12249 6959 12250 6985
rect 11998 6958 12250 6959
rect 12222 6953 12250 6958
rect 12726 6985 12922 6986
rect 12726 6959 12895 6985
rect 12921 6959 12922 6985
rect 12726 6958 12922 6959
rect 11942 6874 11970 6902
rect 12614 6930 12642 6935
rect 12614 6883 12642 6902
rect 12670 6930 12698 6935
rect 12726 6930 12754 6958
rect 12670 6929 12754 6930
rect 12670 6903 12671 6929
rect 12697 6903 12754 6929
rect 12670 6902 12754 6903
rect 11998 6874 12026 6879
rect 11942 6873 12026 6874
rect 11942 6847 11999 6873
rect 12025 6847 12026 6873
rect 11942 6846 12026 6847
rect 11942 6538 11970 6846
rect 11998 6841 12026 6846
rect 12278 6874 12306 6879
rect 12278 6827 12306 6846
rect 11942 6505 11970 6510
rect 12222 6761 12250 6767
rect 12222 6735 12223 6761
rect 12249 6735 12250 6761
rect 12222 6537 12250 6735
rect 12222 6511 12223 6537
rect 12249 6511 12250 6537
rect 12222 6505 12250 6511
rect 11662 6449 11690 6454
rect 11830 6482 11858 6487
rect 11830 6435 11858 6454
rect 11438 6202 11466 6207
rect 11382 6201 11466 6202
rect 11382 6175 11439 6201
rect 11465 6175 11466 6201
rect 11382 6174 11466 6175
rect 11438 6169 11466 6174
rect 10766 6001 10794 6006
rect 11214 6034 11242 6039
rect 11214 4214 11242 6006
rect 12670 4214 12698 6902
rect 12782 6874 12810 6879
rect 12782 6827 12810 6846
rect 12894 6874 12922 6958
rect 13062 6930 13090 6935
rect 13062 6883 13090 6902
rect 12894 6841 12922 6846
rect 13118 6650 13146 7295
rect 13286 7154 13314 8414
rect 13454 8409 13482 8414
rect 14910 8385 14938 8806
rect 18830 8834 18858 8839
rect 18830 8787 18858 8806
rect 18942 8441 18970 9142
rect 20006 9114 20034 9119
rect 20006 9067 20034 9086
rect 20006 8889 20034 8895
rect 20006 8863 20007 8889
rect 20033 8863 20034 8889
rect 20006 8778 20034 8863
rect 20006 8745 20034 8750
rect 18942 8415 18943 8441
rect 18969 8415 18970 8441
rect 18942 8409 18970 8415
rect 20006 8442 20034 8447
rect 14910 8359 14911 8385
rect 14937 8359 14938 8385
rect 14910 8353 14938 8359
rect 20006 8385 20034 8414
rect 20006 8359 20007 8385
rect 20033 8359 20034 8385
rect 20006 8353 20034 8359
rect 17598 8246 17730 8251
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17598 8213 17730 8218
rect 17598 7462 17730 7467
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17598 7429 17730 7434
rect 13342 7154 13370 7159
rect 13286 7153 13370 7154
rect 13286 7127 13343 7153
rect 13369 7127 13370 7153
rect 13286 7126 13370 7127
rect 13174 6874 13202 6879
rect 13202 6846 13314 6874
rect 13174 6841 13202 6846
rect 12950 6622 13146 6650
rect 12950 4214 12978 6622
rect 13286 6537 13314 6846
rect 13286 6511 13287 6537
rect 13313 6511 13314 6537
rect 13286 6505 13314 6511
rect 13342 6538 13370 7126
rect 14294 6930 14322 6935
rect 13510 6538 13538 6543
rect 13342 6537 13538 6538
rect 13342 6511 13511 6537
rect 13537 6511 13538 6537
rect 13342 6510 13538 6511
rect 13342 6482 13370 6510
rect 13510 6505 13538 6510
rect 13342 6449 13370 6454
rect 10934 4186 11242 4214
rect 12614 4186 12698 4214
rect 12894 4186 12978 4214
rect 10934 2169 10962 4186
rect 10934 2143 10935 2169
rect 10961 2143 10962 2169
rect 10934 2137 10962 2143
rect 10710 1751 10711 1777
rect 10737 1751 10738 1777
rect 10710 1745 10738 1751
rect 10766 2058 10794 2063
rect 8414 1722 8442 1727
rect 8414 400 8442 1694
rect 9030 1722 9058 1727
rect 9030 1665 9058 1694
rect 9030 1639 9031 1665
rect 9057 1639 9058 1665
rect 9030 1633 9058 1639
rect 9918 1582 10050 1587
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 9918 1549 10050 1554
rect 10766 400 10794 2030
rect 11382 2058 11410 2063
rect 11382 2011 11410 2030
rect 12614 1777 12642 4186
rect 12894 2169 12922 4186
rect 12894 2143 12895 2169
rect 12921 2143 12922 2169
rect 12894 2137 12922 2143
rect 12614 1751 12615 1777
rect 12641 1751 12642 1777
rect 12614 1745 12642 1751
rect 12782 2058 12810 2063
rect 12446 1722 12474 1727
rect 11214 1666 11242 1671
rect 11102 1665 11242 1666
rect 11102 1639 11215 1665
rect 11241 1639 11242 1665
rect 11102 1638 11242 1639
rect 11102 400 11130 1638
rect 11214 1633 11242 1638
rect 12446 400 12474 1694
rect 12782 400 12810 2030
rect 13398 2058 13426 2063
rect 13398 2011 13426 2030
rect 13062 1833 13090 1839
rect 13062 1807 13063 1833
rect 13089 1807 13090 1833
rect 13062 1722 13090 1807
rect 13062 1689 13090 1694
rect 13118 1834 13146 1839
rect 13118 400 13146 1806
rect 14294 1777 14322 6902
rect 17598 6678 17730 6683
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17598 6645 17730 6650
rect 17598 5894 17730 5899
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17598 5861 17730 5866
rect 17598 5110 17730 5115
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17598 5077 17730 5082
rect 17598 4326 17730 4331
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17598 4293 17730 4298
rect 17598 3542 17730 3547
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17598 3509 17730 3514
rect 17598 2758 17730 2763
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17598 2725 17730 2730
rect 17598 1974 17730 1979
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17598 1941 17730 1946
rect 14686 1834 14714 1839
rect 14686 1787 14714 1806
rect 14294 1751 14295 1777
rect 14321 1751 14322 1777
rect 14294 1745 14322 1751
rect 8400 0 8456 400
rect 10752 0 10808 400
rect 11088 0 11144 400
rect 12432 0 12488 400
rect 12768 0 12824 400
rect 13104 0 13160 400
<< via2 >>
rect 2238 19221 2266 19222
rect 2238 19195 2239 19221
rect 2239 19195 2265 19221
rect 2265 19195 2266 19221
rect 2238 19194 2266 19195
rect 2290 19221 2318 19222
rect 2290 19195 2291 19221
rect 2291 19195 2317 19221
rect 2317 19195 2318 19221
rect 2290 19194 2318 19195
rect 2342 19221 2370 19222
rect 2342 19195 2343 19221
rect 2343 19195 2369 19221
rect 2369 19195 2370 19221
rect 2342 19194 2370 19195
rect 8750 19110 8778 19138
rect 9310 19137 9338 19138
rect 9310 19111 9311 19137
rect 9311 19111 9337 19137
rect 9337 19111 9338 19137
rect 9310 19110 9338 19111
rect 2238 18437 2266 18438
rect 2238 18411 2239 18437
rect 2239 18411 2265 18437
rect 2265 18411 2266 18437
rect 2238 18410 2266 18411
rect 2290 18437 2318 18438
rect 2290 18411 2291 18437
rect 2291 18411 2317 18437
rect 2317 18411 2318 18437
rect 2290 18410 2318 18411
rect 2342 18437 2370 18438
rect 2342 18411 2343 18437
rect 2343 18411 2369 18437
rect 2369 18411 2370 18437
rect 2342 18410 2370 18411
rect 2238 17653 2266 17654
rect 2238 17627 2239 17653
rect 2239 17627 2265 17653
rect 2265 17627 2266 17653
rect 2238 17626 2266 17627
rect 2290 17653 2318 17654
rect 2290 17627 2291 17653
rect 2291 17627 2317 17653
rect 2317 17627 2318 17653
rect 2290 17626 2318 17627
rect 2342 17653 2370 17654
rect 2342 17627 2343 17653
rect 2343 17627 2369 17653
rect 2369 17627 2370 17653
rect 2342 17626 2370 17627
rect 2238 16869 2266 16870
rect 2238 16843 2239 16869
rect 2239 16843 2265 16869
rect 2265 16843 2266 16869
rect 2238 16842 2266 16843
rect 2290 16869 2318 16870
rect 2290 16843 2291 16869
rect 2291 16843 2317 16869
rect 2317 16843 2318 16869
rect 2290 16842 2318 16843
rect 2342 16869 2370 16870
rect 2342 16843 2343 16869
rect 2343 16843 2369 16869
rect 2369 16843 2370 16869
rect 2342 16842 2370 16843
rect 2238 16085 2266 16086
rect 2238 16059 2239 16085
rect 2239 16059 2265 16085
rect 2265 16059 2266 16085
rect 2238 16058 2266 16059
rect 2290 16085 2318 16086
rect 2290 16059 2291 16085
rect 2291 16059 2317 16085
rect 2317 16059 2318 16085
rect 2290 16058 2318 16059
rect 2342 16085 2370 16086
rect 2342 16059 2343 16085
rect 2343 16059 2369 16085
rect 2369 16059 2370 16085
rect 2342 16058 2370 16059
rect 10094 19110 10122 19138
rect 10878 19137 10906 19138
rect 10878 19111 10879 19137
rect 10879 19111 10905 19137
rect 10905 19111 10906 19137
rect 10878 19110 10906 19111
rect 11774 19110 11802 19138
rect 9918 18829 9946 18830
rect 9918 18803 9919 18829
rect 9919 18803 9945 18829
rect 9945 18803 9946 18829
rect 9918 18802 9946 18803
rect 9970 18829 9998 18830
rect 9970 18803 9971 18829
rect 9971 18803 9997 18829
rect 9997 18803 9998 18829
rect 9970 18802 9998 18803
rect 10022 18829 10050 18830
rect 10022 18803 10023 18829
rect 10023 18803 10049 18829
rect 10049 18803 10050 18829
rect 10022 18802 10050 18803
rect 9422 18718 9450 18746
rect 10038 18745 10066 18746
rect 10038 18719 10039 18745
rect 10039 18719 10065 18745
rect 10065 18719 10066 18745
rect 10038 18718 10066 18719
rect 9918 18045 9946 18046
rect 9918 18019 9919 18045
rect 9919 18019 9945 18045
rect 9945 18019 9946 18045
rect 9918 18018 9946 18019
rect 9970 18045 9998 18046
rect 9970 18019 9971 18045
rect 9971 18019 9997 18045
rect 9997 18019 9998 18045
rect 9970 18018 9998 18019
rect 10022 18045 10050 18046
rect 10022 18019 10023 18045
rect 10023 18019 10049 18045
rect 10049 18019 10050 18045
rect 10022 18018 10050 18019
rect 9918 17261 9946 17262
rect 9918 17235 9919 17261
rect 9919 17235 9945 17261
rect 9945 17235 9946 17261
rect 9918 17234 9946 17235
rect 9970 17261 9998 17262
rect 9970 17235 9971 17261
rect 9971 17235 9997 17261
rect 9997 17235 9998 17261
rect 9970 17234 9998 17235
rect 10022 17261 10050 17262
rect 10022 17235 10023 17261
rect 10023 17235 10049 17261
rect 10049 17235 10050 17261
rect 10022 17234 10050 17235
rect 9918 16477 9946 16478
rect 9918 16451 9919 16477
rect 9919 16451 9945 16477
rect 9945 16451 9946 16477
rect 9918 16450 9946 16451
rect 9970 16477 9998 16478
rect 9970 16451 9971 16477
rect 9971 16451 9997 16477
rect 9997 16451 9998 16477
rect 9970 16450 9998 16451
rect 10022 16477 10050 16478
rect 10022 16451 10023 16477
rect 10023 16451 10049 16477
rect 10049 16451 10050 16477
rect 10022 16450 10050 16451
rect 17598 19221 17626 19222
rect 17598 19195 17599 19221
rect 17599 19195 17625 19221
rect 17625 19195 17626 19221
rect 17598 19194 17626 19195
rect 17650 19221 17678 19222
rect 17650 19195 17651 19221
rect 17651 19195 17677 19221
rect 17677 19195 17678 19221
rect 17650 19194 17678 19195
rect 17702 19221 17730 19222
rect 17702 19195 17703 19221
rect 17703 19195 17729 19221
rect 17729 19195 17730 19221
rect 17702 19194 17730 19195
rect 12782 19137 12810 19138
rect 12782 19111 12783 19137
rect 12783 19111 12809 19137
rect 12809 19111 12810 19137
rect 12782 19110 12810 19111
rect 12110 18718 12138 18746
rect 13118 18745 13146 18746
rect 13118 18719 13119 18745
rect 13119 18719 13145 18745
rect 13145 18719 13146 18745
rect 13118 18718 13146 18719
rect 2238 15301 2266 15302
rect 2238 15275 2239 15301
rect 2239 15275 2265 15301
rect 2265 15275 2266 15301
rect 2238 15274 2266 15275
rect 2290 15301 2318 15302
rect 2290 15275 2291 15301
rect 2291 15275 2317 15301
rect 2317 15275 2318 15301
rect 2290 15274 2318 15275
rect 2342 15301 2370 15302
rect 2342 15275 2343 15301
rect 2343 15275 2369 15301
rect 2369 15275 2370 15301
rect 2342 15274 2370 15275
rect 2238 14517 2266 14518
rect 2238 14491 2239 14517
rect 2239 14491 2265 14517
rect 2265 14491 2266 14517
rect 2238 14490 2266 14491
rect 2290 14517 2318 14518
rect 2290 14491 2291 14517
rect 2291 14491 2317 14517
rect 2317 14491 2318 14517
rect 2290 14490 2318 14491
rect 2342 14517 2370 14518
rect 2342 14491 2343 14517
rect 2343 14491 2369 14517
rect 2369 14491 2370 14517
rect 2342 14490 2370 14491
rect 2086 13790 2114 13818
rect 966 12249 994 12250
rect 966 12223 967 12249
rect 967 12223 993 12249
rect 993 12223 994 12249
rect 966 12222 994 12223
rect 966 11774 994 11802
rect 2238 13733 2266 13734
rect 2238 13707 2239 13733
rect 2239 13707 2265 13733
rect 2265 13707 2266 13733
rect 2238 13706 2266 13707
rect 2290 13733 2318 13734
rect 2290 13707 2291 13733
rect 2291 13707 2317 13733
rect 2317 13707 2318 13733
rect 2290 13706 2318 13707
rect 2342 13733 2370 13734
rect 2342 13707 2343 13733
rect 2343 13707 2369 13733
rect 2369 13707 2370 13733
rect 2342 13706 2370 13707
rect 8078 13454 8106 13482
rect 8470 13454 8498 13482
rect 8414 13062 8442 13090
rect 2238 12949 2266 12950
rect 2238 12923 2239 12949
rect 2239 12923 2265 12949
rect 2265 12923 2266 12949
rect 2238 12922 2266 12923
rect 2290 12949 2318 12950
rect 2290 12923 2291 12949
rect 2291 12923 2317 12949
rect 2317 12923 2318 12949
rect 2290 12922 2318 12923
rect 2342 12949 2370 12950
rect 2342 12923 2343 12949
rect 2343 12923 2369 12949
rect 2369 12923 2370 12949
rect 2342 12922 2370 12923
rect 9142 13873 9170 13874
rect 9142 13847 9143 13873
rect 9143 13847 9169 13873
rect 9169 13847 9170 13873
rect 9142 13846 9170 13847
rect 9918 15693 9946 15694
rect 9918 15667 9919 15693
rect 9919 15667 9945 15693
rect 9945 15667 9946 15693
rect 9918 15666 9946 15667
rect 9970 15693 9998 15694
rect 9970 15667 9971 15693
rect 9971 15667 9997 15693
rect 9997 15667 9998 15693
rect 9970 15666 9998 15667
rect 10022 15693 10050 15694
rect 10022 15667 10023 15693
rect 10023 15667 10049 15693
rect 10049 15667 10050 15693
rect 10022 15666 10050 15667
rect 9918 14909 9946 14910
rect 9918 14883 9919 14909
rect 9919 14883 9945 14909
rect 9945 14883 9946 14909
rect 9918 14882 9946 14883
rect 9970 14909 9998 14910
rect 9970 14883 9971 14909
rect 9971 14883 9997 14909
rect 9997 14883 9998 14909
rect 9970 14882 9998 14883
rect 10022 14909 10050 14910
rect 10022 14883 10023 14909
rect 10023 14883 10049 14909
rect 10049 14883 10050 14909
rect 10022 14882 10050 14883
rect 9918 14125 9946 14126
rect 9918 14099 9919 14125
rect 9919 14099 9945 14125
rect 9945 14099 9946 14125
rect 9918 14098 9946 14099
rect 9970 14125 9998 14126
rect 9970 14099 9971 14125
rect 9971 14099 9997 14125
rect 9997 14099 9998 14125
rect 9970 14098 9998 14099
rect 10022 14125 10050 14126
rect 10022 14099 10023 14125
rect 10023 14099 10049 14125
rect 10049 14099 10050 14125
rect 10022 14098 10050 14099
rect 9926 13846 9954 13874
rect 8862 13454 8890 13482
rect 2142 12361 2170 12362
rect 2142 12335 2143 12361
rect 2143 12335 2169 12361
rect 2169 12335 2170 12361
rect 2142 12334 2170 12335
rect 6902 12334 6930 12362
rect 7182 12334 7210 12362
rect 2238 12165 2266 12166
rect 2238 12139 2239 12165
rect 2239 12139 2265 12165
rect 2265 12139 2266 12165
rect 2238 12138 2266 12139
rect 2290 12165 2318 12166
rect 2290 12139 2291 12165
rect 2291 12139 2317 12165
rect 2317 12139 2318 12165
rect 2290 12138 2318 12139
rect 2342 12165 2370 12166
rect 2342 12139 2343 12165
rect 2343 12139 2369 12165
rect 2369 12139 2370 12165
rect 2342 12138 2370 12139
rect 6790 11662 6818 11690
rect 2142 11494 2170 11522
rect 5670 11550 5698 11578
rect 8414 12446 8442 12474
rect 8302 12361 8330 12362
rect 8302 12335 8303 12361
rect 8303 12335 8329 12361
rect 8329 12335 8330 12361
rect 8302 12334 8330 12335
rect 8638 12278 8666 12306
rect 7686 11718 7714 11746
rect 7574 11689 7602 11690
rect 7574 11663 7575 11689
rect 7575 11663 7601 11689
rect 7601 11663 7602 11689
rect 7574 11662 7602 11663
rect 9702 13481 9730 13482
rect 9702 13455 9703 13481
rect 9703 13455 9729 13481
rect 9729 13455 9730 13481
rect 9702 13454 9730 13455
rect 9366 13145 9394 13146
rect 9366 13119 9367 13145
rect 9367 13119 9393 13145
rect 9393 13119 9394 13145
rect 9366 13118 9394 13119
rect 9086 12558 9114 12586
rect 9142 12473 9170 12474
rect 9142 12447 9143 12473
rect 9143 12447 9169 12473
rect 9169 12447 9170 12473
rect 9142 12446 9170 12447
rect 8750 12361 8778 12362
rect 8750 12335 8751 12361
rect 8751 12335 8777 12361
rect 8777 12335 8778 12361
rect 8750 12334 8778 12335
rect 8918 11969 8946 11970
rect 8918 11943 8919 11969
rect 8919 11943 8945 11969
rect 8945 11943 8946 11969
rect 8918 11942 8946 11943
rect 8078 11830 8106 11858
rect 7910 11718 7938 11746
rect 8918 11857 8946 11858
rect 8918 11831 8919 11857
rect 8919 11831 8945 11857
rect 8945 11831 8946 11857
rect 8918 11830 8946 11831
rect 8302 11718 8330 11746
rect 7630 11633 7658 11634
rect 7630 11607 7631 11633
rect 7631 11607 7657 11633
rect 7657 11607 7658 11633
rect 7630 11606 7658 11607
rect 7406 11577 7434 11578
rect 7406 11551 7407 11577
rect 7407 11551 7433 11577
rect 7433 11551 7434 11577
rect 7406 11550 7434 11551
rect 2238 11381 2266 11382
rect 2238 11355 2239 11381
rect 2239 11355 2265 11381
rect 2265 11355 2266 11381
rect 2238 11354 2266 11355
rect 2290 11381 2318 11382
rect 2290 11355 2291 11381
rect 2291 11355 2317 11381
rect 2317 11355 2318 11381
rect 2290 11354 2318 11355
rect 2342 11381 2370 11382
rect 2342 11355 2343 11381
rect 2343 11355 2369 11381
rect 2369 11355 2370 11381
rect 2342 11354 2370 11355
rect 6454 10793 6482 10794
rect 6454 10767 6455 10793
rect 6455 10767 6481 10793
rect 6481 10767 6482 10793
rect 6454 10766 6482 10767
rect 2238 10597 2266 10598
rect 2238 10571 2239 10597
rect 2239 10571 2265 10597
rect 2265 10571 2266 10597
rect 2238 10570 2266 10571
rect 2290 10597 2318 10598
rect 2290 10571 2291 10597
rect 2291 10571 2317 10597
rect 2317 10571 2318 10597
rect 2290 10570 2318 10571
rect 2342 10597 2370 10598
rect 2342 10571 2343 10597
rect 2343 10571 2369 10597
rect 2369 10571 2370 10597
rect 2342 10570 2370 10571
rect 6510 10374 6538 10402
rect 5390 10345 5418 10346
rect 5390 10319 5391 10345
rect 5391 10319 5417 10345
rect 5417 10319 5418 10345
rect 5390 10318 5418 10319
rect 5054 10094 5082 10122
rect 5390 10009 5418 10010
rect 5390 9983 5391 10009
rect 5391 9983 5417 10009
rect 5417 9983 5418 10009
rect 5390 9982 5418 9983
rect 2086 9926 2114 9954
rect 7518 11326 7546 11354
rect 7966 11382 7994 11410
rect 8302 11270 8330 11298
rect 8358 11606 8386 11634
rect 7686 10878 7714 10906
rect 7294 10793 7322 10794
rect 7294 10767 7295 10793
rect 7295 10767 7321 10793
rect 7321 10767 7322 10793
rect 7294 10766 7322 10767
rect 6790 10401 6818 10402
rect 6790 10375 6791 10401
rect 6791 10375 6817 10401
rect 6817 10375 6818 10401
rect 6790 10374 6818 10375
rect 7238 10430 7266 10458
rect 7294 10345 7322 10346
rect 7294 10319 7295 10345
rect 7295 10319 7321 10345
rect 7321 10319 7322 10345
rect 7294 10318 7322 10319
rect 6958 10150 6986 10178
rect 6902 10094 6930 10122
rect 6734 9982 6762 10010
rect 2238 9813 2266 9814
rect 2238 9787 2239 9813
rect 2239 9787 2265 9813
rect 2265 9787 2266 9813
rect 2238 9786 2266 9787
rect 2290 9813 2318 9814
rect 2290 9787 2291 9813
rect 2291 9787 2317 9813
rect 2317 9787 2318 9813
rect 2290 9786 2318 9787
rect 2342 9813 2370 9814
rect 2342 9787 2343 9813
rect 2343 9787 2369 9813
rect 2369 9787 2370 9813
rect 2342 9786 2370 9787
rect 6734 9366 6762 9394
rect 7462 10094 7490 10122
rect 7294 9617 7322 9618
rect 7294 9591 7295 9617
rect 7295 9591 7321 9617
rect 7321 9591 7322 9617
rect 7294 9590 7322 9591
rect 2238 9029 2266 9030
rect 2238 9003 2239 9029
rect 2239 9003 2265 9029
rect 2265 9003 2266 9029
rect 2238 9002 2266 9003
rect 2290 9029 2318 9030
rect 2290 9003 2291 9029
rect 2291 9003 2317 9029
rect 2317 9003 2318 9029
rect 2290 9002 2318 9003
rect 2342 9029 2370 9030
rect 2342 9003 2343 9029
rect 2343 9003 2369 9029
rect 2369 9003 2370 9029
rect 2342 9002 2370 9003
rect 966 8889 994 8890
rect 966 8863 967 8889
rect 967 8863 993 8889
rect 993 8863 994 8889
rect 966 8862 994 8863
rect 2142 8833 2170 8834
rect 2142 8807 2143 8833
rect 2143 8807 2169 8833
rect 2169 8807 2170 8833
rect 2142 8806 2170 8807
rect 4998 8806 5026 8834
rect 966 8078 994 8106
rect 6398 8833 6426 8834
rect 6398 8807 6399 8833
rect 6399 8807 6425 8833
rect 6425 8807 6426 8833
rect 6398 8806 6426 8807
rect 6734 8806 6762 8834
rect 4998 8414 5026 8442
rect 5782 8694 5810 8722
rect 7126 9366 7154 9394
rect 7406 9478 7434 9506
rect 7462 9254 7490 9282
rect 2238 8245 2266 8246
rect 2238 8219 2239 8245
rect 2239 8219 2265 8245
rect 2265 8219 2266 8245
rect 2238 8218 2266 8219
rect 2290 8245 2318 8246
rect 2290 8219 2291 8245
rect 2291 8219 2317 8245
rect 2317 8219 2318 8245
rect 2290 8218 2318 8219
rect 2342 8245 2370 8246
rect 2342 8219 2343 8245
rect 2343 8219 2369 8245
rect 2369 8219 2370 8245
rect 2342 8218 2370 8219
rect 6398 7910 6426 7938
rect 2142 7574 2170 7602
rect 5334 7742 5362 7770
rect 7350 8862 7378 8890
rect 7406 8750 7434 8778
rect 7126 8721 7154 8722
rect 7126 8695 7127 8721
rect 7127 8695 7153 8721
rect 7153 8695 7154 8721
rect 7126 8694 7154 8695
rect 7126 8470 7154 8498
rect 7070 8441 7098 8442
rect 7070 8415 7071 8441
rect 7071 8415 7097 8441
rect 7097 8415 7098 8441
rect 7070 8414 7098 8415
rect 8806 11214 8834 11242
rect 8134 10849 8162 10850
rect 8134 10823 8135 10849
rect 8135 10823 8161 10849
rect 8161 10823 8162 10849
rect 8134 10822 8162 10823
rect 8414 10849 8442 10850
rect 8414 10823 8415 10849
rect 8415 10823 8441 10849
rect 8441 10823 8442 10849
rect 8414 10822 8442 10823
rect 8022 10793 8050 10794
rect 8022 10767 8023 10793
rect 8023 10767 8049 10793
rect 8049 10767 8050 10793
rect 8022 10766 8050 10767
rect 7742 10457 7770 10458
rect 7742 10431 7743 10457
rect 7743 10431 7769 10457
rect 7769 10431 7770 10457
rect 7742 10430 7770 10431
rect 8918 10905 8946 10906
rect 8918 10879 8919 10905
rect 8919 10879 8945 10905
rect 8945 10879 8946 10905
rect 8918 10878 8946 10879
rect 8470 10710 8498 10738
rect 8022 10094 8050 10122
rect 8078 10318 8106 10346
rect 8246 9953 8274 9954
rect 8246 9927 8247 9953
rect 8247 9927 8273 9953
rect 8273 9927 8274 9953
rect 8246 9926 8274 9927
rect 8302 9702 8330 9730
rect 7574 9113 7602 9114
rect 7574 9087 7575 9113
rect 7575 9087 7601 9113
rect 7601 9087 7602 9113
rect 7574 9086 7602 9087
rect 8190 9198 8218 9226
rect 7854 8553 7882 8554
rect 7854 8527 7855 8553
rect 7855 8527 7881 8553
rect 7881 8527 7882 8553
rect 7854 8526 7882 8527
rect 7910 9142 7938 9170
rect 9198 11913 9226 11914
rect 9198 11887 9199 11913
rect 9199 11887 9225 11913
rect 9225 11887 9226 11913
rect 9198 11886 9226 11887
rect 9534 13089 9562 13090
rect 9534 13063 9535 13089
rect 9535 13063 9561 13089
rect 9561 13063 9562 13089
rect 9534 13062 9562 13063
rect 9918 13341 9946 13342
rect 9918 13315 9919 13341
rect 9919 13315 9945 13341
rect 9945 13315 9946 13341
rect 9918 13314 9946 13315
rect 9970 13341 9998 13342
rect 9970 13315 9971 13341
rect 9971 13315 9997 13341
rect 9997 13315 9998 13341
rect 9970 13314 9998 13315
rect 10022 13341 10050 13342
rect 10022 13315 10023 13341
rect 10023 13315 10049 13341
rect 10049 13315 10050 13341
rect 10022 13314 10050 13315
rect 10094 13118 10122 13146
rect 10934 14265 10962 14266
rect 10934 14239 10935 14265
rect 10935 14239 10961 14265
rect 10961 14239 10962 14265
rect 10934 14238 10962 14239
rect 17598 18437 17626 18438
rect 17598 18411 17599 18437
rect 17599 18411 17625 18437
rect 17625 18411 17626 18437
rect 17598 18410 17626 18411
rect 17650 18437 17678 18438
rect 17650 18411 17651 18437
rect 17651 18411 17677 18437
rect 17677 18411 17678 18437
rect 17650 18410 17678 18411
rect 17702 18437 17730 18438
rect 17702 18411 17703 18437
rect 17703 18411 17729 18437
rect 17729 18411 17730 18437
rect 17702 18410 17730 18411
rect 17598 17653 17626 17654
rect 17598 17627 17599 17653
rect 17599 17627 17625 17653
rect 17625 17627 17626 17653
rect 17598 17626 17626 17627
rect 17650 17653 17678 17654
rect 17650 17627 17651 17653
rect 17651 17627 17677 17653
rect 17677 17627 17678 17653
rect 17650 17626 17678 17627
rect 17702 17653 17730 17654
rect 17702 17627 17703 17653
rect 17703 17627 17729 17653
rect 17729 17627 17730 17653
rect 17702 17626 17730 17627
rect 17598 16869 17626 16870
rect 17598 16843 17599 16869
rect 17599 16843 17625 16869
rect 17625 16843 17626 16869
rect 17598 16842 17626 16843
rect 17650 16869 17678 16870
rect 17650 16843 17651 16869
rect 17651 16843 17677 16869
rect 17677 16843 17678 16869
rect 17650 16842 17678 16843
rect 17702 16869 17730 16870
rect 17702 16843 17703 16869
rect 17703 16843 17729 16869
rect 17729 16843 17730 16869
rect 17702 16842 17730 16843
rect 17598 16085 17626 16086
rect 17598 16059 17599 16085
rect 17599 16059 17625 16085
rect 17625 16059 17626 16085
rect 17598 16058 17626 16059
rect 17650 16085 17678 16086
rect 17650 16059 17651 16085
rect 17651 16059 17677 16085
rect 17677 16059 17678 16085
rect 17650 16058 17678 16059
rect 17702 16085 17730 16086
rect 17702 16059 17703 16085
rect 17703 16059 17729 16085
rect 17729 16059 17730 16085
rect 17702 16058 17730 16059
rect 17598 15301 17626 15302
rect 17598 15275 17599 15301
rect 17599 15275 17625 15301
rect 17625 15275 17626 15301
rect 17598 15274 17626 15275
rect 17650 15301 17678 15302
rect 17650 15275 17651 15301
rect 17651 15275 17677 15301
rect 17677 15275 17678 15301
rect 17650 15274 17678 15275
rect 17702 15301 17730 15302
rect 17702 15275 17703 15301
rect 17703 15275 17729 15301
rect 17729 15275 17730 15301
rect 17702 15274 17730 15275
rect 17598 14517 17626 14518
rect 17598 14491 17599 14517
rect 17599 14491 17625 14517
rect 17625 14491 17626 14517
rect 17598 14490 17626 14491
rect 17650 14517 17678 14518
rect 17650 14491 17651 14517
rect 17651 14491 17677 14517
rect 17677 14491 17678 14517
rect 17650 14490 17678 14491
rect 17702 14517 17730 14518
rect 17702 14491 17703 14517
rect 17703 14491 17729 14517
rect 17729 14491 17730 14517
rect 17702 14490 17730 14491
rect 11830 14238 11858 14266
rect 10430 13510 10458 13538
rect 11886 13566 11914 13594
rect 10934 13537 10962 13538
rect 10934 13511 10935 13537
rect 10935 13511 10961 13537
rect 10961 13511 10962 13537
rect 10934 13510 10962 13511
rect 17598 13733 17626 13734
rect 17598 13707 17599 13733
rect 17599 13707 17625 13733
rect 17625 13707 17626 13733
rect 17598 13706 17626 13707
rect 17650 13733 17678 13734
rect 17650 13707 17651 13733
rect 17651 13707 17677 13733
rect 17677 13707 17678 13733
rect 17650 13706 17678 13707
rect 17702 13733 17730 13734
rect 17702 13707 17703 13733
rect 17703 13707 17729 13733
rect 17729 13707 17730 13733
rect 17702 13706 17730 13707
rect 12334 13593 12362 13594
rect 12334 13567 12335 13593
rect 12335 13567 12361 13593
rect 12361 13567 12362 13593
rect 12334 13566 12362 13567
rect 12110 13510 12138 13538
rect 12558 13537 12586 13538
rect 12558 13511 12559 13537
rect 12559 13511 12585 13537
rect 12585 13511 12586 13537
rect 12558 13510 12586 13511
rect 12894 13537 12922 13538
rect 12894 13511 12895 13537
rect 12895 13511 12921 13537
rect 12921 13511 12922 13537
rect 12894 13510 12922 13511
rect 14350 13510 14378 13538
rect 14574 13510 14602 13538
rect 10878 13201 10906 13202
rect 10878 13175 10879 13201
rect 10879 13175 10905 13201
rect 10905 13175 10906 13201
rect 10878 13174 10906 13175
rect 9646 12446 9674 12474
rect 9702 12614 9730 12642
rect 9310 11886 9338 11914
rect 9198 11718 9226 11746
rect 9086 11662 9114 11690
rect 9086 11297 9114 11298
rect 9086 11271 9087 11297
rect 9087 11271 9113 11297
rect 9113 11271 9114 11297
rect 9086 11270 9114 11271
rect 9198 11241 9226 11242
rect 9198 11215 9199 11241
rect 9199 11215 9225 11241
rect 9225 11215 9226 11241
rect 9198 11214 9226 11215
rect 9086 10793 9114 10794
rect 9086 10767 9087 10793
rect 9087 10767 9113 10793
rect 9113 10767 9114 10793
rect 9086 10766 9114 10767
rect 8974 10710 9002 10738
rect 8750 10094 8778 10122
rect 8526 9926 8554 9954
rect 8414 9702 8442 9730
rect 8358 9142 8386 9170
rect 8806 10009 8834 10010
rect 8806 9983 8807 10009
rect 8807 9983 8833 10009
rect 8833 9983 8834 10009
rect 8806 9982 8834 9983
rect 8862 9254 8890 9282
rect 8638 9142 8666 9170
rect 8582 8777 8610 8778
rect 8582 8751 8583 8777
rect 8583 8751 8609 8777
rect 8609 8751 8610 8777
rect 8582 8750 8610 8751
rect 8414 8470 8442 8498
rect 8694 8918 8722 8946
rect 9310 11185 9338 11186
rect 9310 11159 9311 11185
rect 9311 11159 9337 11185
rect 9337 11159 9338 11185
rect 9310 11158 9338 11159
rect 9366 11438 9394 11466
rect 9254 10121 9282 10122
rect 9254 10095 9255 10121
rect 9255 10095 9281 10121
rect 9281 10095 9282 10121
rect 9254 10094 9282 10095
rect 9030 9366 9058 9394
rect 8974 9254 9002 9282
rect 8750 8553 8778 8554
rect 8750 8527 8751 8553
rect 8751 8527 8777 8553
rect 8777 8527 8778 8553
rect 8750 8526 8778 8527
rect 7182 7993 7210 7994
rect 7182 7967 7183 7993
rect 7183 7967 7209 7993
rect 7209 7967 7210 7993
rect 7182 7966 7210 7967
rect 7686 7993 7714 7994
rect 7686 7967 7687 7993
rect 7687 7967 7713 7993
rect 7713 7967 7714 7993
rect 7686 7966 7714 7967
rect 7070 7937 7098 7938
rect 7070 7911 7071 7937
rect 7071 7911 7097 7937
rect 7097 7911 7098 7937
rect 7070 7910 7098 7911
rect 6790 7742 6818 7770
rect 5334 7601 5362 7602
rect 5334 7575 5335 7601
rect 5335 7575 5361 7601
rect 5361 7575 5362 7601
rect 5334 7574 5362 7575
rect 2238 7461 2266 7462
rect 2238 7435 2239 7461
rect 2239 7435 2265 7461
rect 2265 7435 2266 7461
rect 2238 7434 2266 7435
rect 2290 7461 2318 7462
rect 2290 7435 2291 7461
rect 2291 7435 2317 7461
rect 2317 7435 2318 7461
rect 2290 7434 2318 7435
rect 2342 7461 2370 7462
rect 2342 7435 2343 7461
rect 2343 7435 2369 7461
rect 2369 7435 2370 7461
rect 2342 7434 2370 7435
rect 8470 7518 8498 7546
rect 7014 7294 7042 7322
rect 7294 7294 7322 7322
rect 2238 6677 2266 6678
rect 2238 6651 2239 6677
rect 2239 6651 2265 6677
rect 2265 6651 2266 6677
rect 2238 6650 2266 6651
rect 2290 6677 2318 6678
rect 2290 6651 2291 6677
rect 2291 6651 2317 6677
rect 2317 6651 2318 6677
rect 2290 6650 2318 6651
rect 2342 6677 2370 6678
rect 2342 6651 2343 6677
rect 2343 6651 2369 6677
rect 2369 6651 2370 6677
rect 2342 6650 2370 6651
rect 8246 7294 8274 7322
rect 9198 9198 9226 9226
rect 9198 8806 9226 8834
rect 9310 9702 9338 9730
rect 9534 11662 9562 11690
rect 9646 11662 9674 11690
rect 9590 11633 9618 11634
rect 9590 11607 9591 11633
rect 9591 11607 9617 11633
rect 9617 11607 9618 11633
rect 9590 11606 9618 11607
rect 9870 12697 9898 12698
rect 9870 12671 9871 12697
rect 9871 12671 9897 12697
rect 9897 12671 9898 12697
rect 9870 12670 9898 12671
rect 9926 12614 9954 12642
rect 9918 12557 9946 12558
rect 9918 12531 9919 12557
rect 9919 12531 9945 12557
rect 9945 12531 9946 12557
rect 9918 12530 9946 12531
rect 9970 12557 9998 12558
rect 9970 12531 9971 12557
rect 9971 12531 9997 12557
rect 9997 12531 9998 12557
rect 9970 12530 9998 12531
rect 10022 12557 10050 12558
rect 10022 12531 10023 12557
rect 10023 12531 10049 12557
rect 10049 12531 10050 12557
rect 10022 12530 10050 12531
rect 10038 12446 10066 12474
rect 10262 12390 10290 12418
rect 10318 12670 10346 12698
rect 10094 12334 10122 12362
rect 10430 12473 10458 12474
rect 10430 12447 10431 12473
rect 10431 12447 10457 12473
rect 10457 12447 10458 12473
rect 10430 12446 10458 12447
rect 10094 11942 10122 11970
rect 9758 11886 9786 11914
rect 9702 11465 9730 11466
rect 9702 11439 9703 11465
rect 9703 11439 9729 11465
rect 9729 11439 9730 11465
rect 9702 11438 9730 11439
rect 9422 11326 9450 11354
rect 9478 11214 9506 11242
rect 9422 10009 9450 10010
rect 9422 9983 9423 10009
rect 9423 9983 9449 10009
rect 9449 9983 9450 10009
rect 9422 9982 9450 9983
rect 9646 9702 9674 9730
rect 9702 9926 9730 9954
rect 9310 9225 9338 9226
rect 9310 9199 9311 9225
rect 9311 9199 9337 9225
rect 9337 9199 9338 9225
rect 9310 9198 9338 9199
rect 9534 9478 9562 9506
rect 9534 9366 9562 9394
rect 9702 9366 9730 9394
rect 9478 8974 9506 9002
rect 9590 8918 9618 8946
rect 9478 8833 9506 8834
rect 9478 8807 9479 8833
rect 9479 8807 9505 8833
rect 9505 8807 9506 8833
rect 9478 8806 9506 8807
rect 9198 8470 9226 8498
rect 9198 8358 9226 8386
rect 9534 8385 9562 8386
rect 9534 8359 9535 8385
rect 9535 8359 9561 8385
rect 9561 8359 9562 8385
rect 9534 8358 9562 8359
rect 9926 11913 9954 11914
rect 9926 11887 9927 11913
rect 9927 11887 9953 11913
rect 9953 11887 9954 11913
rect 9926 11886 9954 11887
rect 9918 11773 9946 11774
rect 9918 11747 9919 11773
rect 9919 11747 9945 11773
rect 9945 11747 9946 11773
rect 9918 11746 9946 11747
rect 9970 11773 9998 11774
rect 9970 11747 9971 11773
rect 9971 11747 9997 11773
rect 9997 11747 9998 11773
rect 9970 11746 9998 11747
rect 10022 11773 10050 11774
rect 10022 11747 10023 11773
rect 10023 11747 10049 11773
rect 10049 11747 10050 11773
rect 10022 11746 10050 11747
rect 9814 11214 9842 11242
rect 9982 11214 10010 11242
rect 9926 11185 9954 11186
rect 9926 11159 9927 11185
rect 9927 11159 9953 11185
rect 9953 11159 9954 11185
rect 9926 11158 9954 11159
rect 10094 11270 10122 11298
rect 10094 11185 10122 11186
rect 10094 11159 10095 11185
rect 10095 11159 10121 11185
rect 10121 11159 10122 11185
rect 10094 11158 10122 11159
rect 9982 11102 10010 11130
rect 10822 13118 10850 13146
rect 11158 13145 11186 13146
rect 11158 13119 11159 13145
rect 11159 13119 11185 13145
rect 11185 13119 11186 13145
rect 11158 13118 11186 13119
rect 11382 13145 11410 13146
rect 11382 13119 11383 13145
rect 11383 13119 11409 13145
rect 11409 13119 11410 13145
rect 11382 13118 11410 13119
rect 11774 13145 11802 13146
rect 11774 13119 11775 13145
rect 11775 13119 11801 13145
rect 11801 13119 11802 13145
rect 11774 13118 11802 13119
rect 11438 12838 11466 12866
rect 10654 12697 10682 12698
rect 10654 12671 10655 12697
rect 10655 12671 10681 12697
rect 10681 12671 10682 12697
rect 10654 12670 10682 12671
rect 10654 12446 10682 12474
rect 11942 12838 11970 12866
rect 10710 12417 10738 12418
rect 10710 12391 10711 12417
rect 10711 12391 10737 12417
rect 10737 12391 10738 12417
rect 10710 12390 10738 12391
rect 10878 12361 10906 12362
rect 10878 12335 10879 12361
rect 10879 12335 10905 12361
rect 10905 12335 10906 12361
rect 10878 12334 10906 12335
rect 11270 12361 11298 12362
rect 11270 12335 11271 12361
rect 11271 12335 11297 12361
rect 11297 12335 11298 12361
rect 11270 12334 11298 12335
rect 18830 13537 18858 13538
rect 18830 13511 18831 13537
rect 18831 13511 18857 13537
rect 18857 13511 18858 13537
rect 18830 13510 18858 13511
rect 14070 12838 14098 12866
rect 13734 12782 13762 12810
rect 13286 12753 13314 12754
rect 13286 12727 13287 12753
rect 13287 12727 13313 12753
rect 13313 12727 13314 12753
rect 13286 12726 13314 12727
rect 13566 12697 13594 12698
rect 13566 12671 13567 12697
rect 13567 12671 13593 12697
rect 13593 12671 13594 12697
rect 13566 12670 13594 12671
rect 13230 12641 13258 12642
rect 13230 12615 13231 12641
rect 13231 12615 13257 12641
rect 13257 12615 13258 12641
rect 13230 12614 13258 12615
rect 13454 12641 13482 12642
rect 13454 12615 13455 12641
rect 13455 12615 13481 12641
rect 13481 12615 13482 12641
rect 13454 12614 13482 12615
rect 13678 12614 13706 12642
rect 12950 12278 12978 12306
rect 13398 12278 13426 12306
rect 10598 11886 10626 11914
rect 10374 11577 10402 11578
rect 10374 11551 10375 11577
rect 10375 11551 10401 11577
rect 10401 11551 10402 11577
rect 10374 11550 10402 11551
rect 10430 11438 10458 11466
rect 10206 11270 10234 11298
rect 10262 11326 10290 11354
rect 9918 10989 9946 10990
rect 9918 10963 9919 10989
rect 9919 10963 9945 10989
rect 9945 10963 9946 10989
rect 9918 10962 9946 10963
rect 9970 10989 9998 10990
rect 9970 10963 9971 10989
rect 9971 10963 9997 10989
rect 9997 10963 9998 10989
rect 9970 10962 9998 10963
rect 10022 10989 10050 10990
rect 10022 10963 10023 10989
rect 10023 10963 10049 10989
rect 10049 10963 10050 10989
rect 10022 10962 10050 10963
rect 10262 10878 10290 10906
rect 10038 10401 10066 10402
rect 10038 10375 10039 10401
rect 10039 10375 10065 10401
rect 10065 10375 10066 10401
rect 10038 10374 10066 10375
rect 10094 10262 10122 10290
rect 10318 10766 10346 10794
rect 9918 10205 9946 10206
rect 9918 10179 9919 10205
rect 9919 10179 9945 10205
rect 9945 10179 9946 10205
rect 9918 10178 9946 10179
rect 9970 10205 9998 10206
rect 9970 10179 9971 10205
rect 9971 10179 9997 10205
rect 9997 10179 9998 10205
rect 9970 10178 9998 10179
rect 10022 10205 10050 10206
rect 10022 10179 10023 10205
rect 10023 10179 10049 10205
rect 10049 10179 10050 10205
rect 10022 10178 10050 10179
rect 10150 9646 10178 9674
rect 9918 9421 9946 9422
rect 9918 9395 9919 9421
rect 9919 9395 9945 9421
rect 9945 9395 9946 9421
rect 9918 9394 9946 9395
rect 9970 9421 9998 9422
rect 9970 9395 9971 9421
rect 9971 9395 9997 9421
rect 9997 9395 9998 9421
rect 9970 9394 9998 9395
rect 10022 9421 10050 9422
rect 10022 9395 10023 9421
rect 10023 9395 10049 9421
rect 10049 9395 10050 9421
rect 10022 9394 10050 9395
rect 9814 9310 9842 9338
rect 9870 9254 9898 9282
rect 9814 9225 9842 9226
rect 9814 9199 9815 9225
rect 9815 9199 9841 9225
rect 9841 9199 9842 9225
rect 9814 9198 9842 9199
rect 9758 8889 9786 8890
rect 9758 8863 9759 8889
rect 9759 8863 9785 8889
rect 9785 8863 9786 8889
rect 9758 8862 9786 8863
rect 9926 8833 9954 8834
rect 9926 8807 9927 8833
rect 9927 8807 9953 8833
rect 9953 8807 9954 8833
rect 9926 8806 9954 8807
rect 10486 10766 10514 10794
rect 10430 10318 10458 10346
rect 10206 9590 10234 9618
rect 10374 9702 10402 9730
rect 10206 9254 10234 9282
rect 10542 9478 10570 9506
rect 11662 11830 11690 11858
rect 10934 11494 10962 11522
rect 10822 11270 10850 11298
rect 10710 11158 10738 11186
rect 10654 11129 10682 11130
rect 10654 11103 10655 11129
rect 10655 11103 10681 11129
rect 10681 11103 10682 11129
rect 10654 11102 10682 11103
rect 10822 11073 10850 11074
rect 10822 11047 10823 11073
rect 10823 11047 10849 11073
rect 10849 11047 10850 11073
rect 10822 11046 10850 11047
rect 10710 10766 10738 10794
rect 10990 11102 11018 11130
rect 11830 11382 11858 11410
rect 10654 9646 10682 9674
rect 10598 9310 10626 9338
rect 9918 8637 9946 8638
rect 9918 8611 9919 8637
rect 9919 8611 9945 8637
rect 9945 8611 9946 8637
rect 9918 8610 9946 8611
rect 9970 8637 9998 8638
rect 9970 8611 9971 8637
rect 9971 8611 9997 8637
rect 9997 8611 9998 8637
rect 9970 8610 9998 8611
rect 10022 8637 10050 8638
rect 10022 8611 10023 8637
rect 10023 8611 10049 8637
rect 10049 8611 10050 8637
rect 10022 8610 10050 8611
rect 10878 10457 10906 10458
rect 10878 10431 10879 10457
rect 10879 10431 10905 10457
rect 10905 10431 10906 10457
rect 10878 10430 10906 10431
rect 10822 10289 10850 10290
rect 10822 10263 10823 10289
rect 10823 10263 10849 10289
rect 10849 10263 10850 10289
rect 10822 10262 10850 10263
rect 10766 9254 10794 9282
rect 10822 10038 10850 10066
rect 10654 9142 10682 9170
rect 10206 8750 10234 8778
rect 10262 8470 10290 8498
rect 10206 8302 10234 8330
rect 9702 8022 9730 8050
rect 9590 7910 9618 7938
rect 8862 7518 8890 7546
rect 8862 7294 8890 7322
rect 8358 6566 8386 6594
rect 10206 7910 10234 7938
rect 9918 7853 9946 7854
rect 9918 7827 9919 7853
rect 9919 7827 9945 7853
rect 9945 7827 9946 7853
rect 9918 7826 9946 7827
rect 9970 7853 9998 7854
rect 9970 7827 9971 7853
rect 9971 7827 9997 7853
rect 9997 7827 9998 7853
rect 9970 7826 9998 7827
rect 10022 7853 10050 7854
rect 10022 7827 10023 7853
rect 10023 7827 10049 7853
rect 10049 7827 10050 7853
rect 10022 7826 10050 7827
rect 10934 10038 10962 10066
rect 11046 10766 11074 10794
rect 11270 10401 11298 10402
rect 11270 10375 11271 10401
rect 11271 10375 11297 10401
rect 11297 10375 11298 10401
rect 11270 10374 11298 10375
rect 11326 10094 11354 10122
rect 11774 11129 11802 11130
rect 11774 11103 11775 11129
rect 11775 11103 11801 11129
rect 11801 11103 11802 11129
rect 11774 11102 11802 11103
rect 11662 10793 11690 10794
rect 11662 10767 11663 10793
rect 11663 10767 11689 10793
rect 11689 10767 11690 10793
rect 11662 10766 11690 10767
rect 11886 11326 11914 11354
rect 12054 11857 12082 11858
rect 12054 11831 12055 11857
rect 12055 11831 12081 11857
rect 12081 11831 12082 11857
rect 12054 11830 12082 11831
rect 12670 11521 12698 11522
rect 12670 11495 12671 11521
rect 12671 11495 12697 11521
rect 12697 11495 12698 11521
rect 12670 11494 12698 11495
rect 13286 11494 13314 11522
rect 14462 12726 14490 12754
rect 14574 12838 14602 12866
rect 14630 12782 14658 12810
rect 14350 12614 14378 12642
rect 14630 12641 14658 12642
rect 14630 12615 14631 12641
rect 14631 12615 14657 12641
rect 14657 12615 14658 12641
rect 14630 12614 14658 12615
rect 14014 12390 14042 12418
rect 17598 12949 17626 12950
rect 17598 12923 17599 12949
rect 17599 12923 17625 12949
rect 17625 12923 17626 12949
rect 17598 12922 17626 12923
rect 17650 12949 17678 12950
rect 17650 12923 17651 12949
rect 17651 12923 17677 12949
rect 17677 12923 17678 12949
rect 17650 12922 17678 12923
rect 17702 12949 17730 12950
rect 17702 12923 17703 12949
rect 17703 12923 17729 12949
rect 17729 12923 17730 12949
rect 17702 12922 17730 12923
rect 20006 13118 20034 13146
rect 19950 12782 19978 12810
rect 18942 12614 18970 12642
rect 18830 12446 18858 12474
rect 20006 12446 20034 12474
rect 14630 12278 14658 12306
rect 14910 12390 14938 12418
rect 15246 12417 15274 12418
rect 15246 12391 15247 12417
rect 15247 12391 15273 12417
rect 15273 12391 15274 12417
rect 15246 12390 15274 12391
rect 18830 12361 18858 12362
rect 18830 12335 18831 12361
rect 18831 12335 18857 12361
rect 18857 12335 18858 12361
rect 18830 12334 18858 12335
rect 17598 12165 17626 12166
rect 17598 12139 17599 12165
rect 17599 12139 17625 12165
rect 17625 12139 17626 12165
rect 17598 12138 17626 12139
rect 17650 12165 17678 12166
rect 17650 12139 17651 12165
rect 17651 12139 17677 12165
rect 17677 12139 17678 12165
rect 17650 12138 17678 12139
rect 17702 12165 17730 12166
rect 17702 12139 17703 12165
rect 17703 12139 17729 12165
rect 17729 12139 17730 12165
rect 17702 12138 17730 12139
rect 20006 12110 20034 12138
rect 12334 11438 12362 11466
rect 11998 11102 12026 11130
rect 12726 11102 12754 11130
rect 11550 10038 11578 10066
rect 10990 9646 11018 9674
rect 10934 9561 10962 9562
rect 10934 9535 10935 9561
rect 10935 9535 10961 9561
rect 10961 9535 10962 9561
rect 10934 9534 10962 9535
rect 11438 9982 11466 10010
rect 11438 9561 11466 9562
rect 11438 9535 11439 9561
rect 11439 9535 11465 9561
rect 11465 9535 11466 9561
rect 11438 9534 11466 9535
rect 11046 9366 11074 9394
rect 10878 9086 10906 9114
rect 10318 8414 10346 8442
rect 11102 8833 11130 8834
rect 11102 8807 11103 8833
rect 11103 8807 11129 8833
rect 11129 8807 11130 8833
rect 11102 8806 11130 8807
rect 11270 9310 11298 9338
rect 11382 9113 11410 9114
rect 11382 9087 11383 9113
rect 11383 9087 11409 9113
rect 11409 9087 11410 9113
rect 11382 9086 11410 9087
rect 11270 8526 11298 8554
rect 11382 8497 11410 8498
rect 11382 8471 11383 8497
rect 11383 8471 11409 8497
rect 11409 8471 11410 8497
rect 11382 8470 11410 8471
rect 10990 8302 11018 8330
rect 10598 8049 10626 8050
rect 10598 8023 10599 8049
rect 10599 8023 10625 8049
rect 10625 8023 10626 8049
rect 10598 8022 10626 8023
rect 9870 7574 9898 7602
rect 9030 7294 9058 7322
rect 9814 7518 9842 7546
rect 10206 7601 10234 7602
rect 10206 7575 10207 7601
rect 10207 7575 10233 7601
rect 10233 7575 10234 7601
rect 10206 7574 10234 7575
rect 10318 7574 10346 7602
rect 10990 8022 11018 8050
rect 10878 7966 10906 7994
rect 10934 7937 10962 7938
rect 10934 7911 10935 7937
rect 10935 7911 10961 7937
rect 10961 7911 10962 7937
rect 10934 7910 10962 7911
rect 10094 7321 10122 7322
rect 10094 7295 10095 7321
rect 10095 7295 10121 7321
rect 10121 7295 10122 7321
rect 10094 7294 10122 7295
rect 9918 7069 9946 7070
rect 9918 7043 9919 7069
rect 9919 7043 9945 7069
rect 9945 7043 9946 7069
rect 9918 7042 9946 7043
rect 9970 7069 9998 7070
rect 9970 7043 9971 7069
rect 9971 7043 9997 7069
rect 9997 7043 9998 7069
rect 9970 7042 9998 7043
rect 10022 7069 10050 7070
rect 10022 7043 10023 7069
rect 10023 7043 10049 7069
rect 10049 7043 10050 7069
rect 10022 7042 10050 7043
rect 9758 6734 9786 6762
rect 8918 6593 8946 6594
rect 8918 6567 8919 6593
rect 8919 6567 8945 6593
rect 8945 6567 8946 6593
rect 8918 6566 8946 6567
rect 9198 6537 9226 6538
rect 9198 6511 9199 6537
rect 9199 6511 9225 6537
rect 9225 6511 9226 6537
rect 9198 6510 9226 6511
rect 9918 6285 9946 6286
rect 9918 6259 9919 6285
rect 9919 6259 9945 6285
rect 9945 6259 9946 6285
rect 9918 6258 9946 6259
rect 9970 6285 9998 6286
rect 9970 6259 9971 6285
rect 9971 6259 9997 6285
rect 9997 6259 9998 6285
rect 9970 6258 9998 6259
rect 10022 6285 10050 6286
rect 10022 6259 10023 6285
rect 10023 6259 10049 6285
rect 10049 6259 10050 6285
rect 10022 6258 10050 6259
rect 10710 6790 10738 6818
rect 2238 5893 2266 5894
rect 2238 5867 2239 5893
rect 2239 5867 2265 5893
rect 2265 5867 2266 5893
rect 2238 5866 2266 5867
rect 2290 5893 2318 5894
rect 2290 5867 2291 5893
rect 2291 5867 2317 5893
rect 2317 5867 2318 5893
rect 2290 5866 2318 5867
rect 2342 5893 2370 5894
rect 2342 5867 2343 5893
rect 2343 5867 2369 5893
rect 2369 5867 2370 5893
rect 2342 5866 2370 5867
rect 2238 5109 2266 5110
rect 2238 5083 2239 5109
rect 2239 5083 2265 5109
rect 2265 5083 2266 5109
rect 2238 5082 2266 5083
rect 2290 5109 2318 5110
rect 2290 5083 2291 5109
rect 2291 5083 2317 5109
rect 2317 5083 2318 5109
rect 2290 5082 2318 5083
rect 2342 5109 2370 5110
rect 2342 5083 2343 5109
rect 2343 5083 2369 5109
rect 2369 5083 2370 5109
rect 2342 5082 2370 5083
rect 2238 4325 2266 4326
rect 2238 4299 2239 4325
rect 2239 4299 2265 4325
rect 2265 4299 2266 4325
rect 2238 4298 2266 4299
rect 2290 4325 2318 4326
rect 2290 4299 2291 4325
rect 2291 4299 2317 4325
rect 2317 4299 2318 4325
rect 2290 4298 2318 4299
rect 2342 4325 2370 4326
rect 2342 4299 2343 4325
rect 2343 4299 2369 4325
rect 2369 4299 2370 4325
rect 2342 4298 2370 4299
rect 9918 5501 9946 5502
rect 9918 5475 9919 5501
rect 9919 5475 9945 5501
rect 9945 5475 9946 5501
rect 9918 5474 9946 5475
rect 9970 5501 9998 5502
rect 9970 5475 9971 5501
rect 9971 5475 9997 5501
rect 9997 5475 9998 5501
rect 9970 5474 9998 5475
rect 10022 5501 10050 5502
rect 10022 5475 10023 5501
rect 10023 5475 10049 5501
rect 10049 5475 10050 5501
rect 10022 5474 10050 5475
rect 9918 4717 9946 4718
rect 9918 4691 9919 4717
rect 9919 4691 9945 4717
rect 9945 4691 9946 4717
rect 9918 4690 9946 4691
rect 9970 4717 9998 4718
rect 9970 4691 9971 4717
rect 9971 4691 9997 4717
rect 9997 4691 9998 4717
rect 9970 4690 9998 4691
rect 10022 4717 10050 4718
rect 10022 4691 10023 4717
rect 10023 4691 10049 4717
rect 10049 4691 10050 4717
rect 10022 4690 10050 4691
rect 2238 3541 2266 3542
rect 2238 3515 2239 3541
rect 2239 3515 2265 3541
rect 2265 3515 2266 3541
rect 2238 3514 2266 3515
rect 2290 3541 2318 3542
rect 2290 3515 2291 3541
rect 2291 3515 2317 3541
rect 2317 3515 2318 3541
rect 2290 3514 2318 3515
rect 2342 3541 2370 3542
rect 2342 3515 2343 3541
rect 2343 3515 2369 3541
rect 2369 3515 2370 3541
rect 2342 3514 2370 3515
rect 2238 2757 2266 2758
rect 2238 2731 2239 2757
rect 2239 2731 2265 2757
rect 2265 2731 2266 2757
rect 2238 2730 2266 2731
rect 2290 2757 2318 2758
rect 2290 2731 2291 2757
rect 2291 2731 2317 2757
rect 2317 2731 2318 2757
rect 2290 2730 2318 2731
rect 2342 2757 2370 2758
rect 2342 2731 2343 2757
rect 2343 2731 2369 2757
rect 2369 2731 2370 2757
rect 2342 2730 2370 2731
rect 2238 1973 2266 1974
rect 2238 1947 2239 1973
rect 2239 1947 2265 1973
rect 2265 1947 2266 1973
rect 2238 1946 2266 1947
rect 2290 1973 2318 1974
rect 2290 1947 2291 1973
rect 2291 1947 2317 1973
rect 2317 1947 2318 1973
rect 2290 1946 2318 1947
rect 2342 1973 2370 1974
rect 2342 1947 2343 1973
rect 2343 1947 2369 1973
rect 2369 1947 2370 1973
rect 2342 1946 2370 1947
rect 9918 3933 9946 3934
rect 9918 3907 9919 3933
rect 9919 3907 9945 3933
rect 9945 3907 9946 3933
rect 9918 3906 9946 3907
rect 9970 3933 9998 3934
rect 9970 3907 9971 3933
rect 9971 3907 9997 3933
rect 9997 3907 9998 3933
rect 9970 3906 9998 3907
rect 10022 3933 10050 3934
rect 10022 3907 10023 3933
rect 10023 3907 10049 3933
rect 10049 3907 10050 3933
rect 10022 3906 10050 3907
rect 9918 3149 9946 3150
rect 9918 3123 9919 3149
rect 9919 3123 9945 3149
rect 9945 3123 9946 3149
rect 9918 3122 9946 3123
rect 9970 3149 9998 3150
rect 9970 3123 9971 3149
rect 9971 3123 9997 3149
rect 9997 3123 9998 3149
rect 9970 3122 9998 3123
rect 10022 3149 10050 3150
rect 10022 3123 10023 3149
rect 10023 3123 10049 3149
rect 10049 3123 10050 3149
rect 10022 3122 10050 3123
rect 9918 2365 9946 2366
rect 9918 2339 9919 2365
rect 9919 2339 9945 2365
rect 9945 2339 9946 2365
rect 9918 2338 9946 2339
rect 9970 2365 9998 2366
rect 9970 2339 9971 2365
rect 9971 2339 9997 2365
rect 9997 2339 9998 2365
rect 9970 2338 9998 2339
rect 10022 2365 10050 2366
rect 10022 2339 10023 2365
rect 10023 2339 10049 2365
rect 10049 2339 10050 2365
rect 10022 2338 10050 2339
rect 11550 9505 11578 9506
rect 11550 9479 11551 9505
rect 11551 9479 11577 9505
rect 11577 9479 11578 9505
rect 11550 9478 11578 9479
rect 11550 9366 11578 9394
rect 11550 8358 11578 8386
rect 11438 8022 11466 8050
rect 10878 7601 10906 7602
rect 10878 7575 10879 7601
rect 10879 7575 10905 7601
rect 10905 7575 10906 7601
rect 10878 7574 10906 7575
rect 10822 6790 10850 6818
rect 11158 6817 11186 6818
rect 11158 6791 11159 6817
rect 11159 6791 11185 6817
rect 11185 6791 11186 6817
rect 11158 6790 11186 6791
rect 11382 6734 11410 6762
rect 10822 6510 10850 6538
rect 11046 6537 11074 6538
rect 11046 6511 11047 6537
rect 11047 6511 11073 6537
rect 11073 6511 11074 6537
rect 11046 6510 11074 6511
rect 11382 6454 11410 6482
rect 11886 9702 11914 9730
rect 11830 9366 11858 9394
rect 11830 9281 11858 9282
rect 11830 9255 11831 9281
rect 11831 9255 11857 9281
rect 11857 9255 11858 9281
rect 11830 9254 11858 9255
rect 11830 9086 11858 9114
rect 13118 11129 13146 11130
rect 13118 11103 13119 11129
rect 13119 11103 13145 11129
rect 13145 11103 13146 11129
rect 13118 11102 13146 11103
rect 13678 11102 13706 11130
rect 12054 10737 12082 10738
rect 12054 10711 12055 10737
rect 12055 10711 12081 10737
rect 12081 10711 12082 10737
rect 12054 10710 12082 10711
rect 12222 10710 12250 10738
rect 12110 10681 12138 10682
rect 12110 10655 12111 10681
rect 12111 10655 12137 10681
rect 12137 10655 12138 10681
rect 12110 10654 12138 10655
rect 12670 10737 12698 10738
rect 12670 10711 12671 10737
rect 12671 10711 12697 10737
rect 12697 10711 12698 10737
rect 12670 10710 12698 10711
rect 12614 10654 12642 10682
rect 12614 10374 12642 10402
rect 12670 10430 12698 10458
rect 12838 10009 12866 10010
rect 12838 9983 12839 10009
rect 12839 9983 12865 10009
rect 12865 9983 12866 10009
rect 12838 9982 12866 9983
rect 12950 9646 12978 9674
rect 13286 9673 13314 9674
rect 13286 9647 13287 9673
rect 13287 9647 13313 9673
rect 13313 9647 13314 9673
rect 13286 9646 13314 9647
rect 12726 9086 12754 9114
rect 12950 9478 12978 9506
rect 13958 11662 13986 11690
rect 18830 11577 18858 11578
rect 18830 11551 18831 11577
rect 18831 11551 18857 11577
rect 18857 11551 18858 11577
rect 18830 11550 18858 11551
rect 20006 11465 20034 11466
rect 20006 11439 20007 11465
rect 20007 11439 20033 11465
rect 20033 11439 20034 11465
rect 20006 11438 20034 11439
rect 17598 11381 17626 11382
rect 17598 11355 17599 11381
rect 17599 11355 17625 11381
rect 17625 11355 17626 11381
rect 17598 11354 17626 11355
rect 17650 11381 17678 11382
rect 17650 11355 17651 11381
rect 17651 11355 17677 11381
rect 17677 11355 17678 11381
rect 17650 11354 17678 11355
rect 17702 11381 17730 11382
rect 17702 11355 17703 11381
rect 17703 11355 17729 11381
rect 17729 11355 17730 11381
rect 17702 11354 17730 11355
rect 14126 11185 14154 11186
rect 14126 11159 14127 11185
rect 14127 11159 14153 11185
rect 14153 11159 14154 11185
rect 14126 11158 14154 11159
rect 14518 11185 14546 11186
rect 14518 11159 14519 11185
rect 14519 11159 14545 11185
rect 14545 11159 14546 11185
rect 14518 11158 14546 11159
rect 18830 11185 18858 11186
rect 18830 11159 18831 11185
rect 18831 11159 18857 11185
rect 18857 11159 18858 11185
rect 18830 11158 18858 11159
rect 13846 11129 13874 11130
rect 13846 11103 13847 11129
rect 13847 11103 13873 11129
rect 13873 11103 13874 11129
rect 13846 11102 13874 11103
rect 14630 11073 14658 11074
rect 14630 11047 14631 11073
rect 14631 11047 14657 11073
rect 14657 11047 14658 11073
rect 14630 11046 14658 11047
rect 20006 11102 20034 11130
rect 14686 10766 14714 10794
rect 14574 10401 14602 10402
rect 14574 10375 14575 10401
rect 14575 10375 14601 10401
rect 14601 10375 14602 10401
rect 14574 10374 14602 10375
rect 15078 11046 15106 11074
rect 17598 10597 17626 10598
rect 17598 10571 17599 10597
rect 17599 10571 17625 10597
rect 17625 10571 17626 10597
rect 17598 10570 17626 10571
rect 17650 10597 17678 10598
rect 17650 10571 17651 10597
rect 17651 10571 17677 10597
rect 17677 10571 17678 10597
rect 17650 10570 17678 10571
rect 17702 10597 17730 10598
rect 17702 10571 17703 10597
rect 17703 10571 17729 10597
rect 17729 10571 17730 10597
rect 17702 10570 17730 10571
rect 14686 10374 14714 10402
rect 15022 10401 15050 10402
rect 15022 10375 15023 10401
rect 15023 10375 15049 10401
rect 15049 10375 15050 10401
rect 15022 10374 15050 10375
rect 14014 10262 14042 10290
rect 14630 10289 14658 10290
rect 14630 10263 14631 10289
rect 14631 10263 14657 10289
rect 14657 10263 14658 10289
rect 14630 10262 14658 10263
rect 13566 9702 13594 9730
rect 11942 8918 11970 8946
rect 12950 8889 12978 8890
rect 12950 8863 12951 8889
rect 12951 8863 12977 8889
rect 12977 8863 12978 8889
rect 12950 8862 12978 8863
rect 13342 8918 13370 8946
rect 13510 8750 13538 8778
rect 13790 9702 13818 9730
rect 14294 9534 14322 9562
rect 13734 8918 13762 8946
rect 13846 8974 13874 9002
rect 14182 9505 14210 9506
rect 14182 9479 14183 9505
rect 14183 9479 14209 9505
rect 14209 9479 14210 9505
rect 14182 9478 14210 9479
rect 15078 10094 15106 10122
rect 18830 10094 18858 10122
rect 17598 9813 17626 9814
rect 17598 9787 17599 9813
rect 17599 9787 17625 9813
rect 17625 9787 17626 9813
rect 17598 9786 17626 9787
rect 17650 9813 17678 9814
rect 17650 9787 17651 9813
rect 17651 9787 17677 9813
rect 17677 9787 17678 9813
rect 17650 9786 17678 9787
rect 17702 9813 17730 9814
rect 17702 9787 17703 9813
rect 17703 9787 17729 9813
rect 17729 9787 17730 9813
rect 17702 9786 17730 9787
rect 19950 10430 19978 10458
rect 20006 10094 20034 10122
rect 18942 9646 18970 9674
rect 14686 9534 14714 9562
rect 14294 9254 14322 9282
rect 14238 9142 14266 9170
rect 14126 8777 14154 8778
rect 14126 8751 14127 8777
rect 14127 8751 14153 8777
rect 14153 8751 14154 8777
rect 14126 8750 14154 8751
rect 14910 9478 14938 9506
rect 14854 9169 14882 9170
rect 14854 9143 14855 9169
rect 14855 9143 14881 9169
rect 14881 9143 14882 9169
rect 14854 9142 14882 9143
rect 17598 9029 17626 9030
rect 17598 9003 17599 9029
rect 17599 9003 17625 9029
rect 17625 9003 17626 9029
rect 17598 9002 17626 9003
rect 17650 9029 17678 9030
rect 17650 9003 17651 9029
rect 17651 9003 17677 9029
rect 17677 9003 17678 9029
rect 17650 9002 17678 9003
rect 17702 9029 17730 9030
rect 17702 9003 17703 9029
rect 17703 9003 17729 9029
rect 17729 9003 17730 9029
rect 17702 9002 17730 9003
rect 18830 8918 18858 8946
rect 18942 9142 18970 9170
rect 14910 8806 14938 8834
rect 11942 8358 11970 8386
rect 11886 7910 11914 7938
rect 12502 8049 12530 8050
rect 12502 8023 12503 8049
rect 12503 8023 12529 8049
rect 12529 8023 12530 8049
rect 12502 8022 12530 8023
rect 11942 7686 11970 7714
rect 12446 7937 12474 7938
rect 12446 7911 12447 7937
rect 12447 7911 12473 7937
rect 12473 7911 12474 7937
rect 12446 7910 12474 7911
rect 13118 7910 13146 7938
rect 12166 7686 12194 7714
rect 11942 6902 11970 6930
rect 12614 6929 12642 6930
rect 12614 6903 12615 6929
rect 12615 6903 12641 6929
rect 12641 6903 12642 6929
rect 12614 6902 12642 6903
rect 12278 6873 12306 6874
rect 12278 6847 12279 6873
rect 12279 6847 12305 6873
rect 12305 6847 12306 6873
rect 12278 6846 12306 6847
rect 11942 6510 11970 6538
rect 11662 6454 11690 6482
rect 11830 6481 11858 6482
rect 11830 6455 11831 6481
rect 11831 6455 11857 6481
rect 11857 6455 11858 6481
rect 11830 6454 11858 6455
rect 10766 6006 10794 6034
rect 11214 6033 11242 6034
rect 11214 6007 11215 6033
rect 11215 6007 11241 6033
rect 11241 6007 11242 6033
rect 11214 6006 11242 6007
rect 12782 6873 12810 6874
rect 12782 6847 12783 6873
rect 12783 6847 12809 6873
rect 12809 6847 12810 6873
rect 12782 6846 12810 6847
rect 13062 6929 13090 6930
rect 13062 6903 13063 6929
rect 13063 6903 13089 6929
rect 13089 6903 13090 6929
rect 13062 6902 13090 6903
rect 12894 6846 12922 6874
rect 18830 8833 18858 8834
rect 18830 8807 18831 8833
rect 18831 8807 18857 8833
rect 18857 8807 18858 8833
rect 18830 8806 18858 8807
rect 20006 9113 20034 9114
rect 20006 9087 20007 9113
rect 20007 9087 20033 9113
rect 20033 9087 20034 9113
rect 20006 9086 20034 9087
rect 20006 8750 20034 8778
rect 20006 8414 20034 8442
rect 17598 8245 17626 8246
rect 17598 8219 17599 8245
rect 17599 8219 17625 8245
rect 17625 8219 17626 8245
rect 17598 8218 17626 8219
rect 17650 8245 17678 8246
rect 17650 8219 17651 8245
rect 17651 8219 17677 8245
rect 17677 8219 17678 8245
rect 17650 8218 17678 8219
rect 17702 8245 17730 8246
rect 17702 8219 17703 8245
rect 17703 8219 17729 8245
rect 17729 8219 17730 8245
rect 17702 8218 17730 8219
rect 17598 7461 17626 7462
rect 17598 7435 17599 7461
rect 17599 7435 17625 7461
rect 17625 7435 17626 7461
rect 17598 7434 17626 7435
rect 17650 7461 17678 7462
rect 17650 7435 17651 7461
rect 17651 7435 17677 7461
rect 17677 7435 17678 7461
rect 17650 7434 17678 7435
rect 17702 7461 17730 7462
rect 17702 7435 17703 7461
rect 17703 7435 17729 7461
rect 17729 7435 17730 7461
rect 17702 7434 17730 7435
rect 13174 6846 13202 6874
rect 14294 6902 14322 6930
rect 13342 6454 13370 6482
rect 10766 2030 10794 2058
rect 8414 1694 8442 1722
rect 9030 1694 9058 1722
rect 9918 1581 9946 1582
rect 9918 1555 9919 1581
rect 9919 1555 9945 1581
rect 9945 1555 9946 1581
rect 9918 1554 9946 1555
rect 9970 1581 9998 1582
rect 9970 1555 9971 1581
rect 9971 1555 9997 1581
rect 9997 1555 9998 1581
rect 9970 1554 9998 1555
rect 10022 1581 10050 1582
rect 10022 1555 10023 1581
rect 10023 1555 10049 1581
rect 10049 1555 10050 1581
rect 10022 1554 10050 1555
rect 11382 2057 11410 2058
rect 11382 2031 11383 2057
rect 11383 2031 11409 2057
rect 11409 2031 11410 2057
rect 11382 2030 11410 2031
rect 12782 2030 12810 2058
rect 12446 1694 12474 1722
rect 13398 2057 13426 2058
rect 13398 2031 13399 2057
rect 13399 2031 13425 2057
rect 13425 2031 13426 2057
rect 13398 2030 13426 2031
rect 13062 1694 13090 1722
rect 13118 1806 13146 1834
rect 17598 6677 17626 6678
rect 17598 6651 17599 6677
rect 17599 6651 17625 6677
rect 17625 6651 17626 6677
rect 17598 6650 17626 6651
rect 17650 6677 17678 6678
rect 17650 6651 17651 6677
rect 17651 6651 17677 6677
rect 17677 6651 17678 6677
rect 17650 6650 17678 6651
rect 17702 6677 17730 6678
rect 17702 6651 17703 6677
rect 17703 6651 17729 6677
rect 17729 6651 17730 6677
rect 17702 6650 17730 6651
rect 17598 5893 17626 5894
rect 17598 5867 17599 5893
rect 17599 5867 17625 5893
rect 17625 5867 17626 5893
rect 17598 5866 17626 5867
rect 17650 5893 17678 5894
rect 17650 5867 17651 5893
rect 17651 5867 17677 5893
rect 17677 5867 17678 5893
rect 17650 5866 17678 5867
rect 17702 5893 17730 5894
rect 17702 5867 17703 5893
rect 17703 5867 17729 5893
rect 17729 5867 17730 5893
rect 17702 5866 17730 5867
rect 17598 5109 17626 5110
rect 17598 5083 17599 5109
rect 17599 5083 17625 5109
rect 17625 5083 17626 5109
rect 17598 5082 17626 5083
rect 17650 5109 17678 5110
rect 17650 5083 17651 5109
rect 17651 5083 17677 5109
rect 17677 5083 17678 5109
rect 17650 5082 17678 5083
rect 17702 5109 17730 5110
rect 17702 5083 17703 5109
rect 17703 5083 17729 5109
rect 17729 5083 17730 5109
rect 17702 5082 17730 5083
rect 17598 4325 17626 4326
rect 17598 4299 17599 4325
rect 17599 4299 17625 4325
rect 17625 4299 17626 4325
rect 17598 4298 17626 4299
rect 17650 4325 17678 4326
rect 17650 4299 17651 4325
rect 17651 4299 17677 4325
rect 17677 4299 17678 4325
rect 17650 4298 17678 4299
rect 17702 4325 17730 4326
rect 17702 4299 17703 4325
rect 17703 4299 17729 4325
rect 17729 4299 17730 4325
rect 17702 4298 17730 4299
rect 17598 3541 17626 3542
rect 17598 3515 17599 3541
rect 17599 3515 17625 3541
rect 17625 3515 17626 3541
rect 17598 3514 17626 3515
rect 17650 3541 17678 3542
rect 17650 3515 17651 3541
rect 17651 3515 17677 3541
rect 17677 3515 17678 3541
rect 17650 3514 17678 3515
rect 17702 3541 17730 3542
rect 17702 3515 17703 3541
rect 17703 3515 17729 3541
rect 17729 3515 17730 3541
rect 17702 3514 17730 3515
rect 17598 2757 17626 2758
rect 17598 2731 17599 2757
rect 17599 2731 17625 2757
rect 17625 2731 17626 2757
rect 17598 2730 17626 2731
rect 17650 2757 17678 2758
rect 17650 2731 17651 2757
rect 17651 2731 17677 2757
rect 17677 2731 17678 2757
rect 17650 2730 17678 2731
rect 17702 2757 17730 2758
rect 17702 2731 17703 2757
rect 17703 2731 17729 2757
rect 17729 2731 17730 2757
rect 17702 2730 17730 2731
rect 17598 1973 17626 1974
rect 17598 1947 17599 1973
rect 17599 1947 17625 1973
rect 17625 1947 17626 1973
rect 17598 1946 17626 1947
rect 17650 1973 17678 1974
rect 17650 1947 17651 1973
rect 17651 1947 17677 1973
rect 17677 1947 17678 1973
rect 17650 1946 17678 1947
rect 17702 1973 17730 1974
rect 17702 1947 17703 1973
rect 17703 1947 17729 1973
rect 17729 1947 17730 1973
rect 17702 1946 17730 1947
rect 14686 1833 14714 1834
rect 14686 1807 14687 1833
rect 14687 1807 14713 1833
rect 14713 1807 14714 1833
rect 14686 1806 14714 1807
<< metal3 >>
rect 2233 19194 2238 19222
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2370 19194 2375 19222
rect 17593 19194 17598 19222
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17730 19194 17735 19222
rect 8745 19110 8750 19138
rect 8778 19110 9310 19138
rect 9338 19110 9343 19138
rect 10089 19110 10094 19138
rect 10122 19110 10878 19138
rect 10906 19110 10911 19138
rect 11769 19110 11774 19138
rect 11802 19110 12782 19138
rect 12810 19110 12815 19138
rect 9913 18802 9918 18830
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 10050 18802 10055 18830
rect 9417 18718 9422 18746
rect 9450 18718 10038 18746
rect 10066 18718 10071 18746
rect 12105 18718 12110 18746
rect 12138 18718 13118 18746
rect 13146 18718 13151 18746
rect 2233 18410 2238 18438
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2370 18410 2375 18438
rect 17593 18410 17598 18438
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17730 18410 17735 18438
rect 9913 18018 9918 18046
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 10050 18018 10055 18046
rect 2233 17626 2238 17654
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2370 17626 2375 17654
rect 17593 17626 17598 17654
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17730 17626 17735 17654
rect 9913 17234 9918 17262
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 10050 17234 10055 17262
rect 2233 16842 2238 16870
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2370 16842 2375 16870
rect 17593 16842 17598 16870
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17730 16842 17735 16870
rect 9913 16450 9918 16478
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 10050 16450 10055 16478
rect 2233 16058 2238 16086
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2370 16058 2375 16086
rect 17593 16058 17598 16086
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17730 16058 17735 16086
rect 9913 15666 9918 15694
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 10050 15666 10055 15694
rect 2233 15274 2238 15302
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2370 15274 2375 15302
rect 17593 15274 17598 15302
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17730 15274 17735 15302
rect 9913 14882 9918 14910
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 10050 14882 10055 14910
rect 2233 14490 2238 14518
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2370 14490 2375 14518
rect 17593 14490 17598 14518
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17730 14490 17735 14518
rect 10929 14238 10934 14266
rect 10962 14238 11830 14266
rect 11858 14238 11863 14266
rect 9913 14098 9918 14126
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 10050 14098 10055 14126
rect 9137 13846 9142 13874
rect 9170 13846 9926 13874
rect 9954 13846 9959 13874
rect 0 13818 400 13832
rect 0 13790 2086 13818
rect 2114 13790 2119 13818
rect 0 13776 400 13790
rect 2233 13706 2238 13734
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2370 13706 2375 13734
rect 17593 13706 17598 13734
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17730 13706 17735 13734
rect 11881 13566 11886 13594
rect 11914 13566 12334 13594
rect 12362 13566 12367 13594
rect 10425 13510 10430 13538
rect 10458 13510 10934 13538
rect 10962 13510 12110 13538
rect 12138 13510 12558 13538
rect 12586 13510 12894 13538
rect 12922 13510 12927 13538
rect 14345 13510 14350 13538
rect 14378 13510 14574 13538
rect 14602 13510 18830 13538
rect 18858 13510 18863 13538
rect 8073 13454 8078 13482
rect 8106 13454 8470 13482
rect 8498 13454 8862 13482
rect 8890 13454 9702 13482
rect 9730 13454 9735 13482
rect 9913 13314 9918 13342
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 10050 13314 10055 13342
rect 10094 13174 10878 13202
rect 10906 13174 10911 13202
rect 10094 13146 10122 13174
rect 20600 13146 21000 13160
rect 9361 13118 9366 13146
rect 9394 13118 10094 13146
rect 10122 13118 10127 13146
rect 10817 13118 10822 13146
rect 10850 13118 11158 13146
rect 11186 13118 11191 13146
rect 11377 13118 11382 13146
rect 11410 13118 11774 13146
rect 11802 13118 11807 13146
rect 20001 13118 20006 13146
rect 20034 13118 21000 13146
rect 20600 13104 21000 13118
rect 8409 13062 8414 13090
rect 8442 13062 9534 13090
rect 9562 13062 9567 13090
rect 2233 12922 2238 12950
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2370 12922 2375 12950
rect 17593 12922 17598 12950
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17730 12922 17735 12950
rect 11433 12838 11438 12866
rect 11466 12838 11942 12866
rect 11970 12838 14070 12866
rect 14098 12838 14574 12866
rect 14602 12838 14607 12866
rect 20600 12810 21000 12824
rect 13729 12782 13734 12810
rect 13762 12782 14630 12810
rect 14658 12782 14663 12810
rect 19945 12782 19950 12810
rect 19978 12782 21000 12810
rect 20600 12768 21000 12782
rect 9702 12726 11970 12754
rect 13281 12726 13286 12754
rect 13314 12726 14462 12754
rect 14490 12726 14495 12754
rect 9702 12642 9730 12726
rect 11942 12698 11970 12726
rect 9865 12670 9870 12698
rect 9898 12670 10318 12698
rect 10346 12670 10654 12698
rect 10682 12670 10687 12698
rect 11942 12670 13566 12698
rect 13594 12670 13599 12698
rect 9697 12614 9702 12642
rect 9730 12614 9735 12642
rect 9814 12614 9926 12642
rect 9954 12614 9959 12642
rect 13225 12614 13230 12642
rect 13258 12614 13454 12642
rect 13482 12614 13678 12642
rect 13706 12614 13711 12642
rect 14345 12614 14350 12642
rect 14378 12614 14630 12642
rect 14658 12614 18942 12642
rect 18970 12614 18975 12642
rect 9814 12586 9842 12614
rect 9081 12558 9086 12586
rect 9114 12558 9842 12586
rect 9913 12530 9918 12558
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 10050 12530 10055 12558
rect 20600 12474 21000 12488
rect 8409 12446 8414 12474
rect 8442 12446 9142 12474
rect 9170 12446 9175 12474
rect 9641 12446 9646 12474
rect 9674 12446 10038 12474
rect 10066 12446 10430 12474
rect 10458 12446 10654 12474
rect 10682 12446 10687 12474
rect 15946 12446 18830 12474
rect 18858 12446 18863 12474
rect 20001 12446 20006 12474
rect 20034 12446 21000 12474
rect 15946 12418 15974 12446
rect 20600 12432 21000 12446
rect 10257 12390 10262 12418
rect 10290 12390 10710 12418
rect 10738 12390 10743 12418
rect 14009 12390 14014 12418
rect 14042 12390 14910 12418
rect 14938 12390 14943 12418
rect 15241 12390 15246 12418
rect 15274 12390 15974 12418
rect 14910 12362 14938 12390
rect 2137 12334 2142 12362
rect 2170 12334 6902 12362
rect 6930 12334 6935 12362
rect 7177 12334 7182 12362
rect 7210 12334 8302 12362
rect 8330 12334 8750 12362
rect 8778 12334 8783 12362
rect 10089 12334 10094 12362
rect 10122 12334 10878 12362
rect 10906 12334 11270 12362
rect 11298 12334 11303 12362
rect 14910 12334 18830 12362
rect 18858 12334 18863 12362
rect 6902 12306 6930 12334
rect 6902 12278 8638 12306
rect 8666 12278 8671 12306
rect 12945 12278 12950 12306
rect 12978 12278 13398 12306
rect 13426 12278 14630 12306
rect 14658 12278 14663 12306
rect 961 12222 966 12250
rect 994 12222 999 12250
rect 0 12138 400 12152
rect 966 12138 994 12222
rect 2233 12138 2238 12166
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2370 12138 2375 12166
rect 17593 12138 17598 12166
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17730 12138 17735 12166
rect 20600 12138 21000 12152
rect 0 12110 994 12138
rect 20001 12110 20006 12138
rect 20034 12110 21000 12138
rect 0 12096 400 12110
rect 20600 12096 21000 12110
rect 8913 11942 8918 11970
rect 8946 11942 10094 11970
rect 10122 11942 10127 11970
rect 9193 11886 9198 11914
rect 9226 11886 9310 11914
rect 9338 11886 9758 11914
rect 9786 11886 9791 11914
rect 9921 11886 9926 11914
rect 9954 11886 10598 11914
rect 10626 11886 10631 11914
rect 8073 11830 8078 11858
rect 8106 11830 8918 11858
rect 8946 11830 8951 11858
rect 11657 11830 11662 11858
rect 11690 11830 12054 11858
rect 12082 11830 12087 11858
rect 0 11802 400 11816
rect 0 11774 966 11802
rect 994 11774 999 11802
rect 0 11760 400 11774
rect 9913 11746 9918 11774
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 10050 11746 10055 11774
rect 7681 11718 7686 11746
rect 7714 11718 7910 11746
rect 7938 11718 8302 11746
rect 8330 11718 9198 11746
rect 9226 11718 9231 11746
rect 6785 11662 6790 11690
rect 6818 11662 7574 11690
rect 7602 11662 7607 11690
rect 9081 11662 9086 11690
rect 9114 11662 9534 11690
rect 9562 11662 9567 11690
rect 9641 11662 9646 11690
rect 9674 11662 13958 11690
rect 13986 11662 13991 11690
rect 7625 11606 7630 11634
rect 7658 11606 8358 11634
rect 8386 11606 9590 11634
rect 9618 11606 9623 11634
rect 4186 11550 5670 11578
rect 5698 11550 7406 11578
rect 7434 11550 7439 11578
rect 10355 11550 10374 11578
rect 10402 11550 10407 11578
rect 15946 11550 18830 11578
rect 18858 11550 18863 11578
rect 4186 11522 4214 11550
rect 2137 11494 2142 11522
rect 2170 11494 4214 11522
rect 10929 11494 10934 11522
rect 10962 11494 12670 11522
rect 12698 11494 13286 11522
rect 13314 11494 13319 11522
rect 15946 11466 15974 11550
rect 20600 11466 21000 11480
rect 9361 11438 9366 11466
rect 9394 11438 9702 11466
rect 9730 11438 10430 11466
rect 10458 11438 10463 11466
rect 12329 11438 12334 11466
rect 12362 11438 15974 11466
rect 20001 11438 20006 11466
rect 20034 11438 21000 11466
rect 20600 11424 21000 11438
rect 7546 11382 7966 11410
rect 7994 11382 11830 11410
rect 11858 11382 11863 11410
rect 2233 11354 2238 11382
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2370 11354 2375 11382
rect 7513 11326 7518 11354
rect 7546 11326 7574 11382
rect 17593 11354 17598 11382
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17730 11354 17735 11382
rect 9417 11326 9422 11354
rect 9450 11326 10262 11354
rect 10290 11326 11886 11354
rect 11914 11326 11919 11354
rect 8297 11270 8302 11298
rect 8330 11270 9086 11298
rect 9114 11270 9119 11298
rect 10075 11270 10094 11298
rect 10122 11270 10127 11298
rect 10201 11270 10206 11298
rect 10234 11270 10822 11298
rect 10850 11270 10855 11298
rect 8801 11214 8806 11242
rect 8834 11214 9198 11242
rect 9226 11214 9231 11242
rect 9473 11214 9478 11242
rect 9506 11214 9814 11242
rect 9842 11214 9982 11242
rect 10010 11214 10015 11242
rect 9305 11158 9310 11186
rect 9338 11158 9926 11186
rect 9954 11158 9959 11186
rect 10089 11158 10094 11186
rect 10122 11158 10710 11186
rect 10738 11158 10743 11186
rect 14121 11158 14126 11186
rect 14154 11158 14518 11186
rect 14546 11158 14551 11186
rect 15946 11158 18830 11186
rect 18858 11158 18863 11186
rect 9977 11102 9982 11130
rect 10010 11102 10654 11130
rect 10682 11102 10990 11130
rect 11018 11102 11023 11130
rect 11769 11102 11774 11130
rect 11802 11102 11998 11130
rect 12026 11102 12726 11130
rect 12754 11102 12759 11130
rect 13113 11102 13118 11130
rect 13146 11102 13678 11130
rect 13706 11102 13846 11130
rect 13874 11102 13879 11130
rect 11774 11074 11802 11102
rect 15946 11074 15974 11158
rect 20600 11130 21000 11144
rect 20001 11102 20006 11130
rect 20034 11102 21000 11130
rect 20600 11088 21000 11102
rect 10817 11046 10822 11074
rect 10850 11046 11802 11074
rect 14625 11046 14630 11074
rect 14658 11046 15078 11074
rect 15106 11046 15974 11074
rect 9913 10962 9918 10990
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 10050 10962 10055 10990
rect 7681 10878 7686 10906
rect 7714 10878 8918 10906
rect 8946 10878 10094 10906
rect 10122 10878 10127 10906
rect 10257 10878 10262 10906
rect 10290 10878 10374 10906
rect 10402 10878 10407 10906
rect 8129 10822 8134 10850
rect 8162 10822 8414 10850
rect 8442 10822 10346 10850
rect 10318 10794 10346 10822
rect 6449 10766 6454 10794
rect 6482 10766 7294 10794
rect 7322 10766 7327 10794
rect 8017 10766 8022 10794
rect 8050 10766 9086 10794
rect 9114 10766 9119 10794
rect 10313 10766 10318 10794
rect 10346 10766 10486 10794
rect 10514 10766 10710 10794
rect 10738 10766 10743 10794
rect 11041 10766 11046 10794
rect 11074 10766 11662 10794
rect 11690 10766 14686 10794
rect 14714 10766 14719 10794
rect 8465 10710 8470 10738
rect 8498 10710 8974 10738
rect 9002 10710 12054 10738
rect 12082 10710 12087 10738
rect 12217 10710 12222 10738
rect 12250 10710 12670 10738
rect 12698 10710 12703 10738
rect 12105 10654 12110 10682
rect 12138 10654 12614 10682
rect 12642 10654 12647 10682
rect 2233 10570 2238 10598
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2370 10570 2375 10598
rect 17593 10570 17598 10598
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17730 10570 17735 10598
rect 20600 10458 21000 10472
rect 7233 10430 7238 10458
rect 7266 10430 7742 10458
rect 7770 10430 7775 10458
rect 10873 10430 10878 10458
rect 10906 10430 12670 10458
rect 12698 10430 12703 10458
rect 19945 10430 19950 10458
rect 19978 10430 21000 10458
rect 20600 10416 21000 10430
rect 6505 10374 6510 10402
rect 6538 10374 6790 10402
rect 6818 10374 6823 10402
rect 10033 10374 10038 10402
rect 10066 10374 11270 10402
rect 11298 10374 11303 10402
rect 12609 10374 12614 10402
rect 12642 10374 14574 10402
rect 14602 10374 14607 10402
rect 14681 10374 14686 10402
rect 14714 10374 15022 10402
rect 15050 10374 15055 10402
rect 5385 10318 5390 10346
rect 5418 10318 7294 10346
rect 7322 10318 8078 10346
rect 8106 10318 10430 10346
rect 10458 10318 10463 10346
rect 10089 10262 10094 10290
rect 10122 10262 10822 10290
rect 10850 10262 10855 10290
rect 14009 10262 14014 10290
rect 14042 10262 14630 10290
rect 14658 10262 14663 10290
rect 9913 10178 9918 10206
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 10050 10178 10055 10206
rect 6953 10150 6958 10178
rect 6986 10150 7490 10178
rect 7462 10122 7490 10150
rect 20600 10122 21000 10136
rect 5049 10094 5054 10122
rect 5082 10094 6902 10122
rect 6930 10094 6935 10122
rect 7457 10094 7462 10122
rect 7490 10094 8022 10122
rect 8050 10094 8055 10122
rect 8745 10094 8750 10122
rect 8778 10094 9254 10122
rect 9282 10094 11326 10122
rect 11354 10094 11359 10122
rect 15073 10094 15078 10122
rect 15106 10094 18830 10122
rect 18858 10094 18863 10122
rect 20001 10094 20006 10122
rect 20034 10094 21000 10122
rect 20600 10080 21000 10094
rect 10817 10038 10822 10066
rect 10850 10038 10934 10066
rect 10962 10038 11550 10066
rect 11578 10038 11583 10066
rect 5385 9982 5390 10010
rect 5418 9982 6734 10010
rect 6762 9982 6767 10010
rect 7546 9982 8806 10010
rect 8834 9982 9422 10010
rect 9450 9982 9455 10010
rect 11433 9982 11438 10010
rect 11466 9982 12838 10010
rect 12866 9982 12871 10010
rect 7546 9954 7574 9982
rect 2081 9926 2086 9954
rect 2114 9926 7574 9954
rect 8241 9926 8246 9954
rect 8274 9926 8526 9954
rect 8554 9926 9702 9954
rect 9730 9926 9735 9954
rect 2233 9786 2238 9814
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2370 9786 2375 9814
rect 17593 9786 17598 9814
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17730 9786 17735 9814
rect 8297 9702 8302 9730
rect 8330 9702 8414 9730
rect 8442 9702 9310 9730
rect 9338 9702 9646 9730
rect 9674 9702 10374 9730
rect 10402 9702 10407 9730
rect 11881 9702 11886 9730
rect 11914 9702 13566 9730
rect 13594 9702 13790 9730
rect 13818 9702 13823 9730
rect 10145 9646 10150 9674
rect 10178 9646 10654 9674
rect 10682 9646 10990 9674
rect 11018 9646 11023 9674
rect 12945 9646 12950 9674
rect 12978 9646 13286 9674
rect 13314 9646 18942 9674
rect 18970 9646 18975 9674
rect 7289 9590 7294 9618
rect 7322 9590 10206 9618
rect 10234 9590 10239 9618
rect 10929 9534 10934 9562
rect 10962 9534 11438 9562
rect 11466 9534 11471 9562
rect 14289 9534 14294 9562
rect 14322 9534 14686 9562
rect 14714 9534 14719 9562
rect 7401 9478 7406 9506
rect 7434 9478 9534 9506
rect 9562 9478 10542 9506
rect 10570 9478 10575 9506
rect 11545 9478 11550 9506
rect 11578 9478 12950 9506
rect 12978 9478 12983 9506
rect 14177 9478 14182 9506
rect 14210 9478 14910 9506
rect 14938 9478 14943 9506
rect 9913 9394 9918 9422
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 10050 9394 10055 9422
rect 6729 9366 6734 9394
rect 6762 9366 7126 9394
rect 7154 9366 7574 9394
rect 9025 9366 9030 9394
rect 9058 9366 9534 9394
rect 9562 9366 9702 9394
rect 9730 9366 9735 9394
rect 11041 9366 11046 9394
rect 11074 9366 11550 9394
rect 11578 9366 11830 9394
rect 11858 9366 11863 9394
rect 7546 9338 7574 9366
rect 7546 9310 9814 9338
rect 9842 9310 10598 9338
rect 10626 9310 10631 9338
rect 11265 9310 11270 9338
rect 11298 9310 13454 9338
rect 13426 9282 13454 9310
rect 7457 9254 7462 9282
rect 7490 9254 8862 9282
rect 8890 9254 8974 9282
rect 9002 9254 9007 9282
rect 9865 9254 9870 9282
rect 9898 9254 10206 9282
rect 10234 9254 10239 9282
rect 10761 9254 10766 9282
rect 10794 9254 11830 9282
rect 11858 9254 11863 9282
rect 13426 9254 14294 9282
rect 14322 9254 14327 9282
rect 8185 9198 8190 9226
rect 8218 9198 9198 9226
rect 9226 9198 9231 9226
rect 9305 9198 9310 9226
rect 9338 9198 9814 9226
rect 9842 9198 9847 9226
rect 7905 9142 7910 9170
rect 7938 9142 8358 9170
rect 8386 9142 8638 9170
rect 8666 9142 8671 9170
rect 10649 9142 10654 9170
rect 10682 9142 11410 9170
rect 14233 9142 14238 9170
rect 14266 9142 14854 9170
rect 14882 9142 18942 9170
rect 18970 9142 18975 9170
rect 11382 9114 11410 9142
rect 20600 9114 21000 9128
rect 7569 9086 7574 9114
rect 7602 9086 10878 9114
rect 10906 9086 10911 9114
rect 11377 9086 11382 9114
rect 11410 9086 11830 9114
rect 11858 9086 12726 9114
rect 12754 9086 12759 9114
rect 20001 9086 20006 9114
rect 20034 9086 21000 9114
rect 20600 9072 21000 9086
rect 2233 9002 2238 9030
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2370 9002 2375 9030
rect 17593 9002 17598 9030
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17730 9002 17735 9030
rect 9473 8974 9478 9002
rect 9506 8974 13846 9002
rect 13874 8974 13879 9002
rect 8689 8918 8694 8946
rect 8722 8918 9590 8946
rect 9618 8918 9623 8946
rect 11937 8918 11942 8946
rect 11970 8918 13342 8946
rect 13370 8918 13734 8946
rect 13762 8918 13767 8946
rect 15946 8918 18830 8946
rect 18858 8918 18863 8946
rect 15946 8890 15974 8918
rect 961 8862 966 8890
rect 994 8862 999 8890
rect 7345 8862 7350 8890
rect 7378 8862 9758 8890
rect 9786 8862 9791 8890
rect 12945 8862 12950 8890
rect 12978 8862 15974 8890
rect 0 8778 400 8792
rect 966 8778 994 8862
rect 2137 8806 2142 8834
rect 2170 8806 4998 8834
rect 5026 8806 5031 8834
rect 6393 8806 6398 8834
rect 6426 8806 6734 8834
rect 6762 8806 6767 8834
rect 9193 8806 9198 8834
rect 9226 8806 9478 8834
rect 9506 8806 9511 8834
rect 9921 8806 9926 8834
rect 9954 8806 11102 8834
rect 11130 8806 11135 8834
rect 14905 8806 14910 8834
rect 14938 8806 18830 8834
rect 18858 8806 18863 8834
rect 20600 8778 21000 8792
rect 0 8750 994 8778
rect 7401 8750 7406 8778
rect 7434 8750 8582 8778
rect 8610 8750 10206 8778
rect 10234 8750 10239 8778
rect 13505 8750 13510 8778
rect 13538 8750 14126 8778
rect 14154 8750 14159 8778
rect 20001 8750 20006 8778
rect 20034 8750 21000 8778
rect 0 8736 400 8750
rect 20600 8736 21000 8750
rect 5777 8694 5782 8722
rect 5810 8694 7126 8722
rect 7154 8694 7159 8722
rect 9913 8610 9918 8638
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 10050 8610 10055 8638
rect 7546 8526 7854 8554
rect 7882 8526 7887 8554
rect 8745 8526 8750 8554
rect 8778 8526 11270 8554
rect 11298 8526 11303 8554
rect 7546 8498 7574 8526
rect 7121 8470 7126 8498
rect 7154 8470 7574 8498
rect 8409 8470 8414 8498
rect 8442 8470 9198 8498
rect 9226 8470 9231 8498
rect 10257 8470 10262 8498
rect 10290 8470 11382 8498
rect 11410 8470 11415 8498
rect 20600 8442 21000 8456
rect 4993 8414 4998 8442
rect 5026 8414 7070 8442
rect 7098 8414 7103 8442
rect 9534 8414 10318 8442
rect 10346 8414 10351 8442
rect 20001 8414 20006 8442
rect 20034 8414 21000 8442
rect 9534 8386 9562 8414
rect 20600 8400 21000 8414
rect 9193 8358 9198 8386
rect 9226 8358 9534 8386
rect 9562 8358 9567 8386
rect 11545 8358 11550 8386
rect 11578 8358 11942 8386
rect 11970 8358 11975 8386
rect 10201 8302 10206 8330
rect 10234 8302 10990 8330
rect 11018 8302 11023 8330
rect 2233 8218 2238 8246
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2370 8218 2375 8246
rect 17593 8218 17598 8246
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17730 8218 17735 8246
rect 0 8106 400 8120
rect 0 8078 966 8106
rect 994 8078 999 8106
rect 0 8064 400 8078
rect 9697 8022 9702 8050
rect 9730 8022 10598 8050
rect 10626 8022 10631 8050
rect 10985 8022 10990 8050
rect 11018 8022 11438 8050
rect 11466 8022 12502 8050
rect 12530 8022 12535 8050
rect 7177 7966 7182 7994
rect 7210 7966 7686 7994
rect 7714 7966 10878 7994
rect 10906 7966 10911 7994
rect 6393 7910 6398 7938
rect 6426 7910 7070 7938
rect 7098 7910 7103 7938
rect 9585 7910 9590 7938
rect 9618 7910 10206 7938
rect 10234 7910 10239 7938
rect 10929 7910 10934 7938
rect 10962 7910 11886 7938
rect 11914 7910 11919 7938
rect 12441 7910 12446 7938
rect 12474 7910 13118 7938
rect 13146 7910 13151 7938
rect 9913 7826 9918 7854
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 10050 7826 10055 7854
rect 5329 7742 5334 7770
rect 5362 7742 6790 7770
rect 6818 7742 6823 7770
rect 11937 7686 11942 7714
rect 11970 7686 12166 7714
rect 12194 7686 12199 7714
rect 2137 7574 2142 7602
rect 2170 7574 5334 7602
rect 5362 7574 5367 7602
rect 9865 7574 9870 7602
rect 9898 7574 10206 7602
rect 10234 7574 10239 7602
rect 10313 7574 10318 7602
rect 10346 7574 10878 7602
rect 10906 7574 10911 7602
rect 8465 7518 8470 7546
rect 8498 7518 8862 7546
rect 8890 7518 9814 7546
rect 9842 7518 9847 7546
rect 2233 7434 2238 7462
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2370 7434 2375 7462
rect 17593 7434 17598 7462
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17730 7434 17735 7462
rect 7009 7294 7014 7322
rect 7042 7294 7294 7322
rect 7322 7294 8246 7322
rect 8274 7294 8862 7322
rect 8890 7294 9030 7322
rect 9058 7294 10094 7322
rect 10122 7294 10127 7322
rect 9913 7042 9918 7070
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 10050 7042 10055 7070
rect 11937 6902 11942 6930
rect 11970 6902 12614 6930
rect 12642 6902 12647 6930
rect 13057 6902 13062 6930
rect 13090 6902 14294 6930
rect 14322 6902 14327 6930
rect 12273 6846 12278 6874
rect 12306 6846 12782 6874
rect 12810 6846 12815 6874
rect 12889 6846 12894 6874
rect 12922 6846 13174 6874
rect 13202 6846 13207 6874
rect 10705 6790 10710 6818
rect 10738 6790 10822 6818
rect 10850 6790 11158 6818
rect 11186 6790 11191 6818
rect 9753 6734 9758 6762
rect 9786 6734 11382 6762
rect 11410 6734 11415 6762
rect 2233 6650 2238 6678
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2370 6650 2375 6678
rect 17593 6650 17598 6678
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17730 6650 17735 6678
rect 8353 6566 8358 6594
rect 8386 6566 8918 6594
rect 8946 6566 8951 6594
rect 9193 6510 9198 6538
rect 9226 6510 10822 6538
rect 10850 6510 11046 6538
rect 11074 6510 11942 6538
rect 11970 6510 11975 6538
rect 11377 6454 11382 6482
rect 11410 6454 11662 6482
rect 11690 6454 11830 6482
rect 11858 6454 13342 6482
rect 13370 6454 13375 6482
rect 9913 6258 9918 6286
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 10050 6258 10055 6286
rect 10761 6006 10766 6034
rect 10794 6006 11214 6034
rect 11242 6006 11247 6034
rect 2233 5866 2238 5894
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2370 5866 2375 5894
rect 17593 5866 17598 5894
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17730 5866 17735 5894
rect 9913 5474 9918 5502
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 10050 5474 10055 5502
rect 2233 5082 2238 5110
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2370 5082 2375 5110
rect 17593 5082 17598 5110
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17730 5082 17735 5110
rect 9913 4690 9918 4718
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 10050 4690 10055 4718
rect 2233 4298 2238 4326
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2370 4298 2375 4326
rect 17593 4298 17598 4326
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17730 4298 17735 4326
rect 9913 3906 9918 3934
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 10050 3906 10055 3934
rect 2233 3514 2238 3542
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2370 3514 2375 3542
rect 17593 3514 17598 3542
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17730 3514 17735 3542
rect 9913 3122 9918 3150
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 10050 3122 10055 3150
rect 2233 2730 2238 2758
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2370 2730 2375 2758
rect 17593 2730 17598 2758
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17730 2730 17735 2758
rect 9913 2338 9918 2366
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 10050 2338 10055 2366
rect 10761 2030 10766 2058
rect 10794 2030 11382 2058
rect 11410 2030 11415 2058
rect 12777 2030 12782 2058
rect 12810 2030 13398 2058
rect 13426 2030 13431 2058
rect 2233 1946 2238 1974
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2370 1946 2375 1974
rect 17593 1946 17598 1974
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17730 1946 17735 1974
rect 13113 1806 13118 1834
rect 13146 1806 14686 1834
rect 14714 1806 14719 1834
rect 8409 1694 8414 1722
rect 8442 1694 9030 1722
rect 9058 1694 9063 1722
rect 12441 1694 12446 1722
rect 12474 1694 13062 1722
rect 13090 1694 13095 1722
rect 9913 1554 9918 1582
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 10050 1554 10055 1582
<< via3 >>
rect 2238 19194 2266 19222
rect 2290 19194 2318 19222
rect 2342 19194 2370 19222
rect 17598 19194 17626 19222
rect 17650 19194 17678 19222
rect 17702 19194 17730 19222
rect 9918 18802 9946 18830
rect 9970 18802 9998 18830
rect 10022 18802 10050 18830
rect 2238 18410 2266 18438
rect 2290 18410 2318 18438
rect 2342 18410 2370 18438
rect 17598 18410 17626 18438
rect 17650 18410 17678 18438
rect 17702 18410 17730 18438
rect 9918 18018 9946 18046
rect 9970 18018 9998 18046
rect 10022 18018 10050 18046
rect 2238 17626 2266 17654
rect 2290 17626 2318 17654
rect 2342 17626 2370 17654
rect 17598 17626 17626 17654
rect 17650 17626 17678 17654
rect 17702 17626 17730 17654
rect 9918 17234 9946 17262
rect 9970 17234 9998 17262
rect 10022 17234 10050 17262
rect 2238 16842 2266 16870
rect 2290 16842 2318 16870
rect 2342 16842 2370 16870
rect 17598 16842 17626 16870
rect 17650 16842 17678 16870
rect 17702 16842 17730 16870
rect 9918 16450 9946 16478
rect 9970 16450 9998 16478
rect 10022 16450 10050 16478
rect 2238 16058 2266 16086
rect 2290 16058 2318 16086
rect 2342 16058 2370 16086
rect 17598 16058 17626 16086
rect 17650 16058 17678 16086
rect 17702 16058 17730 16086
rect 9918 15666 9946 15694
rect 9970 15666 9998 15694
rect 10022 15666 10050 15694
rect 2238 15274 2266 15302
rect 2290 15274 2318 15302
rect 2342 15274 2370 15302
rect 17598 15274 17626 15302
rect 17650 15274 17678 15302
rect 17702 15274 17730 15302
rect 9918 14882 9946 14910
rect 9970 14882 9998 14910
rect 10022 14882 10050 14910
rect 2238 14490 2266 14518
rect 2290 14490 2318 14518
rect 2342 14490 2370 14518
rect 17598 14490 17626 14518
rect 17650 14490 17678 14518
rect 17702 14490 17730 14518
rect 9918 14098 9946 14126
rect 9970 14098 9998 14126
rect 10022 14098 10050 14126
rect 2238 13706 2266 13734
rect 2290 13706 2318 13734
rect 2342 13706 2370 13734
rect 17598 13706 17626 13734
rect 17650 13706 17678 13734
rect 17702 13706 17730 13734
rect 9918 13314 9946 13342
rect 9970 13314 9998 13342
rect 10022 13314 10050 13342
rect 2238 12922 2266 12950
rect 2290 12922 2318 12950
rect 2342 12922 2370 12950
rect 17598 12922 17626 12950
rect 17650 12922 17678 12950
rect 17702 12922 17730 12950
rect 9918 12530 9946 12558
rect 9970 12530 9998 12558
rect 10022 12530 10050 12558
rect 2238 12138 2266 12166
rect 2290 12138 2318 12166
rect 2342 12138 2370 12166
rect 17598 12138 17626 12166
rect 17650 12138 17678 12166
rect 17702 12138 17730 12166
rect 9918 11746 9946 11774
rect 9970 11746 9998 11774
rect 10022 11746 10050 11774
rect 10374 11550 10402 11578
rect 2238 11354 2266 11382
rect 2290 11354 2318 11382
rect 2342 11354 2370 11382
rect 17598 11354 17626 11382
rect 17650 11354 17678 11382
rect 17702 11354 17730 11382
rect 10094 11270 10122 11298
rect 9918 10962 9946 10990
rect 9970 10962 9998 10990
rect 10022 10962 10050 10990
rect 10094 10878 10122 10906
rect 10374 10878 10402 10906
rect 2238 10570 2266 10598
rect 2290 10570 2318 10598
rect 2342 10570 2370 10598
rect 17598 10570 17626 10598
rect 17650 10570 17678 10598
rect 17702 10570 17730 10598
rect 9918 10178 9946 10206
rect 9970 10178 9998 10206
rect 10022 10178 10050 10206
rect 2238 9786 2266 9814
rect 2290 9786 2318 9814
rect 2342 9786 2370 9814
rect 17598 9786 17626 9814
rect 17650 9786 17678 9814
rect 17702 9786 17730 9814
rect 9918 9394 9946 9422
rect 9970 9394 9998 9422
rect 10022 9394 10050 9422
rect 2238 9002 2266 9030
rect 2290 9002 2318 9030
rect 2342 9002 2370 9030
rect 17598 9002 17626 9030
rect 17650 9002 17678 9030
rect 17702 9002 17730 9030
rect 9918 8610 9946 8638
rect 9970 8610 9998 8638
rect 10022 8610 10050 8638
rect 2238 8218 2266 8246
rect 2290 8218 2318 8246
rect 2342 8218 2370 8246
rect 17598 8218 17626 8246
rect 17650 8218 17678 8246
rect 17702 8218 17730 8246
rect 9918 7826 9946 7854
rect 9970 7826 9998 7854
rect 10022 7826 10050 7854
rect 2238 7434 2266 7462
rect 2290 7434 2318 7462
rect 2342 7434 2370 7462
rect 17598 7434 17626 7462
rect 17650 7434 17678 7462
rect 17702 7434 17730 7462
rect 9918 7042 9946 7070
rect 9970 7042 9998 7070
rect 10022 7042 10050 7070
rect 2238 6650 2266 6678
rect 2290 6650 2318 6678
rect 2342 6650 2370 6678
rect 17598 6650 17626 6678
rect 17650 6650 17678 6678
rect 17702 6650 17730 6678
rect 9918 6258 9946 6286
rect 9970 6258 9998 6286
rect 10022 6258 10050 6286
rect 2238 5866 2266 5894
rect 2290 5866 2318 5894
rect 2342 5866 2370 5894
rect 17598 5866 17626 5894
rect 17650 5866 17678 5894
rect 17702 5866 17730 5894
rect 9918 5474 9946 5502
rect 9970 5474 9998 5502
rect 10022 5474 10050 5502
rect 2238 5082 2266 5110
rect 2290 5082 2318 5110
rect 2342 5082 2370 5110
rect 17598 5082 17626 5110
rect 17650 5082 17678 5110
rect 17702 5082 17730 5110
rect 9918 4690 9946 4718
rect 9970 4690 9998 4718
rect 10022 4690 10050 4718
rect 2238 4298 2266 4326
rect 2290 4298 2318 4326
rect 2342 4298 2370 4326
rect 17598 4298 17626 4326
rect 17650 4298 17678 4326
rect 17702 4298 17730 4326
rect 9918 3906 9946 3934
rect 9970 3906 9998 3934
rect 10022 3906 10050 3934
rect 2238 3514 2266 3542
rect 2290 3514 2318 3542
rect 2342 3514 2370 3542
rect 17598 3514 17626 3542
rect 17650 3514 17678 3542
rect 17702 3514 17730 3542
rect 9918 3122 9946 3150
rect 9970 3122 9998 3150
rect 10022 3122 10050 3150
rect 2238 2730 2266 2758
rect 2290 2730 2318 2758
rect 2342 2730 2370 2758
rect 17598 2730 17626 2758
rect 17650 2730 17678 2758
rect 17702 2730 17730 2758
rect 9918 2338 9946 2366
rect 9970 2338 9998 2366
rect 10022 2338 10050 2366
rect 2238 1946 2266 1974
rect 2290 1946 2318 1974
rect 2342 1946 2370 1974
rect 17598 1946 17626 1974
rect 17650 1946 17678 1974
rect 17702 1946 17730 1974
rect 9918 1554 9946 1582
rect 9970 1554 9998 1582
rect 10022 1554 10050 1582
<< metal4 >>
rect 2224 19222 2384 19238
rect 2224 19194 2238 19222
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2370 19194 2384 19222
rect 2224 18438 2384 19194
rect 2224 18410 2238 18438
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2370 18410 2384 18438
rect 2224 17654 2384 18410
rect 2224 17626 2238 17654
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2370 17626 2384 17654
rect 2224 16870 2384 17626
rect 2224 16842 2238 16870
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2370 16842 2384 16870
rect 2224 16086 2384 16842
rect 2224 16058 2238 16086
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2370 16058 2384 16086
rect 2224 15302 2384 16058
rect 2224 15274 2238 15302
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2370 15274 2384 15302
rect 2224 14518 2384 15274
rect 2224 14490 2238 14518
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2370 14490 2384 14518
rect 2224 13734 2384 14490
rect 2224 13706 2238 13734
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2370 13706 2384 13734
rect 2224 12950 2384 13706
rect 2224 12922 2238 12950
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2370 12922 2384 12950
rect 2224 12166 2384 12922
rect 2224 12138 2238 12166
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2370 12138 2384 12166
rect 2224 11382 2384 12138
rect 2224 11354 2238 11382
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2370 11354 2384 11382
rect 2224 10598 2384 11354
rect 2224 10570 2238 10598
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2370 10570 2384 10598
rect 2224 9814 2384 10570
rect 2224 9786 2238 9814
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2370 9786 2384 9814
rect 2224 9030 2384 9786
rect 2224 9002 2238 9030
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2370 9002 2384 9030
rect 2224 8246 2384 9002
rect 2224 8218 2238 8246
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2370 8218 2384 8246
rect 2224 7462 2384 8218
rect 2224 7434 2238 7462
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2370 7434 2384 7462
rect 2224 6678 2384 7434
rect 2224 6650 2238 6678
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2370 6650 2384 6678
rect 2224 5894 2384 6650
rect 2224 5866 2238 5894
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2370 5866 2384 5894
rect 2224 5110 2384 5866
rect 2224 5082 2238 5110
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2370 5082 2384 5110
rect 2224 4326 2384 5082
rect 2224 4298 2238 4326
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2370 4298 2384 4326
rect 2224 3542 2384 4298
rect 2224 3514 2238 3542
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2370 3514 2384 3542
rect 2224 2758 2384 3514
rect 2224 2730 2238 2758
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2370 2730 2384 2758
rect 2224 1974 2384 2730
rect 2224 1946 2238 1974
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2370 1946 2384 1974
rect 2224 1538 2384 1946
rect 9904 18830 10064 19238
rect 9904 18802 9918 18830
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 10050 18802 10064 18830
rect 9904 18046 10064 18802
rect 9904 18018 9918 18046
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 10050 18018 10064 18046
rect 9904 17262 10064 18018
rect 9904 17234 9918 17262
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 10050 17234 10064 17262
rect 9904 16478 10064 17234
rect 9904 16450 9918 16478
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 10050 16450 10064 16478
rect 9904 15694 10064 16450
rect 9904 15666 9918 15694
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 10050 15666 10064 15694
rect 9904 14910 10064 15666
rect 9904 14882 9918 14910
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 10050 14882 10064 14910
rect 9904 14126 10064 14882
rect 9904 14098 9918 14126
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 10050 14098 10064 14126
rect 9904 13342 10064 14098
rect 9904 13314 9918 13342
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 10050 13314 10064 13342
rect 9904 12558 10064 13314
rect 9904 12530 9918 12558
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 10050 12530 10064 12558
rect 9904 11774 10064 12530
rect 9904 11746 9918 11774
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 10050 11746 10064 11774
rect 9904 10990 10064 11746
rect 17584 19222 17744 19238
rect 17584 19194 17598 19222
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17730 19194 17744 19222
rect 17584 18438 17744 19194
rect 17584 18410 17598 18438
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17730 18410 17744 18438
rect 17584 17654 17744 18410
rect 17584 17626 17598 17654
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17730 17626 17744 17654
rect 17584 16870 17744 17626
rect 17584 16842 17598 16870
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17730 16842 17744 16870
rect 17584 16086 17744 16842
rect 17584 16058 17598 16086
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17730 16058 17744 16086
rect 17584 15302 17744 16058
rect 17584 15274 17598 15302
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17730 15274 17744 15302
rect 17584 14518 17744 15274
rect 17584 14490 17598 14518
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17730 14490 17744 14518
rect 17584 13734 17744 14490
rect 17584 13706 17598 13734
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17730 13706 17744 13734
rect 17584 12950 17744 13706
rect 17584 12922 17598 12950
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17730 12922 17744 12950
rect 17584 12166 17744 12922
rect 17584 12138 17598 12166
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17730 12138 17744 12166
rect 10374 11578 10402 11583
rect 9904 10962 9918 10990
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 10050 10962 10064 10990
rect 9904 10206 10064 10962
rect 10094 11298 10122 11303
rect 10094 10906 10122 11270
rect 10094 10873 10122 10878
rect 10374 10906 10402 11550
rect 10374 10873 10402 10878
rect 17584 11382 17744 12138
rect 17584 11354 17598 11382
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17730 11354 17744 11382
rect 9904 10178 9918 10206
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 10050 10178 10064 10206
rect 9904 9422 10064 10178
rect 9904 9394 9918 9422
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 10050 9394 10064 9422
rect 9904 8638 10064 9394
rect 9904 8610 9918 8638
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 10050 8610 10064 8638
rect 9904 7854 10064 8610
rect 9904 7826 9918 7854
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 10050 7826 10064 7854
rect 9904 7070 10064 7826
rect 9904 7042 9918 7070
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 10050 7042 10064 7070
rect 9904 6286 10064 7042
rect 9904 6258 9918 6286
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 10050 6258 10064 6286
rect 9904 5502 10064 6258
rect 9904 5474 9918 5502
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 10050 5474 10064 5502
rect 9904 4718 10064 5474
rect 9904 4690 9918 4718
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 10050 4690 10064 4718
rect 9904 3934 10064 4690
rect 9904 3906 9918 3934
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 10050 3906 10064 3934
rect 9904 3150 10064 3906
rect 9904 3122 9918 3150
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 10050 3122 10064 3150
rect 9904 2366 10064 3122
rect 9904 2338 9918 2366
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 10050 2338 10064 2366
rect 9904 1582 10064 2338
rect 9904 1554 9918 1582
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 10050 1554 10064 1582
rect 9904 1538 10064 1554
rect 17584 10598 17744 11354
rect 17584 10570 17598 10598
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17730 10570 17744 10598
rect 17584 9814 17744 10570
rect 17584 9786 17598 9814
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17730 9786 17744 9814
rect 17584 9030 17744 9786
rect 17584 9002 17598 9030
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17730 9002 17744 9030
rect 17584 8246 17744 9002
rect 17584 8218 17598 8246
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17730 8218 17744 8246
rect 17584 7462 17744 8218
rect 17584 7434 17598 7462
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17730 7434 17744 7462
rect 17584 6678 17744 7434
rect 17584 6650 17598 6678
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17730 6650 17744 6678
rect 17584 5894 17744 6650
rect 17584 5866 17598 5894
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17730 5866 17744 5894
rect 17584 5110 17744 5866
rect 17584 5082 17598 5110
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17730 5082 17744 5110
rect 17584 4326 17744 5082
rect 17584 4298 17598 4326
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17730 4298 17744 4326
rect 17584 3542 17744 4298
rect 17584 3514 17598 3542
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17730 3514 17744 3542
rect 17584 2758 17744 3514
rect 17584 2730 17598 2758
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17730 2730 17744 2758
rect 17584 1974 17744 2730
rect 17584 1946 17598 1974
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17730 1946 17744 1974
rect 17584 1538 17744 1946
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _115_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8624 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _116_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 11480 0 -1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _117_
timestamp 1698175906
transform 1 0 10584 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _118_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 6944 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _119_
timestamp 1698175906
transform -1 0 7560 0 1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _120_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 6720 0 1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _121_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8064 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _122_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 9352 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _123_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 8512 0 -1 10192
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _124_
timestamp 1698175906
transform 1 0 11984 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _125_
timestamp 1698175906
transform -1 0 10360 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _126_
timestamp 1698175906
transform -1 0 11200 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _127_
timestamp 1698175906
transform 1 0 9016 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _128_
timestamp 1698175906
transform 1 0 9016 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _129_
timestamp 1698175906
transform 1 0 10248 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _130_
timestamp 1698175906
transform -1 0 10472 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _131_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 11536 0 -1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _132_
timestamp 1698175906
transform 1 0 7896 0 -1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _133_
timestamp 1698175906
transform -1 0 11144 0 -1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _134_
timestamp 1698175906
transform 1 0 10472 0 -1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _135_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 11032 0 1 10192
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _136_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 12544 0 -1 10192
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _137_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 12544 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _138_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10808 0 -1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _139_
timestamp 1698175906
transform 1 0 11536 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _140_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 9072 0 1 6272
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _141_
timestamp 1698175906
transform 1 0 7280 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _142_
timestamp 1698175906
transform -1 0 9352 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _143_
timestamp 1698175906
transform -1 0 8512 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _144_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8792 0 1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _145_
timestamp 1698175906
transform -1 0 8512 0 -1 7056
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _146_
timestamp 1698175906
transform 1 0 8456 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _147_
timestamp 1698175906
transform 1 0 9744 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _148_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 9912 0 -1 8624
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _149_
timestamp 1698175906
transform 1 0 7224 0 1 9408
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _150_
timestamp 1698175906
transform 1 0 7336 0 -1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _151_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 6104 0 -1 10976
box -43 -43 715 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _152_
timestamp 1698175906
transform 1 0 6552 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _153_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10584 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _154_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10528 0 -1 7840
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _155_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 10416 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _156_
timestamp 1698175906
transform 1 0 8680 0 -1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _157_
timestamp 1698175906
transform 1 0 7224 0 -1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _158_
timestamp 1698175906
transform -1 0 8512 0 -1 10976
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _159_
timestamp 1698175906
transform -1 0 8008 0 -1 8624
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _160_
timestamp 1698175906
transform -1 0 7840 0 1 7840
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _161_
timestamp 1698175906
transform 1 0 11032 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _162_
timestamp 1698175906
transform 1 0 8624 0 -1 8624
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _163_
timestamp 1698175906
transform -1 0 8904 0 -1 7840
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _164_
timestamp 1698175906
transform 1 0 8848 0 -1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _165_
timestamp 1698175906
transform -1 0 10920 0 1 6272
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _166_
timestamp 1698175906
transform -1 0 10864 0 1 7056
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _167_
timestamp 1698175906
transform -1 0 10472 0 1 10976
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _168_
timestamp 1698175906
transform 1 0 11928 0 1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _169_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 11984 0 1 10976
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _170_
timestamp 1698175906
transform -1 0 6944 0 1 7840
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _171_
timestamp 1698175906
transform -1 0 10248 0 1 8624
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _172_
timestamp 1698175906
transform 1 0 6944 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _173_
timestamp 1698175906
transform -1 0 14392 0 1 8624
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _174_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 10808 0 -1 10976
box -43 -43 771 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _175_
timestamp 1698175906
transform 1 0 11312 0 -1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _176_
timestamp 1698175906
transform -1 0 13664 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _177_
timestamp 1698175906
transform 1 0 14952 0 1 10192
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _178_
timestamp 1698175906
transform 1 0 14504 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _179_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 7336 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _180_
timestamp 1698175906
transform -1 0 7784 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _181_
timestamp 1698175906
transform 1 0 6888 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _182_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 7000 0 1 8624
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _183_
timestamp 1698175906
transform 1 0 5656 0 -1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _184_
timestamp 1698175906
transform -1 0 11760 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _185_
timestamp 1698175906
transform 1 0 11648 0 -1 9408
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _186_
timestamp 1698175906
transform 1 0 12544 0 -1 7056
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _187_
timestamp 1698175906
transform -1 0 12376 0 -1 7056
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _188_
timestamp 1698175906
transform -1 0 12600 0 1 7840
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _189_
timestamp 1698175906
transform 1 0 10584 0 1 7840
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _190_
timestamp 1698175906
transform 1 0 11872 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _191_
timestamp 1698175906
transform 1 0 8680 0 1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _192_
timestamp 1698175906
transform -1 0 14336 0 1 9408
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _193_
timestamp 1698175906
transform -1 0 14112 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _194_
timestamp 1698175906
transform 1 0 12880 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _195_
timestamp 1698175906
transform -1 0 14784 0 1 10976
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _196_
timestamp 1698175906
transform 1 0 13776 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _197_
timestamp 1698175906
transform 1 0 8960 0 1 10976
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _198_
timestamp 1698175906
transform 1 0 7336 0 -1 11760
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _199_
timestamp 1698175906
transform -1 0 6888 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _200_
timestamp 1698175906
transform -1 0 10192 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _201_
timestamp 1698175906
transform 1 0 11200 0 -1 12544
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _202_
timestamp 1698175906
transform -1 0 14728 0 -1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _203_
timestamp 1698175906
transform -1 0 13384 0 1 12544
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _204_
timestamp 1698175906
transform 1 0 14504 0 1 12544
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _205_
timestamp 1698175906
transform -1 0 13776 0 1 12544
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _206_
timestamp 1698175906
transform -1 0 14168 0 1 12544
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _207_
timestamp 1698175906
transform -1 0 14000 0 1 11760
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _208_
timestamp 1698175906
transform -1 0 10976 0 -1 12544
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _209_
timestamp 1698175906
transform 1 0 10808 0 1 14112
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _210_
timestamp 1698175906
transform 1 0 10304 0 -1 11760
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _211_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 10080 0 -1 10976
box -43 -43 883 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _212_
timestamp 1698175906
transform 1 0 10248 0 -1 12544
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _213_
timestamp 1698175906
transform 1 0 9128 0 1 12544
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _214_
timestamp 1698175906
transform 1 0 10528 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _215_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8904 0 -1 12544
box -43 -43 659 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _216_
timestamp 1698175906
transform -1 0 8512 0 1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _217_
timestamp 1698175906
transform -1 0 9968 0 -1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _218_
timestamp 1698175906
transform -1 0 9968 0 1 12544
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _219_
timestamp 1698175906
transform -1 0 9688 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _220_
timestamp 1698175906
transform -1 0 10304 0 1 14112
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _221_
timestamp 1698175906
transform 1 0 9912 0 -1 11760
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _222_
timestamp 1698175906
transform -1 0 10360 0 1 11760
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _223_
timestamp 1698175906
transform 1 0 9800 0 1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _224_
timestamp 1698175906
transform -1 0 9800 0 -1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _225_
timestamp 1698175906
transform 1 0 8680 0 1 11760
box -43 -43 659 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _226_
timestamp 1698175906
transform -1 0 8176 0 1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _227_
timestamp 1698175906
transform 1 0 10584 0 1 12544
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _228_
timestamp 1698175906
transform -1 0 12040 0 -1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _229_
timestamp 1698175906
transform -1 0 11424 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _230_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 11760 0 1 9408
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _231_
timestamp 1698175906
transform 1 0 7168 0 1 6272
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _232_
timestamp 1698175906
transform 1 0 9632 0 -1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _233_
timestamp 1698175906
transform 1 0 4928 0 1 10192
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _234_
timestamp 1698175906
transform 1 0 4928 0 -1 10192
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _235_
timestamp 1698175906
transform 1 0 6888 0 -1 7840
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _236_
timestamp 1698175906
transform 1 0 8120 0 1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _237_
timestamp 1698175906
transform 1 0 9688 0 -1 6272
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _238_
timestamp 1698175906
transform 1 0 10808 0 -1 11760
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _239_
timestamp 1698175906
transform -1 0 6888 0 -1 7840
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _240_
timestamp 1698175906
transform 1 0 13328 0 -1 9408
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _241_
timestamp 1698175906
transform 1 0 13552 0 -1 10192
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _242_
timestamp 1698175906
transform -1 0 6552 0 1 8624
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _243_
timestamp 1698175906
transform 1 0 11424 0 1 8624
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _244_
timestamp 1698175906
transform 1 0 11760 0 1 6272
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _245_
timestamp 1698175906
transform 1 0 11592 0 1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _246_
timestamp 1698175906
transform 1 0 13384 0 -1 8624
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _247_
timestamp 1698175906
transform 1 0 13552 0 -1 10976
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _248_
timestamp 1698175906
transform -1 0 7224 0 -1 11760
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _249_
timestamp 1698175906
transform 1 0 12768 0 1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _250_
timestamp 1698175906
transform 1 0 12824 0 -1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _251_
timestamp 1698175906
transform 1 0 13384 0 -1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _252_
timestamp 1698175906
transform 1 0 10304 0 -1 14112
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _253_
timestamp 1698175906
transform 1 0 7112 0 1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _254_
timestamp 1698175906
transform 1 0 7952 0 1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _255_
timestamp 1698175906
transform 1 0 8680 0 -1 14112
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _256_
timestamp 1698175906
transform -1 0 8456 0 -1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _257_
timestamp 1698175906
transform 1 0 10808 0 1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _258_
timestamp 1698175906
transform 1 0 15008 0 -1 12544
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _259_
timestamp 1698175906
transform 1 0 12824 0 -1 7056
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__140__A2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9184 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__165__A2
timestamp 1698175906
transform 1 0 11032 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__186__A2
timestamp 1698175906
transform 1 0 11984 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__198__B1
timestamp 1698175906
transform 1 0 7952 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__230__CLK
timestamp 1698175906
transform 1 0 13496 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__231__CLK
timestamp 1698175906
transform -1 0 8904 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__232__CLK
timestamp 1698175906
transform 1 0 11368 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__233__CLK
timestamp 1698175906
transform 1 0 6888 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__234__CLK
timestamp 1698175906
transform 1 0 6776 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__235__CLK
timestamp 1698175906
transform 1 0 9016 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__236__CLK
timestamp 1698175906
transform 1 0 10080 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__237__CLK
timestamp 1698175906
transform 1 0 11424 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__238__CLK
timestamp 1698175906
transform 1 0 12656 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__239__CLK
timestamp 1698175906
transform 1 0 6888 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__240__CLK
timestamp 1698175906
transform 1 0 13216 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__241__CLK
timestamp 1698175906
transform 1 0 13440 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__242__CLK
timestamp 1698175906
transform 1 0 6776 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__243__CLK
timestamp 1698175906
transform 1 0 13048 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__244__CLK
timestamp 1698175906
transform 1 0 13496 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__245__CLK
timestamp 1698175906
transform 1 0 13328 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__246__CLK
timestamp 1698175906
transform 1 0 13272 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__247__CLK
timestamp 1698175906
transform 1 0 13440 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__248__CLK
timestamp 1698175906
transform 1 0 7224 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__249__CLK
timestamp 1698175906
transform 1 0 14616 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__250__CLK
timestamp 1698175906
transform 1 0 14840 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__251__CLK
timestamp 1698175906
transform 1 0 13272 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__252__CLK
timestamp 1698175906
transform -1 0 12152 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__253__CLK
timestamp 1698175906
transform 1 0 8848 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__254__CLK
timestamp 1698175906
transform 1 0 9688 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__255__CLK
timestamp 1698175906
transform -1 0 8512 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__256__CLK
timestamp 1698175906
transform 1 0 8736 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__257__CLK
timestamp 1698175906
transform 1 0 12544 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1698175906
transform 1 0 8792 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9352 0 -1 10192
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1698175906
transform -1 0 10360 0 1 10192
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1698175906
transform 1 0 11200 0 1 10192
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 784 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698175906
transform 1 0 2688 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698175906
transform 1 0 4592 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698175906
transform 1 0 6496 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_138 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8400 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_165 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9912 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_169
timestamp 1698175906
transform 1 0 10136 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_172
timestamp 1698175906
transform 1 0 10304 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_176 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10528 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_206
timestamp 1698175906
transform 1 0 12208 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_210
timestamp 1698175906
transform 1 0 12432 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_237
timestamp 1698175906
transform 1 0 13944 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_266
timestamp 1698175906
transform 1 0 15568 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_270
timestamp 1698175906
transform 1 0 15792 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_274
timestamp 1698175906
transform 1 0 16016 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_308
timestamp 1698175906
transform 1 0 17920 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_342
timestamp 1698175906
transform 1 0 19824 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_346
timestamp 1698175906
transform 1 0 20048 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_348
timestamp 1698175906
transform 1 0 20160 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 784 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698175906
transform 1 0 4368 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698175906
transform 1 0 4704 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698175906
transform 1 0 8288 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_142
timestamp 1698175906
transform 1 0 8624 0 -1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_174
timestamp 1698175906
transform 1 0 10416 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_178
timestamp 1698175906
transform 1 0 10640 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_180
timestamp 1698175906
transform 1 0 10752 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_207
timestamp 1698175906
transform 1 0 12264 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_209
timestamp 1698175906
transform 1 0 12376 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_212
timestamp 1698175906
transform 1 0 12544 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_216
timestamp 1698175906
transform 1 0 12768 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_243
timestamp 1698175906
transform 1 0 14280 0 -1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_275
timestamp 1698175906
transform 1 0 16072 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_279
timestamp 1698175906
transform 1 0 16296 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_282
timestamp 1698175906
transform 1 0 16464 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_346
timestamp 1698175906
transform 1 0 20048 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_348
timestamp 1698175906
transform 1 0 20160 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698175906
transform 1 0 784 0 1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698175906
transform 1 0 2576 0 1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698175906
transform 1 0 2744 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698175906
transform 1 0 6328 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_107
timestamp 1698175906
transform 1 0 6664 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_171
timestamp 1698175906
transform 1 0 10248 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_177
timestamp 1698175906
transform 1 0 10584 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_241
timestamp 1698175906
transform 1 0 14168 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698175906
transform 1 0 14504 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698175906
transform 1 0 18088 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_317
timestamp 1698175906
transform 1 0 18424 0 1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698175906
transform 1 0 784 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698175906
transform 1 0 4368 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698175906
transform 1 0 4704 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698175906
transform 1 0 8288 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_142
timestamp 1698175906
transform 1 0 8624 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_206
timestamp 1698175906
transform 1 0 12208 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_212
timestamp 1698175906
transform 1 0 12544 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_276
timestamp 1698175906
transform 1 0 16128 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_282
timestamp 1698175906
transform 1 0 16464 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_346
timestamp 1698175906
transform 1 0 20048 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_348
timestamp 1698175906
transform 1 0 20160 0 -1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698175906
transform 1 0 784 0 1 3136
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698175906
transform 1 0 2576 0 1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698175906
transform 1 0 2744 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698175906
transform 1 0 6328 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_107
timestamp 1698175906
transform 1 0 6664 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698175906
transform 1 0 10248 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_177
timestamp 1698175906
transform 1 0 10584 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_241
timestamp 1698175906
transform 1 0 14168 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698175906
transform 1 0 14504 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698175906
transform 1 0 18088 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_317
timestamp 1698175906
transform 1 0 18424 0 1 3136
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698175906
transform 1 0 784 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698175906
transform 1 0 4368 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698175906
transform 1 0 4704 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698175906
transform 1 0 8288 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_142
timestamp 1698175906
transform 1 0 8624 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_206
timestamp 1698175906
transform 1 0 12208 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_212
timestamp 1698175906
transform 1 0 12544 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698175906
transform 1 0 16128 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_282
timestamp 1698175906
transform 1 0 16464 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_346
timestamp 1698175906
transform 1 0 20048 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_348
timestamp 1698175906
transform 1 0 20160 0 -1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698175906
transform 1 0 784 0 1 3920
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698175906
transform 1 0 2576 0 1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698175906
transform 1 0 2744 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698175906
transform 1 0 6328 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_107
timestamp 1698175906
transform 1 0 6664 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_171
timestamp 1698175906
transform 1 0 10248 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_177
timestamp 1698175906
transform 1 0 10584 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_241
timestamp 1698175906
transform 1 0 14168 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_247
timestamp 1698175906
transform 1 0 14504 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_311
timestamp 1698175906
transform 1 0 18088 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_317
timestamp 1698175906
transform 1 0 18424 0 1 3920
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698175906
transform 1 0 784 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698175906
transform 1 0 4368 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_72
timestamp 1698175906
transform 1 0 4704 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698175906
transform 1 0 8288 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_142
timestamp 1698175906
transform 1 0 8624 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_206
timestamp 1698175906
transform 1 0 12208 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_212
timestamp 1698175906
transform 1 0 12544 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_276
timestamp 1698175906
transform 1 0 16128 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_282
timestamp 1698175906
transform 1 0 16464 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_346
timestamp 1698175906
transform 1 0 20048 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_348
timestamp 1698175906
transform 1 0 20160 0 -1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698175906
transform 1 0 784 0 1 4704
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698175906
transform 1 0 2576 0 1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_37
timestamp 1698175906
transform 1 0 2744 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_101
timestamp 1698175906
transform 1 0 6328 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_107
timestamp 1698175906
transform 1 0 6664 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_171
timestamp 1698175906
transform 1 0 10248 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_177
timestamp 1698175906
transform 1 0 10584 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_241
timestamp 1698175906
transform 1 0 14168 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_247
timestamp 1698175906
transform 1 0 14504 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_311
timestamp 1698175906
transform 1 0 18088 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_317
timestamp 1698175906
transform 1 0 18424 0 1 4704
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698175906
transform 1 0 784 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698175906
transform 1 0 4368 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_72
timestamp 1698175906
transform 1 0 4704 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_136
timestamp 1698175906
transform 1 0 8288 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_142
timestamp 1698175906
transform 1 0 8624 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_206
timestamp 1698175906
transform 1 0 12208 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_212
timestamp 1698175906
transform 1 0 12544 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_276
timestamp 1698175906
transform 1 0 16128 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_282
timestamp 1698175906
transform 1 0 16464 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_346
timestamp 1698175906
transform 1 0 20048 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_348
timestamp 1698175906
transform 1 0 20160 0 -1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698175906
transform 1 0 784 0 1 5488
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698175906
transform 1 0 2576 0 1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_37
timestamp 1698175906
transform 1 0 2744 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698175906
transform 1 0 6328 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_107
timestamp 1698175906
transform 1 0 6664 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_171
timestamp 1698175906
transform 1 0 10248 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_177
timestamp 1698175906
transform 1 0 10584 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_241
timestamp 1698175906
transform 1 0 14168 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_247
timestamp 1698175906
transform 1 0 14504 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_311
timestamp 1698175906
transform 1 0 18088 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_317
timestamp 1698175906
transform 1 0 18424 0 1 5488
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2
timestamp 1698175906
transform 1 0 784 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698175906
transform 1 0 4368 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_72
timestamp 1698175906
transform 1 0 4704 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698175906
transform 1 0 8288 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_142
timestamp 1698175906
transform 1 0 8624 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_144
timestamp 1698175906
transform 1 0 8736 0 -1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_147 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8904 0 -1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_155
timestamp 1698175906
transform 1 0 9352 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_159
timestamp 1698175906
transform 1 0 9576 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_190
timestamp 1698175906
transform 1 0 11312 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_194 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 11536 0 -1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_212
timestamp 1698175906
transform 1 0 12544 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_276
timestamp 1698175906
transform 1 0 16128 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_282
timestamp 1698175906
transform 1 0 16464 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_346
timestamp 1698175906
transform 1 0 20048 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_348
timestamp 1698175906
transform 1 0 20160 0 -1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698175906
transform 1 0 784 0 1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698175906
transform 1 0 2576 0 1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_37
timestamp 1698175906
transform 1 0 2744 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698175906
transform 1 0 6328 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_107
timestamp 1698175906
transform 1 0 6664 0 1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_115
timestamp 1698175906
transform 1 0 7112 0 1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_150
timestamp 1698175906
transform 1 0 9072 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_154
timestamp 1698175906
transform 1 0 9296 0 1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_170
timestamp 1698175906
transform 1 0 10192 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_174
timestamp 1698175906
transform 1 0 10416 0 1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_177
timestamp 1698175906
transform 1 0 10584 0 1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_183
timestamp 1698175906
transform 1 0 10920 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_187
timestamp 1698175906
transform 1 0 11144 0 1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_195
timestamp 1698175906
transform 1 0 11592 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_197
timestamp 1698175906
transform 1 0 11704 0 1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_227
timestamp 1698175906
transform 1 0 13384 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_231
timestamp 1698175906
transform 1 0 13608 0 1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_239
timestamp 1698175906
transform 1 0 14056 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_243
timestamp 1698175906
transform 1 0 14280 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_247
timestamp 1698175906
transform 1 0 14504 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_311
timestamp 1698175906
transform 1 0 18088 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_317
timestamp 1698175906
transform 1 0 18424 0 1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_2
timestamp 1698175906
transform 1 0 784 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_66
timestamp 1698175906
transform 1 0 4368 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_72
timestamp 1698175906
transform 1 0 4704 0 -1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_104
timestamp 1698175906
transform 1 0 6496 0 -1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_120
timestamp 1698175906
transform 1 0 7392 0 -1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_128
timestamp 1698175906
transform 1 0 7840 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_132
timestamp 1698175906
transform 1 0 8064 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_134
timestamp 1698175906
transform 1 0 8176 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_142
timestamp 1698175906
transform 1 0 8624 0 -1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_158
timestamp 1698175906
transform 1 0 9520 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_189
timestamp 1698175906
transform 1 0 11256 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_193
timestamp 1698175906
transform 1 0 11480 0 -1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_201
timestamp 1698175906
transform 1 0 11928 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_209
timestamp 1698175906
transform 1 0 12376 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_223
timestamp 1698175906
transform 1 0 13160 0 -1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_255
timestamp 1698175906
transform 1 0 14952 0 -1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_271
timestamp 1698175906
transform 1 0 15848 0 -1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_279
timestamp 1698175906
transform 1 0 16296 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_282
timestamp 1698175906
transform 1 0 16464 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_346
timestamp 1698175906
transform 1 0 20048 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_348
timestamp 1698175906
transform 1 0 20160 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698175906
transform 1 0 784 0 1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698175906
transform 1 0 2576 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_37
timestamp 1698175906
transform 1 0 2744 0 1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_101
timestamp 1698175906
transform 1 0 6328 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_107
timestamp 1698175906
transform 1 0 6664 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_113
timestamp 1698175906
transform 1 0 7000 0 1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_129
timestamp 1698175906
transform 1 0 7896 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_166
timestamp 1698175906
transform 1 0 9968 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_170
timestamp 1698175906
transform 1 0 10192 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_174
timestamp 1698175906
transform 1 0 10416 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_182
timestamp 1698175906
transform 1 0 10864 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_190
timestamp 1698175906
transform 1 0 11312 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_194
timestamp 1698175906
transform 1 0 11536 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_224
timestamp 1698175906
transform 1 0 13216 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_228
timestamp 1698175906
transform 1 0 13440 0 1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_244
timestamp 1698175906
transform 1 0 14336 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_247
timestamp 1698175906
transform 1 0 14504 0 1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_311
timestamp 1698175906
transform 1 0 18088 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_317
timestamp 1698175906
transform 1 0 18424 0 1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_2
timestamp 1698175906
transform 1 0 784 0 -1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_66
timestamp 1698175906
transform 1 0 4368 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_72
timestamp 1698175906
transform 1 0 4704 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_80
timestamp 1698175906
transform 1 0 5152 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_147
timestamp 1698175906
transform 1 0 8904 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_151
timestamp 1698175906
transform 1 0 9128 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_159
timestamp 1698175906
transform 1 0 9576 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_163
timestamp 1698175906
transform 1 0 9800 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_165
timestamp 1698175906
transform 1 0 9912 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_174
timestamp 1698175906
transform 1 0 10416 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_185
timestamp 1698175906
transform 1 0 11032 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_193
timestamp 1698175906
transform 1 0 11480 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_197
timestamp 1698175906
transform 1 0 11704 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_199
timestamp 1698175906
transform 1 0 11816 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_208
timestamp 1698175906
transform 1 0 12320 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_212
timestamp 1698175906
transform 1 0 12544 0 -1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_276
timestamp 1698175906
transform 1 0 16128 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_282
timestamp 1698175906
transform 1 0 16464 0 -1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_346
timestamp 1698175906
transform 1 0 20048 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_348
timestamp 1698175906
transform 1 0 20160 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_2
timestamp 1698175906
transform 1 0 784 0 1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698175906
transform 1 0 2576 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_37
timestamp 1698175906
transform 1 0 2744 0 1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_101
timestamp 1698175906
transform 1 0 6328 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_120
timestamp 1698175906
transform 1 0 7392 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_122
timestamp 1698175906
transform 1 0 7504 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_128
timestamp 1698175906
transform 1 0 7840 0 1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_160
timestamp 1698175906
transform 1 0 9632 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_164
timestamp 1698175906
transform 1 0 9856 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_173
timestamp 1698175906
transform 1 0 10360 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_184
timestamp 1698175906
transform 1 0 10976 0 1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_200
timestamp 1698175906
transform 1 0 11872 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_213
timestamp 1698175906
transform 1 0 12600 0 1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_247
timestamp 1698175906
transform 1 0 14504 0 1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_311
timestamp 1698175906
transform 1 0 18088 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_317
timestamp 1698175906
transform 1 0 18424 0 1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_28
timestamp 1698175906
transform 1 0 2240 0 -1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_60
timestamp 1698175906
transform 1 0 4032 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_68
timestamp 1698175906
transform 1 0 4480 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_72
timestamp 1698175906
transform 1 0 4704 0 -1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_88
timestamp 1698175906
transform 1 0 5600 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_95
timestamp 1698175906
transform 1 0 5992 0 -1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_125
timestamp 1698175906
transform 1 0 7672 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_131
timestamp 1698175906
transform 1 0 8008 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_139
timestamp 1698175906
transform 1 0 8456 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_165
timestamp 1698175906
transform 1 0 9912 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_187
timestamp 1698175906
transform 1 0 11144 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_189
timestamp 1698175906
transform 1 0 11256 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_196
timestamp 1698175906
transform 1 0 11648 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_204
timestamp 1698175906
transform 1 0 12096 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_208
timestamp 1698175906
transform 1 0 12320 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_212
timestamp 1698175906
transform 1 0 12544 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_220
timestamp 1698175906
transform 1 0 12992 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_223
timestamp 1698175906
transform 1 0 13160 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_256
timestamp 1698175906
transform 1 0 15008 0 -1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_272
timestamp 1698175906
transform 1 0 15904 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_282
timestamp 1698175906
transform 1 0 16464 0 -1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_314
timestamp 1698175906
transform 1 0 18256 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_322
timestamp 1698175906
transform 1 0 18704 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_28
timestamp 1698175906
transform 1 0 2240 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_32
timestamp 1698175906
transform 1 0 2464 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698175906
transform 1 0 2576 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_37
timestamp 1698175906
transform 1 0 2744 0 1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_69
timestamp 1698175906
transform 1 0 4536 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_73
timestamp 1698175906
transform 1 0 4760 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_75
timestamp 1698175906
transform 1 0 4872 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_107
timestamp 1698175906
transform 1 0 6664 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_111
timestamp 1698175906
transform 1 0 6888 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_123
timestamp 1698175906
transform 1 0 7560 0 1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_191
timestamp 1698175906
transform 1 0 11368 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_221
timestamp 1698175906
transform 1 0 13048 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_223
timestamp 1698175906
transform 1 0 13160 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_247
timestamp 1698175906
transform 1 0 14504 0 1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_311
timestamp 1698175906
transform 1 0 18088 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_317
timestamp 1698175906
transform 1 0 18424 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_321
timestamp 1698175906
transform 1 0 18648 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_2
timestamp 1698175906
transform 1 0 784 0 -1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_66
timestamp 1698175906
transform 1 0 4368 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_72
timestamp 1698175906
transform 1 0 4704 0 -1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_104
timestamp 1698175906
transform 1 0 6496 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_108
timestamp 1698175906
transform 1 0 6720 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_110
timestamp 1698175906
transform 1 0 6832 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_127
timestamp 1698175906
transform 1 0 7784 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_131
timestamp 1698175906
transform 1 0 8008 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_194
timestamp 1698175906
transform 1 0 11536 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_205
timestamp 1698175906
transform 1 0 12152 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_209
timestamp 1698175906
transform 1 0 12376 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_212
timestamp 1698175906
transform 1 0 12544 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_220
timestamp 1698175906
transform 1 0 12992 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_255
timestamp 1698175906
transform 1 0 14952 0 -1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_271
timestamp 1698175906
transform 1 0 15848 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_279
timestamp 1698175906
transform 1 0 16296 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_282
timestamp 1698175906
transform 1 0 16464 0 -1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_314
timestamp 1698175906
transform 1 0 18256 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_322
timestamp 1698175906
transform 1 0 18704 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_2
timestamp 1698175906
transform 1 0 784 0 1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698175906
transform 1 0 2576 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_37
timestamp 1698175906
transform 1 0 2744 0 1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_101
timestamp 1698175906
transform 1 0 6328 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_107
timestamp 1698175906
transform 1 0 6664 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_111
timestamp 1698175906
transform 1 0 6888 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_115
timestamp 1698175906
transform 1 0 7112 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_124
timestamp 1698175906
transform 1 0 7616 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_140
timestamp 1698175906
transform 1 0 8512 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_142
timestamp 1698175906
transform 1 0 8624 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_177
timestamp 1698175906
transform 1 0 10584 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_181
timestamp 1698175906
transform 1 0 10808 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_188
timestamp 1698175906
transform 1 0 11200 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_227
timestamp 1698175906
transform 1 0 13384 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_231
timestamp 1698175906
transform 1 0 13608 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_244
timestamp 1698175906
transform 1 0 14336 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_247
timestamp 1698175906
transform 1 0 14504 0 1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_311
timestamp 1698175906
transform 1 0 18088 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_317
timestamp 1698175906
transform 1 0 18424 0 1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_2
timestamp 1698175906
transform 1 0 784 0 -1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_66
timestamp 1698175906
transform 1 0 4368 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_72
timestamp 1698175906
transform 1 0 4704 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_111
timestamp 1698175906
transform 1 0 6888 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_142
timestamp 1698175906
transform 1 0 8624 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_144
timestamp 1698175906
transform 1 0 8736 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_205
timestamp 1698175906
transform 1 0 12152 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_209
timestamp 1698175906
transform 1 0 12376 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_221
timestamp 1698175906
transform 1 0 13048 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_225
timestamp 1698175906
transform 1 0 13272 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_227
timestamp 1698175906
transform 1 0 13384 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_259
timestamp 1698175906
transform 1 0 15176 0 -1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_275
timestamp 1698175906
transform 1 0 16072 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_279
timestamp 1698175906
transform 1 0 16296 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_282
timestamp 1698175906
transform 1 0 16464 0 -1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_346
timestamp 1698175906
transform 1 0 20048 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_348
timestamp 1698175906
transform 1 0 20160 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_2
timestamp 1698175906
transform 1 0 784 0 1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698175906
transform 1 0 2576 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_37
timestamp 1698175906
transform 1 0 2744 0 1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_69
timestamp 1698175906
transform 1 0 4536 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_73
timestamp 1698175906
transform 1 0 4760 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_75
timestamp 1698175906
transform 1 0 4872 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_107
timestamp 1698175906
transform 1 0 6664 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_114
timestamp 1698175906
transform 1 0 7056 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_116
timestamp 1698175906
transform 1 0 7168 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_173
timestamp 1698175906
transform 1 0 10360 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_177
timestamp 1698175906
transform 1 0 10584 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_185
timestamp 1698175906
transform 1 0 11032 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_187
timestamp 1698175906
transform 1 0 11144 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_238
timestamp 1698175906
transform 1 0 14000 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_242
timestamp 1698175906
transform 1 0 14224 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_244
timestamp 1698175906
transform 1 0 14336 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_260
timestamp 1698175906
transform 1 0 15232 0 1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_292
timestamp 1698175906
transform 1 0 17024 0 1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_308
timestamp 1698175906
transform 1 0 17920 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_312
timestamp 1698175906
transform 1 0 18144 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_314
timestamp 1698175906
transform 1 0 18256 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_317
timestamp 1698175906
transform 1 0 18424 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_321
timestamp 1698175906
transform 1 0 18648 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_2
timestamp 1698175906
transform 1 0 784 0 -1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_66
timestamp 1698175906
transform 1 0 4368 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_72
timestamp 1698175906
transform 1 0 4704 0 -1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_88
timestamp 1698175906
transform 1 0 5600 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_96
timestamp 1698175906
transform 1 0 6048 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_109
timestamp 1698175906
transform 1 0 6776 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_113
timestamp 1698175906
transform 1 0 7000 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_123
timestamp 1698175906
transform 1 0 7560 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_127
timestamp 1698175906
transform 1 0 7784 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_142
timestamp 1698175906
transform 1 0 8624 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_193
timestamp 1698175906
transform 1 0 11480 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_206
timestamp 1698175906
transform 1 0 12208 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_220
timestamp 1698175906
transform 1 0 12992 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_259
timestamp 1698175906
transform 1 0 15176 0 -1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_275
timestamp 1698175906
transform 1 0 16072 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_279
timestamp 1698175906
transform 1 0 16296 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_282
timestamp 1698175906
transform 1 0 16464 0 -1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_314
timestamp 1698175906
transform 1 0 18256 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_322
timestamp 1698175906
transform 1 0 18704 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_2
timestamp 1698175906
transform 1 0 784 0 1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698175906
transform 1 0 2576 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_37
timestamp 1698175906
transform 1 0 2744 0 1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_101
timestamp 1698175906
transform 1 0 6328 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_107
timestamp 1698175906
transform 1 0 6664 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_115
timestamp 1698175906
transform 1 0 7112 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_119
timestamp 1698175906
transform 1 0 7336 0 1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_135
timestamp 1698175906
transform 1 0 8232 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_143
timestamp 1698175906
transform 1 0 8680 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_147
timestamp 1698175906
transform 1 0 8904 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_183
timestamp 1698175906
transform 1 0 10920 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_191
timestamp 1698175906
transform 1 0 11368 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_202
timestamp 1698175906
transform 1 0 11984 0 1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_224
timestamp 1698175906
transform 1 0 13216 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_232
timestamp 1698175906
transform 1 0 13664 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_242
timestamp 1698175906
transform 1 0 14224 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_244
timestamp 1698175906
transform 1 0 14336 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_252
timestamp 1698175906
transform 1 0 14784 0 1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_284
timestamp 1698175906
transform 1 0 16576 0 1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_300
timestamp 1698175906
transform 1 0 17472 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_308
timestamp 1698175906
transform 1 0 17920 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_312
timestamp 1698175906
transform 1 0 18144 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_314
timestamp 1698175906
transform 1 0 18256 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_317
timestamp 1698175906
transform 1 0 18424 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_321
timestamp 1698175906
transform 1 0 18648 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_2
timestamp 1698175906
transform 1 0 784 0 -1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_66
timestamp 1698175906
transform 1 0 4368 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_72
timestamp 1698175906
transform 1 0 4704 0 -1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_117
timestamp 1698175906
transform 1 0 7224 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_128
timestamp 1698175906
transform 1 0 7840 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_132
timestamp 1698175906
transform 1 0 8064 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_142
timestamp 1698175906
transform 1 0 8624 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_146
timestamp 1698175906
transform 1 0 8848 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_148
timestamp 1698175906
transform 1 0 8960 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_163
timestamp 1698175906
transform 1 0 9800 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_177
timestamp 1698175906
transform 1 0 10584 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_212
timestamp 1698175906
transform 1 0 12544 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_216
timestamp 1698175906
transform 1 0 12768 0 -1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_282
timestamp 1698175906
transform 1 0 16464 0 -1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_314
timestamp 1698175906
transform 1 0 18256 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_322
timestamp 1698175906
transform 1 0 18704 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_28
timestamp 1698175906
transform 1 0 2240 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_32
timestamp 1698175906
transform 1 0 2464 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698175906
transform 1 0 2576 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_37
timestamp 1698175906
transform 1 0 2744 0 1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_101
timestamp 1698175906
transform 1 0 6328 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_111
timestamp 1698175906
transform 1 0 6888 0 1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_127
timestamp 1698175906
transform 1 0 7784 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_140
timestamp 1698175906
transform 1 0 8512 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_142
timestamp 1698175906
transform 1 0 8624 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_154
timestamp 1698175906
transform 1 0 9296 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_162
timestamp 1698175906
transform 1 0 9744 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_173
timestamp 1698175906
transform 1 0 10360 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_177
timestamp 1698175906
transform 1 0 10584 0 1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_193
timestamp 1698175906
transform 1 0 11480 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_207
timestamp 1698175906
transform 1 0 12264 0 1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_223
timestamp 1698175906
transform 1 0 13160 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_238
timestamp 1698175906
transform 1 0 14000 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_242
timestamp 1698175906
transform 1 0 14224 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_244
timestamp 1698175906
transform 1 0 14336 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_247
timestamp 1698175906
transform 1 0 14504 0 1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_311
timestamp 1698175906
transform 1 0 18088 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_317
timestamp 1698175906
transform 1 0 18424 0 1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_28
timestamp 1698175906
transform 1 0 2240 0 -1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_60
timestamp 1698175906
transform 1 0 4032 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_68
timestamp 1698175906
transform 1 0 4480 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_72
timestamp 1698175906
transform 1 0 4704 0 -1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_104
timestamp 1698175906
transform 1 0 6496 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_108
timestamp 1698175906
transform 1 0 6720 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_139
timestamp 1698175906
transform 1 0 8456 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_142
timestamp 1698175906
transform 1 0 8624 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_146
timestamp 1698175906
transform 1 0 8848 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_158
timestamp 1698175906
transform 1 0 9520 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_166
timestamp 1698175906
transform 1 0 9968 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_170
timestamp 1698175906
transform 1 0 10192 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_184
timestamp 1698175906
transform 1 0 10976 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_194
timestamp 1698175906
transform 1 0 11536 0 -1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_212
timestamp 1698175906
transform 1 0 12544 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_220
timestamp 1698175906
transform 1 0 12992 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_224
timestamp 1698175906
transform 1 0 13216 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_262
timestamp 1698175906
transform 1 0 15344 0 -1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_278
timestamp 1698175906
transform 1 0 16240 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_282
timestamp 1698175906
transform 1 0 16464 0 -1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_314
timestamp 1698175906
transform 1 0 18256 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_322
timestamp 1698175906
transform 1 0 18704 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_2
timestamp 1698175906
transform 1 0 784 0 1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698175906
transform 1 0 2576 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_37
timestamp 1698175906
transform 1 0 2744 0 1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_101
timestamp 1698175906
transform 1 0 6328 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_107
timestamp 1698175906
transform 1 0 6664 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_144
timestamp 1698175906
transform 1 0 8736 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_148
timestamp 1698175906
transform 1 0 8960 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_150
timestamp 1698175906
transform 1 0 9072 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_157
timestamp 1698175906
transform 1 0 9464 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_166
timestamp 1698175906
transform 1 0 9968 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_174
timestamp 1698175906
transform 1 0 10416 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_182
timestamp 1698175906
transform 1 0 10864 0 1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_214
timestamp 1698175906
transform 1 0 12656 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_234
timestamp 1698175906
transform 1 0 13776 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_241
timestamp 1698175906
transform 1 0 14168 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_252
timestamp 1698175906
transform 1 0 14784 0 1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_284
timestamp 1698175906
transform 1 0 16576 0 1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_300
timestamp 1698175906
transform 1 0 17472 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_308
timestamp 1698175906
transform 1 0 17920 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_312
timestamp 1698175906
transform 1 0 18144 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_314
timestamp 1698175906
transform 1 0 18256 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_317
timestamp 1698175906
transform 1 0 18424 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_321
timestamp 1698175906
transform 1 0 18648 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_2
timestamp 1698175906
transform 1 0 784 0 -1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_66
timestamp 1698175906
transform 1 0 4368 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_72
timestamp 1698175906
transform 1 0 4704 0 -1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_136
timestamp 1698175906
transform 1 0 8288 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_142
timestamp 1698175906
transform 1 0 8624 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_150
timestamp 1698175906
transform 1 0 9072 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_152
timestamp 1698175906
transform 1 0 9184 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_166
timestamp 1698175906
transform 1 0 9968 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_174
timestamp 1698175906
transform 1 0 10416 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_192
timestamp 1698175906
transform 1 0 11424 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_196
timestamp 1698175906
transform 1 0 11648 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_203
timestamp 1698175906
transform 1 0 12040 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_207
timestamp 1698175906
transform 1 0 12264 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_209
timestamp 1698175906
transform 1 0 12376 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_212
timestamp 1698175906
transform 1 0 12544 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_216
timestamp 1698175906
transform 1 0 12768 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_251
timestamp 1698175906
transform 1 0 14728 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_255
timestamp 1698175906
transform 1 0 14952 0 -1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_271
timestamp 1698175906
transform 1 0 15848 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_279
timestamp 1698175906
transform 1 0 16296 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_282
timestamp 1698175906
transform 1 0 16464 0 -1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_314
timestamp 1698175906
transform 1 0 18256 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_322
timestamp 1698175906
transform 1 0 18704 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_2
timestamp 1698175906
transform 1 0 784 0 1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698175906
transform 1 0 2576 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_37
timestamp 1698175906
transform 1 0 2744 0 1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_101
timestamp 1698175906
transform 1 0 6328 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_107
timestamp 1698175906
transform 1 0 6664 0 1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_123
timestamp 1698175906
transform 1 0 7560 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_127
timestamp 1698175906
transform 1 0 7784 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_129
timestamp 1698175906
transform 1 0 7896 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_159
timestamp 1698175906
transform 1 0 9576 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_171
timestamp 1698175906
transform 1 0 10248 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_177
timestamp 1698175906
transform 1 0 10584 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_210
timestamp 1698175906
transform 1 0 12432 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_214
timestamp 1698175906
transform 1 0 12656 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_247
timestamp 1698175906
transform 1 0 14504 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_251
timestamp 1698175906
transform 1 0 14728 0 1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_317
timestamp 1698175906
transform 1 0 18424 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_321
timestamp 1698175906
transform 1 0 18648 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_2
timestamp 1698175906
transform 1 0 784 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_66
timestamp 1698175906
transform 1 0 4368 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_72
timestamp 1698175906
transform 1 0 4704 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_136
timestamp 1698175906
transform 1 0 8288 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_142
timestamp 1698175906
transform 1 0 8624 0 -1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_201
timestamp 1698175906
transform 1 0 11928 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_205
timestamp 1698175906
transform 1 0 12152 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_209
timestamp 1698175906
transform 1 0 12376 0 -1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_212
timestamp 1698175906
transform 1 0 12544 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_276
timestamp 1698175906
transform 1 0 16128 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_282
timestamp 1698175906
transform 1 0 16464 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_346
timestamp 1698175906
transform 1 0 20048 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_348
timestamp 1698175906
transform 1 0 20160 0 -1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_2
timestamp 1698175906
transform 1 0 784 0 1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698175906
transform 1 0 2576 0 1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_37
timestamp 1698175906
transform 1 0 2744 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_101
timestamp 1698175906
transform 1 0 6328 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_107
timestamp 1698175906
transform 1 0 6664 0 1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_139
timestamp 1698175906
transform 1 0 8456 0 1 14112
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_155
timestamp 1698175906
transform 1 0 9352 0 1 14112
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_163
timestamp 1698175906
transform 1 0 9800 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_172
timestamp 1698175906
transform 1 0 10304 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_174
timestamp 1698175906
transform 1 0 10416 0 1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_177
timestamp 1698175906
transform 1 0 10584 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_186
timestamp 1698175906
transform 1 0 11088 0 1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_218
timestamp 1698175906
transform 1 0 12880 0 1 14112
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_234
timestamp 1698175906
transform 1 0 13776 0 1 14112
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_242
timestamp 1698175906
transform 1 0 14224 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_244
timestamp 1698175906
transform 1 0 14336 0 1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_247
timestamp 1698175906
transform 1 0 14504 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_311
timestamp 1698175906
transform 1 0 18088 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_317
timestamp 1698175906
transform 1 0 18424 0 1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_2
timestamp 1698175906
transform 1 0 784 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_66
timestamp 1698175906
transform 1 0 4368 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_72
timestamp 1698175906
transform 1 0 4704 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_136
timestamp 1698175906
transform 1 0 8288 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_142
timestamp 1698175906
transform 1 0 8624 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_206
timestamp 1698175906
transform 1 0 12208 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_212
timestamp 1698175906
transform 1 0 12544 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_276
timestamp 1698175906
transform 1 0 16128 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_282
timestamp 1698175906
transform 1 0 16464 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_346
timestamp 1698175906
transform 1 0 20048 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_348
timestamp 1698175906
transform 1 0 20160 0 -1 14896
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698175906
transform 1 0 784 0 1 14896
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698175906
transform 1 0 2576 0 1 14896
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_37
timestamp 1698175906
transform 1 0 2744 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_101
timestamp 1698175906
transform 1 0 6328 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_107
timestamp 1698175906
transform 1 0 6664 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_171
timestamp 1698175906
transform 1 0 10248 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_177
timestamp 1698175906
transform 1 0 10584 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_241
timestamp 1698175906
transform 1 0 14168 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_247
timestamp 1698175906
transform 1 0 14504 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_311
timestamp 1698175906
transform 1 0 18088 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_317
timestamp 1698175906
transform 1 0 18424 0 1 14896
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2
timestamp 1698175906
transform 1 0 784 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_66
timestamp 1698175906
transform 1 0 4368 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_72
timestamp 1698175906
transform 1 0 4704 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_136
timestamp 1698175906
transform 1 0 8288 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_142
timestamp 1698175906
transform 1 0 8624 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_206
timestamp 1698175906
transform 1 0 12208 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_212
timestamp 1698175906
transform 1 0 12544 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_276
timestamp 1698175906
transform 1 0 16128 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_282
timestamp 1698175906
transform 1 0 16464 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_346
timestamp 1698175906
transform 1 0 20048 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_348
timestamp 1698175906
transform 1 0 20160 0 -1 15680
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_2
timestamp 1698175906
transform 1 0 784 0 1 15680
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698175906
transform 1 0 2576 0 1 15680
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_37
timestamp 1698175906
transform 1 0 2744 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_101
timestamp 1698175906
transform 1 0 6328 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_107
timestamp 1698175906
transform 1 0 6664 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_171
timestamp 1698175906
transform 1 0 10248 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_177
timestamp 1698175906
transform 1 0 10584 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_241
timestamp 1698175906
transform 1 0 14168 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_247
timestamp 1698175906
transform 1 0 14504 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_311
timestamp 1698175906
transform 1 0 18088 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_317
timestamp 1698175906
transform 1 0 18424 0 1 15680
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2
timestamp 1698175906
transform 1 0 784 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_66
timestamp 1698175906
transform 1 0 4368 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_72
timestamp 1698175906
transform 1 0 4704 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_136
timestamp 1698175906
transform 1 0 8288 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_142
timestamp 1698175906
transform 1 0 8624 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_206
timestamp 1698175906
transform 1 0 12208 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_212
timestamp 1698175906
transform 1 0 12544 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_276
timestamp 1698175906
transform 1 0 16128 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_282
timestamp 1698175906
transform 1 0 16464 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_346
timestamp 1698175906
transform 1 0 20048 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_348
timestamp 1698175906
transform 1 0 20160 0 -1 16464
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698175906
transform 1 0 784 0 1 16464
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698175906
transform 1 0 2576 0 1 16464
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_37
timestamp 1698175906
transform 1 0 2744 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_101
timestamp 1698175906
transform 1 0 6328 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_107
timestamp 1698175906
transform 1 0 6664 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_171
timestamp 1698175906
transform 1 0 10248 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_177
timestamp 1698175906
transform 1 0 10584 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_241
timestamp 1698175906
transform 1 0 14168 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_247
timestamp 1698175906
transform 1 0 14504 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_311
timestamp 1698175906
transform 1 0 18088 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_317
timestamp 1698175906
transform 1 0 18424 0 1 16464
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_2
timestamp 1698175906
transform 1 0 784 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_66
timestamp 1698175906
transform 1 0 4368 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_72
timestamp 1698175906
transform 1 0 4704 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_136
timestamp 1698175906
transform 1 0 8288 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_142
timestamp 1698175906
transform 1 0 8624 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_206
timestamp 1698175906
transform 1 0 12208 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_212
timestamp 1698175906
transform 1 0 12544 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_276
timestamp 1698175906
transform 1 0 16128 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_282
timestamp 1698175906
transform 1 0 16464 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_346
timestamp 1698175906
transform 1 0 20048 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_348
timestamp 1698175906
transform 1 0 20160 0 -1 17248
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698175906
transform 1 0 784 0 1 17248
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698175906
transform 1 0 2576 0 1 17248
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_37
timestamp 1698175906
transform 1 0 2744 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_101
timestamp 1698175906
transform 1 0 6328 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_107
timestamp 1698175906
transform 1 0 6664 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_171
timestamp 1698175906
transform 1 0 10248 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_177
timestamp 1698175906
transform 1 0 10584 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_241
timestamp 1698175906
transform 1 0 14168 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_247
timestamp 1698175906
transform 1 0 14504 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_311
timestamp 1698175906
transform 1 0 18088 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_317
timestamp 1698175906
transform 1 0 18424 0 1 17248
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2
timestamp 1698175906
transform 1 0 784 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1698175906
transform 1 0 4368 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_72
timestamp 1698175906
transform 1 0 4704 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_136
timestamp 1698175906
transform 1 0 8288 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_142
timestamp 1698175906
transform 1 0 8624 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_206
timestamp 1698175906
transform 1 0 12208 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_212
timestamp 1698175906
transform 1 0 12544 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_276
timestamp 1698175906
transform 1 0 16128 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_282
timestamp 1698175906
transform 1 0 16464 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_346
timestamp 1698175906
transform 1 0 20048 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_348
timestamp 1698175906
transform 1 0 20160 0 -1 18032
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_2
timestamp 1698175906
transform 1 0 784 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698175906
transform 1 0 2576 0 1 18032
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_37
timestamp 1698175906
transform 1 0 2744 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_101
timestamp 1698175906
transform 1 0 6328 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_107
timestamp 1698175906
transform 1 0 6664 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_171
timestamp 1698175906
transform 1 0 10248 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_177
timestamp 1698175906
transform 1 0 10584 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_241
timestamp 1698175906
transform 1 0 14168 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_247
timestamp 1698175906
transform 1 0 14504 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_311
timestamp 1698175906
transform 1 0 18088 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_317
timestamp 1698175906
transform 1 0 18424 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_2
timestamp 1698175906
transform 1 0 784 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_66
timestamp 1698175906
transform 1 0 4368 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_72
timestamp 1698175906
transform 1 0 4704 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_136
timestamp 1698175906
transform 1 0 8288 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_142
timestamp 1698175906
transform 1 0 8624 0 -1 18816
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_150
timestamp 1698175906
transform 1 0 9072 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_154
timestamp 1698175906
transform 1 0 9296 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_156
timestamp 1698175906
transform 1 0 9408 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_183
timestamp 1698175906
transform 1 0 10920 0 -1 18816
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_199
timestamp 1698175906
transform 1 0 11816 0 -1 18816
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_207
timestamp 1698175906
transform 1 0 12264 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_209
timestamp 1698175906
transform 1 0 12376 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_238
timestamp 1698175906
transform 1 0 14000 0 -1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_270
timestamp 1698175906
transform 1 0 15792 0 -1 18816
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_278
timestamp 1698175906
transform 1 0 16240 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_282
timestamp 1698175906
transform 1 0 16464 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_346
timestamp 1698175906
transform 1 0 20048 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_348
timestamp 1698175906
transform 1 0 20160 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_2
timestamp 1698175906
transform 1 0 784 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_36
timestamp 1698175906
transform 1 0 2688 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_70
timestamp 1698175906
transform 1 0 4592 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_104
timestamp 1698175906
transform 1 0 6496 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_138
timestamp 1698175906
transform 1 0 8400 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_142
timestamp 1698175906
transform 1 0 8624 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_198
timestamp 1698175906
transform 1 0 11760 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_202
timestamp 1698175906
transform 1 0 11984 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_232
timestamp 1698175906
transform 1 0 13664 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_236
timestamp 1698175906
transform 1 0 13888 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_240
timestamp 1698175906
transform 1 0 14112 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_274
timestamp 1698175906
transform 1 0 16016 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_308
timestamp 1698175906
transform 1 0 17920 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_342
timestamp 1698175906
transform 1 0 19824 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_346
timestamp 1698175906
transform 1 0 20048 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_348
timestamp 1698175906
transform 1 0 20160 0 1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18760 0 1 13328
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output2
timestamp 1698175906
transform 1 0 9464 0 -1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output3
timestamp 1698175906
transform 1 0 10304 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output4
timestamp 1698175906
transform -1 0 2240 0 -1 12544
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output5
timestamp 1698175906
transform 1 0 12544 0 -1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output6
timestamp 1698175906
transform 1 0 18760 0 -1 9408
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output7
timestamp 1698175906
transform 1 0 18760 0 -1 13328
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output8
timestamp 1698175906
transform 1 0 18760 0 1 12544
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output9
timestamp 1698175906
transform 1 0 12488 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output10
timestamp 1698175906
transform 1 0 18760 0 -1 12544
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output11
timestamp 1698175906
transform 1 0 12824 0 -1 2352
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output12
timestamp 1698175906
transform 1 0 10640 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output13
timestamp 1698175906
transform 1 0 12208 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output14
timestamp 1698175906
transform 1 0 8736 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output15
timestamp 1698175906
transform -1 0 2240 0 1 8624
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output16
timestamp 1698175906
transform 1 0 18760 0 1 10976
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output17
timestamp 1698175906
transform -1 0 2240 0 1 11760
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output18
timestamp 1698175906
transform 1 0 18760 0 1 10192
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output19
timestamp 1698175906
transform 1 0 18760 0 -1 8624
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output20
timestamp 1698175906
transform -1 0 2240 0 -1 8624
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output21
timestamp 1698175906
transform 1 0 18760 0 -1 11760
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output22
timestamp 1698175906
transform 1 0 10808 0 -1 2352
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output23
timestamp 1698175906
transform 1 0 18760 0 1 8624
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output24
timestamp 1698175906
transform 1 0 8456 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output25
timestamp 1698175906
transform 1 0 14112 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output26
timestamp 1698175906
transform 1 0 18760 0 -1 10976
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_45 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 672 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698175906
transform -1 0 20328 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_46
timestamp 1698175906
transform 1 0 672 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698175906
transform -1 0 20328 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_47
timestamp 1698175906
transform 1 0 672 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698175906
transform -1 0 20328 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_48
timestamp 1698175906
transform 1 0 672 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698175906
transform -1 0 20328 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_49
timestamp 1698175906
transform 1 0 672 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698175906
transform -1 0 20328 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_50
timestamp 1698175906
transform 1 0 672 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698175906
transform -1 0 20328 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_51
timestamp 1698175906
transform 1 0 672 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698175906
transform -1 0 20328 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_52
timestamp 1698175906
transform 1 0 672 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698175906
transform -1 0 20328 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_53
timestamp 1698175906
transform 1 0 672 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698175906
transform -1 0 20328 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_54
timestamp 1698175906
transform 1 0 672 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698175906
transform -1 0 20328 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_55
timestamp 1698175906
transform 1 0 672 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698175906
transform -1 0 20328 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_56
timestamp 1698175906
transform 1 0 672 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698175906
transform -1 0 20328 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_57
timestamp 1698175906
transform 1 0 672 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698175906
transform -1 0 20328 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_58
timestamp 1698175906
transform 1 0 672 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698175906
transform -1 0 20328 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_59
timestamp 1698175906
transform 1 0 672 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698175906
transform -1 0 20328 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_60
timestamp 1698175906
transform 1 0 672 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698175906
transform -1 0 20328 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_61
timestamp 1698175906
transform 1 0 672 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698175906
transform -1 0 20328 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_62
timestamp 1698175906
transform 1 0 672 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698175906
transform -1 0 20328 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_63
timestamp 1698175906
transform 1 0 672 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698175906
transform -1 0 20328 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_64
timestamp 1698175906
transform 1 0 672 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698175906
transform -1 0 20328 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_65
timestamp 1698175906
transform 1 0 672 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698175906
transform -1 0 20328 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_66
timestamp 1698175906
transform 1 0 672 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698175906
transform -1 0 20328 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_67
timestamp 1698175906
transform 1 0 672 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698175906
transform -1 0 20328 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_68
timestamp 1698175906
transform 1 0 672 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698175906
transform -1 0 20328 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_69
timestamp 1698175906
transform 1 0 672 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698175906
transform -1 0 20328 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_70
timestamp 1698175906
transform 1 0 672 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698175906
transform -1 0 20328 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_71
timestamp 1698175906
transform 1 0 672 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698175906
transform -1 0 20328 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_72
timestamp 1698175906
transform 1 0 672 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698175906
transform -1 0 20328 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_73
timestamp 1698175906
transform 1 0 672 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698175906
transform -1 0 20328 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_74
timestamp 1698175906
transform 1 0 672 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698175906
transform -1 0 20328 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_75
timestamp 1698175906
transform 1 0 672 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698175906
transform -1 0 20328 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_76
timestamp 1698175906
transform 1 0 672 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698175906
transform -1 0 20328 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_77
timestamp 1698175906
transform 1 0 672 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698175906
transform -1 0 20328 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_78
timestamp 1698175906
transform 1 0 672 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698175906
transform -1 0 20328 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_79
timestamp 1698175906
transform 1 0 672 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698175906
transform -1 0 20328 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_80
timestamp 1698175906
transform 1 0 672 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698175906
transform -1 0 20328 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_81
timestamp 1698175906
transform 1 0 672 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698175906
transform -1 0 20328 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_82
timestamp 1698175906
transform 1 0 672 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698175906
transform -1 0 20328 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_83
timestamp 1698175906
transform 1 0 672 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698175906
transform -1 0 20328 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_84
timestamp 1698175906
transform 1 0 672 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698175906
transform -1 0 20328 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_85
timestamp 1698175906
transform 1 0 672 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698175906
transform -1 0 20328 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_86
timestamp 1698175906
transform 1 0 672 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698175906
transform -1 0 20328 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_87
timestamp 1698175906
transform 1 0 672 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698175906
transform -1 0 20328 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_88
timestamp 1698175906
transform 1 0 672 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698175906
transform -1 0 20328 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_89
timestamp 1698175906
transform 1 0 672 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698175906
transform -1 0 20328 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_90 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 2576 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_91
timestamp 1698175906
transform 1 0 4480 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_92
timestamp 1698175906
transform 1 0 6384 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_93
timestamp 1698175906
transform 1 0 8288 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_94
timestamp 1698175906
transform 1 0 10192 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_95
timestamp 1698175906
transform 1 0 12096 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_96
timestamp 1698175906
transform 1 0 14000 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_97
timestamp 1698175906
transform 1 0 15904 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_98
timestamp 1698175906
transform 1 0 17808 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_99
timestamp 1698175906
transform 1 0 19712 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_100
timestamp 1698175906
transform 1 0 4592 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_101
timestamp 1698175906
transform 1 0 8512 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_102
timestamp 1698175906
transform 1 0 12432 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_103
timestamp 1698175906
transform 1 0 16352 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_104
timestamp 1698175906
transform 1 0 2632 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_105
timestamp 1698175906
transform 1 0 6552 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_106
timestamp 1698175906
transform 1 0 10472 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_107
timestamp 1698175906
transform 1 0 14392 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_108
timestamp 1698175906
transform 1 0 18312 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_109
timestamp 1698175906
transform 1 0 4592 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_110
timestamp 1698175906
transform 1 0 8512 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_111
timestamp 1698175906
transform 1 0 12432 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_112
timestamp 1698175906
transform 1 0 16352 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_113
timestamp 1698175906
transform 1 0 2632 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_114
timestamp 1698175906
transform 1 0 6552 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_115
timestamp 1698175906
transform 1 0 10472 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_116
timestamp 1698175906
transform 1 0 14392 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_117
timestamp 1698175906
transform 1 0 18312 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_118
timestamp 1698175906
transform 1 0 4592 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_119
timestamp 1698175906
transform 1 0 8512 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_120
timestamp 1698175906
transform 1 0 12432 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_121
timestamp 1698175906
transform 1 0 16352 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_122
timestamp 1698175906
transform 1 0 2632 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_123
timestamp 1698175906
transform 1 0 6552 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_124
timestamp 1698175906
transform 1 0 10472 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_125
timestamp 1698175906
transform 1 0 14392 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_126
timestamp 1698175906
transform 1 0 18312 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_127
timestamp 1698175906
transform 1 0 4592 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_128
timestamp 1698175906
transform 1 0 8512 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_129
timestamp 1698175906
transform 1 0 12432 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_130
timestamp 1698175906
transform 1 0 16352 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_131
timestamp 1698175906
transform 1 0 2632 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_132
timestamp 1698175906
transform 1 0 6552 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_133
timestamp 1698175906
transform 1 0 10472 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_134
timestamp 1698175906
transform 1 0 14392 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_135
timestamp 1698175906
transform 1 0 18312 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_136
timestamp 1698175906
transform 1 0 4592 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_137
timestamp 1698175906
transform 1 0 8512 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_138
timestamp 1698175906
transform 1 0 12432 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_139
timestamp 1698175906
transform 1 0 16352 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_140
timestamp 1698175906
transform 1 0 2632 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_141
timestamp 1698175906
transform 1 0 6552 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_142
timestamp 1698175906
transform 1 0 10472 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_143
timestamp 1698175906
transform 1 0 14392 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_144
timestamp 1698175906
transform 1 0 18312 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_145
timestamp 1698175906
transform 1 0 4592 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_146
timestamp 1698175906
transform 1 0 8512 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_147
timestamp 1698175906
transform 1 0 12432 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_148
timestamp 1698175906
transform 1 0 16352 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_149
timestamp 1698175906
transform 1 0 2632 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_150
timestamp 1698175906
transform 1 0 6552 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_151
timestamp 1698175906
transform 1 0 10472 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_152
timestamp 1698175906
transform 1 0 14392 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_153
timestamp 1698175906
transform 1 0 18312 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_154
timestamp 1698175906
transform 1 0 4592 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_155
timestamp 1698175906
transform 1 0 8512 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_156
timestamp 1698175906
transform 1 0 12432 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_157
timestamp 1698175906
transform 1 0 16352 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_158
timestamp 1698175906
transform 1 0 2632 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_159
timestamp 1698175906
transform 1 0 6552 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_160
timestamp 1698175906
transform 1 0 10472 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_161
timestamp 1698175906
transform 1 0 14392 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_162
timestamp 1698175906
transform 1 0 18312 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_163
timestamp 1698175906
transform 1 0 4592 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_164
timestamp 1698175906
transform 1 0 8512 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_165
timestamp 1698175906
transform 1 0 12432 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_166
timestamp 1698175906
transform 1 0 16352 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_167
timestamp 1698175906
transform 1 0 2632 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_168
timestamp 1698175906
transform 1 0 6552 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_169
timestamp 1698175906
transform 1 0 10472 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_170
timestamp 1698175906
transform 1 0 14392 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_171
timestamp 1698175906
transform 1 0 18312 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_172
timestamp 1698175906
transform 1 0 4592 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_173
timestamp 1698175906
transform 1 0 8512 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_174
timestamp 1698175906
transform 1 0 12432 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_175
timestamp 1698175906
transform 1 0 16352 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_176
timestamp 1698175906
transform 1 0 2632 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_177
timestamp 1698175906
transform 1 0 6552 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_178
timestamp 1698175906
transform 1 0 10472 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_179
timestamp 1698175906
transform 1 0 14392 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_180
timestamp 1698175906
transform 1 0 18312 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_181
timestamp 1698175906
transform 1 0 4592 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_182
timestamp 1698175906
transform 1 0 8512 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_183
timestamp 1698175906
transform 1 0 12432 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_184
timestamp 1698175906
transform 1 0 16352 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_185
timestamp 1698175906
transform 1 0 2632 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_186
timestamp 1698175906
transform 1 0 6552 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_187
timestamp 1698175906
transform 1 0 10472 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_188
timestamp 1698175906
transform 1 0 14392 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_189
timestamp 1698175906
transform 1 0 18312 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_190
timestamp 1698175906
transform 1 0 4592 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_191
timestamp 1698175906
transform 1 0 8512 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_192
timestamp 1698175906
transform 1 0 12432 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_193
timestamp 1698175906
transform 1 0 16352 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_194
timestamp 1698175906
transform 1 0 2632 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_195
timestamp 1698175906
transform 1 0 6552 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_196
timestamp 1698175906
transform 1 0 10472 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_197
timestamp 1698175906
transform 1 0 14392 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_198
timestamp 1698175906
transform 1 0 18312 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_199
timestamp 1698175906
transform 1 0 4592 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_200
timestamp 1698175906
transform 1 0 8512 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_201
timestamp 1698175906
transform 1 0 12432 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_202
timestamp 1698175906
transform 1 0 16352 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_203
timestamp 1698175906
transform 1 0 2632 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_204
timestamp 1698175906
transform 1 0 6552 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_205
timestamp 1698175906
transform 1 0 10472 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_206
timestamp 1698175906
transform 1 0 14392 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_207
timestamp 1698175906
transform 1 0 18312 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_208
timestamp 1698175906
transform 1 0 4592 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_209
timestamp 1698175906
transform 1 0 8512 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_210
timestamp 1698175906
transform 1 0 12432 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_211
timestamp 1698175906
transform 1 0 16352 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_212
timestamp 1698175906
transform 1 0 2632 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_213
timestamp 1698175906
transform 1 0 6552 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_214
timestamp 1698175906
transform 1 0 10472 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_215
timestamp 1698175906
transform 1 0 14392 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_216
timestamp 1698175906
transform 1 0 18312 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_217
timestamp 1698175906
transform 1 0 4592 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_218
timestamp 1698175906
transform 1 0 8512 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_219
timestamp 1698175906
transform 1 0 12432 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_220
timestamp 1698175906
transform 1 0 16352 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_221
timestamp 1698175906
transform 1 0 2632 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_222
timestamp 1698175906
transform 1 0 6552 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_223
timestamp 1698175906
transform 1 0 10472 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_224
timestamp 1698175906
transform 1 0 14392 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_225
timestamp 1698175906
transform 1 0 18312 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_226
timestamp 1698175906
transform 1 0 4592 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_227
timestamp 1698175906
transform 1 0 8512 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_228
timestamp 1698175906
transform 1 0 12432 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_229
timestamp 1698175906
transform 1 0 16352 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_230
timestamp 1698175906
transform 1 0 2632 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_231
timestamp 1698175906
transform 1 0 6552 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_232
timestamp 1698175906
transform 1 0 10472 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_233
timestamp 1698175906
transform 1 0 14392 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_234
timestamp 1698175906
transform 1 0 18312 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_235
timestamp 1698175906
transform 1 0 4592 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_236
timestamp 1698175906
transform 1 0 8512 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_237
timestamp 1698175906
transform 1 0 12432 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_238
timestamp 1698175906
transform 1 0 16352 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_239
timestamp 1698175906
transform 1 0 2632 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_240
timestamp 1698175906
transform 1 0 6552 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_241
timestamp 1698175906
transform 1 0 10472 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_242
timestamp 1698175906
transform 1 0 14392 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_243
timestamp 1698175906
transform 1 0 18312 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_244
timestamp 1698175906
transform 1 0 4592 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_245
timestamp 1698175906
transform 1 0 8512 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_246
timestamp 1698175906
transform 1 0 12432 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_247
timestamp 1698175906
transform 1 0 16352 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_248
timestamp 1698175906
transform 1 0 2632 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_249
timestamp 1698175906
transform 1 0 6552 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_250
timestamp 1698175906
transform 1 0 10472 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_251
timestamp 1698175906
transform 1 0 14392 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_252
timestamp 1698175906
transform 1 0 18312 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_253
timestamp 1698175906
transform 1 0 4592 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_254
timestamp 1698175906
transform 1 0 8512 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_255
timestamp 1698175906
transform 1 0 12432 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_256
timestamp 1698175906
transform 1 0 16352 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_257
timestamp 1698175906
transform 1 0 2632 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_258
timestamp 1698175906
transform 1 0 6552 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_259
timestamp 1698175906
transform 1 0 10472 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_260
timestamp 1698175906
transform 1 0 14392 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_261
timestamp 1698175906
transform 1 0 18312 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_262
timestamp 1698175906
transform 1 0 4592 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_263
timestamp 1698175906
transform 1 0 8512 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_264
timestamp 1698175906
transform 1 0 12432 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_265
timestamp 1698175906
transform 1 0 16352 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_266
timestamp 1698175906
transform 1 0 2632 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_267
timestamp 1698175906
transform 1 0 6552 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_268
timestamp 1698175906
transform 1 0 10472 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_269
timestamp 1698175906
transform 1 0 14392 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_270
timestamp 1698175906
transform 1 0 18312 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_271
timestamp 1698175906
transform 1 0 4592 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_272
timestamp 1698175906
transform 1 0 8512 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_273
timestamp 1698175906
transform 1 0 12432 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_274
timestamp 1698175906
transform 1 0 16352 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_275
timestamp 1698175906
transform 1 0 2632 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_276
timestamp 1698175906
transform 1 0 6552 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_277
timestamp 1698175906
transform 1 0 10472 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_278
timestamp 1698175906
transform 1 0 14392 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_279
timestamp 1698175906
transform 1 0 18312 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_280
timestamp 1698175906
transform 1 0 4592 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_281
timestamp 1698175906
transform 1 0 8512 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_282
timestamp 1698175906
transform 1 0 12432 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_283
timestamp 1698175906
transform 1 0 16352 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_284
timestamp 1698175906
transform 1 0 2632 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_285
timestamp 1698175906
transform 1 0 6552 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_286
timestamp 1698175906
transform 1 0 10472 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_287
timestamp 1698175906
transform 1 0 14392 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_288
timestamp 1698175906
transform 1 0 18312 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_289
timestamp 1698175906
transform 1 0 4592 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_290
timestamp 1698175906
transform 1 0 8512 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_291
timestamp 1698175906
transform 1 0 12432 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_292
timestamp 1698175906
transform 1 0 16352 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_293
timestamp 1698175906
transform 1 0 2576 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_294
timestamp 1698175906
transform 1 0 4480 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_295
timestamp 1698175906
transform 1 0 6384 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_296
timestamp 1698175906
transform 1 0 8288 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_297
timestamp 1698175906
transform 1 0 10192 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_298
timestamp 1698175906
transform 1 0 12096 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_299
timestamp 1698175906
transform 1 0 14000 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_300
timestamp 1698175906
transform 1 0 15904 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_301
timestamp 1698175906
transform 1 0 17808 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_302
timestamp 1698175906
transform 1 0 19712 0 1 18816
box -43 -43 155 435
<< labels >>
flabel metal3 s 0 13776 400 13832 0 FreeSans 224 0 0 0 clk
port 0 nsew signal input
flabel metal3 s 20600 13104 21000 13160 0 FreeSans 224 0 0 0 segm[0]
port 1 nsew signal tristate
flabel metal2 s 9408 20600 9464 21000 0 FreeSans 224 90 0 0 segm[10]
port 2 nsew signal tristate
flabel metal2 s 10080 20600 10136 21000 0 FreeSans 224 90 0 0 segm[11]
port 3 nsew signal tristate
flabel metal3 s 0 12096 400 12152 0 FreeSans 224 0 0 0 segm[12]
port 4 nsew signal tristate
flabel metal2 s 12096 20600 12152 21000 0 FreeSans 224 90 0 0 segm[13]
port 5 nsew signal tristate
flabel metal3 s 20600 9072 21000 9128 0 FreeSans 224 0 0 0 segm[1]
port 6 nsew signal tristate
flabel metal3 s 20600 12768 21000 12824 0 FreeSans 224 0 0 0 segm[2]
port 7 nsew signal tristate
flabel metal3 s 20600 12432 21000 12488 0 FreeSans 224 0 0 0 segm[3]
port 8 nsew signal tristate
flabel metal2 s 12432 0 12488 400 0 FreeSans 224 90 0 0 segm[4]
port 9 nsew signal tristate
flabel metal3 s 20600 12096 21000 12152 0 FreeSans 224 0 0 0 segm[5]
port 10 nsew signal tristate
flabel metal2 s 12768 0 12824 400 0 FreeSans 224 90 0 0 segm[6]
port 11 nsew signal tristate
flabel metal2 s 11088 0 11144 400 0 FreeSans 224 90 0 0 segm[7]
port 12 nsew signal tristate
flabel metal2 s 11760 20600 11816 21000 0 FreeSans 224 90 0 0 segm[8]
port 13 nsew signal tristate
flabel metal2 s 8736 20600 8792 21000 0 FreeSans 224 90 0 0 segm[9]
port 14 nsew signal tristate
flabel metal3 s 0 8736 400 8792 0 FreeSans 224 0 0 0 sel[0]
port 15 nsew signal tristate
flabel metal3 s 20600 11088 21000 11144 0 FreeSans 224 0 0 0 sel[10]
port 16 nsew signal tristate
flabel metal3 s 0 11760 400 11816 0 FreeSans 224 0 0 0 sel[11]
port 17 nsew signal tristate
flabel metal3 s 20600 10080 21000 10136 0 FreeSans 224 0 0 0 sel[1]
port 18 nsew signal tristate
flabel metal3 s 20600 8400 21000 8456 0 FreeSans 224 0 0 0 sel[2]
port 19 nsew signal tristate
flabel metal3 s 0 8064 400 8120 0 FreeSans 224 0 0 0 sel[3]
port 20 nsew signal tristate
flabel metal3 s 20600 11424 21000 11480 0 FreeSans 224 0 0 0 sel[4]
port 21 nsew signal tristate
flabel metal2 s 10752 0 10808 400 0 FreeSans 224 90 0 0 sel[5]
port 22 nsew signal tristate
flabel metal3 s 20600 8736 21000 8792 0 FreeSans 224 0 0 0 sel[6]
port 23 nsew signal tristate
flabel metal2 s 8400 0 8456 400 0 FreeSans 224 90 0 0 sel[7]
port 24 nsew signal tristate
flabel metal2 s 13104 0 13160 400 0 FreeSans 224 90 0 0 sel[8]
port 25 nsew signal tristate
flabel metal3 s 20600 10416 21000 10472 0 FreeSans 224 0 0 0 sel[9]
port 26 nsew signal tristate
flabel metal4 s 2224 1538 2384 19238 0 FreeSans 640 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 17584 1538 17744 19238 0 FreeSans 640 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 9904 1538 10064 19238 0 FreeSans 640 90 0 0 vss
port 28 nsew ground bidirectional
rlabel metal1 10500 19208 10500 19208 0 vdd
rlabel metal1 10500 18816 10500 18816 0 vss
rlabel metal2 6412 7812 6412 7812 0 _000_
rlabel metal2 13552 8876 13552 8876 0 _001_
rlabel metal3 14336 10276 14336 10276 0 _002_
rlabel metal2 5908 8652 5908 8652 0 _003_
rlabel metal2 11900 9016 11900 9016 0 _004_
rlabel metal2 12236 6636 12236 6636 0 _005_
rlabel metal2 12040 7644 12040 7644 0 _006_
rlabel metal2 13888 8484 13888 8484 0 _007_
rlabel metal2 13972 10836 13972 10836 0 _008_
rlabel metal2 6748 11732 6748 11732 0 _009_
rlabel metal2 13244 13160 13244 13160 0 _010_
rlabel metal2 13412 12964 13412 12964 0 _011_
rlabel metal2 13860 12180 13860 12180 0 _012_
rlabel metal2 10752 13860 10752 13860 0 _013_
rlabel metal2 8260 12376 8260 12376 0 _014_
rlabel metal3 8988 13076 8988 13076 0 _015_
rlabel metal2 9940 13720 9940 13720 0 _016_
rlabel metal2 7980 12152 7980 12152 0 _017_
rlabel metal2 11284 13356 11284 13356 0 _018_
rlabel metal2 12236 10192 12236 10192 0 _019_
rlabel metal2 7644 6692 7644 6692 0 _020_
rlabel metal2 10108 7028 10108 7028 0 _021_
rlabel metal2 8092 10164 8092 10164 0 _022_
rlabel metal2 7140 9296 7140 9296 0 _023_
rlabel metal2 7364 7812 7364 7812 0 _024_
rlabel metal2 8624 7308 8624 7308 0 _025_
rlabel metal2 10164 6636 10164 6636 0 _026_
rlabel metal2 11284 11284 11284 11284 0 _027_
rlabel metal2 7924 8820 7924 8820 0 _028_
rlabel metal2 7756 8232 7756 8232 0 _029_
rlabel metal2 14308 9044 14308 9044 0 _030_
rlabel metal2 8820 8008 8820 8008 0 _031_
rlabel metal2 10724 7364 10724 7364 0 _032_
rlabel metal2 10780 6888 10780 6888 0 _033_
rlabel metal2 10248 11172 10248 11172 0 _034_
rlabel metal2 11676 11564 11676 11564 0 _035_
rlabel metal2 6804 8120 6804 8120 0 _036_
rlabel metal2 7308 8848 7308 8848 0 _037_
rlabel metal2 13468 8792 13468 8792 0 _038_
rlabel metal2 13636 9268 13636 9268 0 _039_
rlabel metal2 13748 8876 13748 8876 0 _040_
rlabel metal2 14924 10444 14924 10444 0 _041_
rlabel metal2 7196 8960 7196 8960 0 _042_
rlabel metal2 6972 8736 6972 8736 0 _043_
rlabel metal2 7056 8540 7056 8540 0 _044_
rlabel metal2 5796 8568 5796 8568 0 _045_
rlabel metal2 11676 9268 11676 9268 0 _046_
rlabel metal3 12544 6860 12544 6860 0 _047_
rlabel metal2 12124 7812 12124 7812 0 _048_
rlabel metal2 11900 7784 11900 7784 0 _049_
rlabel metal2 13916 8904 13916 8904 0 _050_
rlabel metal2 14084 9156 14084 9156 0 _051_
rlabel metal2 13692 11480 13692 11480 0 _052_
rlabel metal3 14336 11172 14336 11172 0 _053_
rlabel metal2 8316 11564 8316 11564 0 _054_
rlabel metal2 6804 11788 6804 11788 0 _055_
rlabel metal3 11088 12348 11088 12348 0 _056_
rlabel metal2 14084 12796 14084 12796 0 _057_
rlabel metal2 14476 12936 14476 12936 0 _058_
rlabel metal2 14644 12824 14644 12824 0 _059_
rlabel metal2 13916 12292 13916 12292 0 _060_
rlabel metal2 10248 14252 10248 14252 0 _061_
rlabel metal2 10892 13692 10892 13692 0 _062_
rlabel via2 10052 12460 10052 12460 0 _063_
rlabel metal2 10164 11424 10164 11424 0 _064_
rlabel metal2 10612 12796 10612 12796 0 _065_
rlabel metal2 9380 12908 9380 12908 0 _066_
rlabel metal2 8428 12264 8428 12264 0 _067_
rlabel metal2 9632 13244 9632 13244 0 _068_
rlabel metal2 9604 12992 9604 12992 0 _069_
rlabel metal2 10108 14112 10108 14112 0 _070_
rlabel metal2 10276 11788 10276 11788 0 _071_
rlabel metal2 9800 13524 9800 13524 0 _072_
rlabel metal2 9548 11592 9548 11592 0 _073_
rlabel metal2 8092 11872 8092 11872 0 _074_
rlabel metal2 10836 12936 10836 12936 0 _075_
rlabel metal3 11592 13132 11592 13132 0 _076_
rlabel metal3 10304 10108 10304 10108 0 _077_
rlabel metal2 9828 11200 9828 11200 0 _078_
rlabel metal3 12264 11116 12264 11116 0 _079_
rlabel metal2 7448 10276 7448 10276 0 _080_
rlabel metal2 6972 10220 6972 10220 0 _081_
rlabel metal2 10388 9660 10388 9660 0 _082_
rlabel metal2 9548 9296 9548 9296 0 _083_
rlabel metal2 8484 10416 8484 10416 0 _084_
rlabel metal2 12628 10584 12628 10584 0 _085_
rlabel metal2 9940 8764 9940 8764 0 _086_
rlabel metal2 11452 9772 11452 9772 0 _087_
rlabel metal2 9324 11368 9324 11368 0 _088_
rlabel metal3 9576 9212 9576 9212 0 _089_
rlabel metal2 10388 8624 10388 8624 0 _090_
rlabel metal2 10892 10864 10892 10864 0 _091_
rlabel metal2 12124 6972 12124 6972 0 _092_
rlabel metal2 10332 10808 10332 10808 0 _093_
rlabel metal2 10920 8820 10920 8820 0 _094_
rlabel metal2 10948 10192 10948 10192 0 _095_
rlabel metal2 12684 10220 12684 10220 0 _096_
rlabel metal2 12964 10444 12964 10444 0 _097_
rlabel metal2 14700 10752 14700 10752 0 _098_
rlabel metal2 11984 6860 11984 6860 0 _099_
rlabel metal3 8652 6580 8652 6580 0 _100_
rlabel metal2 7476 9240 7476 9240 0 _101_
rlabel metal2 8708 8764 8708 8764 0 _102_
rlabel metal2 8820 11004 8820 11004 0 _103_
rlabel metal2 9828 7420 9828 7420 0 _104_
rlabel metal2 7420 8792 7420 8792 0 _105_
rlabel metal3 10052 7588 10052 7588 0 _106_
rlabel metal2 10248 10780 10248 10780 0 _107_
rlabel metal2 7504 8428 7504 8428 0 _108_
rlabel metal2 10892 7840 10892 7840 0 _109_
rlabel metal2 6692 10360 6692 10360 0 _110_
rlabel metal2 10780 8372 10780 8372 0 _111_
rlabel metal2 10332 7616 10332 7616 0 _112_
rlabel metal2 7140 8400 7140 8400 0 _113_
rlabel metal2 13972 11424 13972 11424 0 _114_
rlabel metal3 1239 13804 1239 13804 0 clk
rlabel metal2 11284 10220 11284 10220 0 clknet_0_clk
rlabel metal3 5992 10108 5992 10108 0 clknet_1_0__leaf_clk
rlabel metal2 13468 12320 13468 12320 0 clknet_1_1__leaf_clk
rlabel metal2 6468 10612 6468 10612 0 dut11.count\[0\]
rlabel metal3 6664 10388 6664 10388 0 dut11.count\[1\]
rlabel metal2 8428 8400 8428 8400 0 dut11.count\[2\]
rlabel metal2 9660 7434 9660 7434 0 dut11.count\[3\]
rlabel metal2 14308 13552 14308 13552 0 net1
rlabel metal2 14924 12348 14924 12348 0 net10
rlabel metal2 12908 3178 12908 3178 0 net11
rlabel metal3 10948 6804 10948 6804 0 net12
rlabel metal3 11396 14252 11396 14252 0 net13
rlabel metal2 8736 15960 8736 15960 0 net14
rlabel metal2 5012 8652 5012 8652 0 net15
rlabel metal2 15092 10892 15092 10892 0 net16
rlabel metal2 2156 11732 2156 11732 0 net17
rlabel metal2 15092 10192 15092 10192 0 net18
rlabel metal2 14252 8960 14252 8960 0 net19
rlabel metal2 9688 13636 9688 13636 0 net2
rlabel metal2 2156 8008 2156 8008 0 net20
rlabel metal3 15960 11508 15960 11508 0 net21
rlabel metal2 10948 3178 10948 3178 0 net22
rlabel metal2 14924 8932 14924 8932 0 net23
rlabel metal2 8540 2982 8540 2982 0 net24
rlabel metal3 13692 6916 13692 6916 0 net25
rlabel metal2 18956 10220 18956 10220 0 net26
rlabel metal2 10192 13860 10192 13860 0 net3
rlabel metal2 6916 12320 6916 12320 0 net4
rlabel metal2 12348 13916 12348 13916 0 net5
rlabel metal3 15960 8904 15960 8904 0 net6
rlabel metal2 14364 12852 14364 12852 0 net7
rlabel metal3 15610 12404 15610 12404 0 net8
rlabel metal2 12628 2982 12628 2982 0 net9
rlabel metal2 20020 13356 20020 13356 0 segm[0]
rlabel metal3 9744 18732 9744 18732 0 segm[10]
rlabel metal2 10108 19873 10108 19873 0 segm[11]
rlabel metal3 679 12124 679 12124 0 segm[12]
rlabel metal2 12124 19677 12124 19677 0 segm[13]
rlabel metal3 20321 9100 20321 9100 0 segm[1]
rlabel metal2 19964 12936 19964 12936 0 segm[2]
rlabel metal2 20020 12628 20020 12628 0 segm[3]
rlabel metal2 12460 1043 12460 1043 0 segm[4]
rlabel metal2 20020 12180 20020 12180 0 segm[5]
rlabel metal2 12796 1211 12796 1211 0 segm[6]
rlabel metal2 11116 1015 11116 1015 0 segm[7]
rlabel metal2 11788 19873 11788 19873 0 segm[8]
rlabel metal2 8764 19873 8764 19873 0 segm[9]
rlabel metal3 679 8764 679 8764 0 sel[0]
rlabel metal2 20020 11172 20020 11172 0 sel[10]
rlabel metal3 679 11788 679 11788 0 sel[11]
rlabel metal2 20020 10276 20020 10276 0 sel[1]
rlabel metal2 20020 8400 20020 8400 0 sel[2]
rlabel metal3 679 8092 679 8092 0 sel[3]
rlabel metal3 20321 11452 20321 11452 0 sel[4]
rlabel metal2 10780 1211 10780 1211 0 sel[5]
rlabel metal2 20020 8820 20020 8820 0 sel[6]
rlabel metal2 8428 1043 8428 1043 0 sel[7]
rlabel metal2 13132 1099 13132 1099 0 sel[8]
rlabel metal2 19964 10584 19964 10584 0 sel[9]
<< properties >>
string FIXED_BBOX 0 0 21000 21000
<< end >>
