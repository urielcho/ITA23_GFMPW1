magic
tech gf180mcuD
magscale 1 5
timestamp 1699641379
<< obsm1 >>
rect 672 1538 20328 19238
<< metal2 >>
rect 7392 20600 7448 21000
rect 7728 20600 7784 21000
rect 8064 20600 8120 21000
rect 9744 20600 9800 21000
rect 10080 20600 10136 21000
rect 11088 20600 11144 21000
rect 11424 20600 11480 21000
rect 9072 0 9128 400
rect 9408 0 9464 400
rect 10416 0 10472 400
rect 11424 0 11480 400
rect 12096 0 12152 400
<< obsm2 >>
rect 854 20570 7362 20600
rect 7478 20570 7698 20600
rect 7814 20570 8034 20600
rect 8150 20570 9714 20600
rect 9830 20570 10050 20600
rect 10166 20570 11058 20600
rect 11174 20570 11394 20600
rect 11510 20570 20034 20600
rect 854 430 20034 20570
rect 854 400 9042 430
rect 9158 400 9378 430
rect 9494 400 10386 430
rect 10502 400 11394 430
rect 11510 400 12066 430
rect 12182 400 20034 430
<< metal3 >>
rect 0 18480 400 18536
rect 0 14112 400 14168
rect 0 13440 400 13496
rect 20600 12768 21000 12824
rect 20600 12432 21000 12488
rect 20600 12096 21000 12152
rect 20600 11760 21000 11816
rect 20600 11088 21000 11144
rect 20600 10752 21000 10808
rect 0 10416 400 10472
rect 20600 10080 21000 10136
rect 20600 9072 21000 9128
rect 0 8400 400 8456
rect 0 8064 400 8120
rect 20600 8064 21000 8120
<< obsm3 >>
rect 400 18566 20600 19222
rect 430 18450 20600 18566
rect 400 14198 20600 18450
rect 430 14082 20600 14198
rect 400 13526 20600 14082
rect 430 13410 20600 13526
rect 400 12854 20600 13410
rect 400 12738 20570 12854
rect 400 12518 20600 12738
rect 400 12402 20570 12518
rect 400 12182 20600 12402
rect 400 12066 20570 12182
rect 400 11846 20600 12066
rect 400 11730 20570 11846
rect 400 11174 20600 11730
rect 400 11058 20570 11174
rect 400 10838 20600 11058
rect 400 10722 20570 10838
rect 400 10502 20600 10722
rect 430 10386 20600 10502
rect 400 10166 20600 10386
rect 400 10050 20570 10166
rect 400 9158 20600 10050
rect 400 9042 20570 9158
rect 400 8486 20600 9042
rect 430 8370 20600 8486
rect 400 8150 20600 8370
rect 430 8034 20570 8150
rect 400 1554 20600 8034
<< metal4 >>
rect 2224 1538 2384 19238
rect 9904 1538 10064 19238
rect 17584 1538 17744 19238
<< obsm4 >>
rect 9422 7569 9874 10127
rect 10094 7569 12810 10127
<< labels >>
rlabel metal3 s 0 14112 400 14168 6 clk
port 1 nsew signal input
rlabel metal3 s 0 18480 400 18536 6 segm[0]
port 2 nsew signal output
rlabel metal2 s 11424 0 11480 400 6 segm[10]
port 3 nsew signal output
rlabel metal3 s 0 13440 400 13496 6 segm[11]
port 4 nsew signal output
rlabel metal2 s 10416 0 10472 400 6 segm[12]
port 5 nsew signal output
rlabel metal3 s 0 8064 400 8120 6 segm[13]
port 6 nsew signal output
rlabel metal3 s 20600 11088 21000 11144 6 segm[1]
port 7 nsew signal output
rlabel metal3 s 20600 12768 21000 12824 6 segm[2]
port 8 nsew signal output
rlabel metal2 s 7392 20600 7448 21000 6 segm[3]
port 9 nsew signal output
rlabel metal3 s 20600 10752 21000 10808 6 segm[4]
port 10 nsew signal output
rlabel metal3 s 20600 11760 21000 11816 6 segm[5]
port 11 nsew signal output
rlabel metal2 s 9744 20600 9800 21000 6 segm[6]
port 12 nsew signal output
rlabel metal2 s 11088 20600 11144 21000 6 segm[7]
port 13 nsew signal output
rlabel metal3 s 0 8400 400 8456 6 segm[8]
port 14 nsew signal output
rlabel metal3 s 0 10416 400 10472 6 segm[9]
port 15 nsew signal output
rlabel metal3 s 20600 9072 21000 9128 6 sel[0]
port 16 nsew signal output
rlabel metal2 s 12096 0 12152 400 6 sel[10]
port 17 nsew signal output
rlabel metal2 s 9072 0 9128 400 6 sel[11]
port 18 nsew signal output
rlabel metal3 s 20600 12096 21000 12152 6 sel[1]
port 19 nsew signal output
rlabel metal3 s 20600 12432 21000 12488 6 sel[2]
port 20 nsew signal output
rlabel metal3 s 20600 8064 21000 8120 6 sel[3]
port 21 nsew signal output
rlabel metal2 s 9408 0 9464 400 6 sel[4]
port 22 nsew signal output
rlabel metal3 s 20600 10080 21000 10136 6 sel[5]
port 23 nsew signal output
rlabel metal2 s 10080 20600 10136 21000 6 sel[6]
port 24 nsew signal output
rlabel metal2 s 8064 20600 8120 21000 6 sel[7]
port 25 nsew signal output
rlabel metal2 s 7728 20600 7784 21000 6 sel[8]
port 26 nsew signal output
rlabel metal2 s 11424 20600 11480 21000 6 sel[9]
port 27 nsew signal output
rlabel metal4 s 2224 1538 2384 19238 6 vdd
port 28 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 19238 6 vdd
port 28 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 19238 6 vss
port 29 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 21000 21000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 482386
string GDS_FILE /home/urielcho/Proyectos_caravel/ITA23_GFMPW1b/openlane/ita19/runs/23_11_10_12_34/results/signoff/ita19.magic.gds
string GDS_START 162218
<< end >>

