// This is the unpowered netlist.
module ita17 (clk,
    segm,
    sel);
 input clk;
 output [13:0] segm;
 output [11:0] sel;

 wire net25;
 wire net26;
 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire \dut17.count[0] ;
 wire \dut17.count[1] ;
 wire \dut17.count[2] ;
 wire \dut17.count[3] ;
 wire net1;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;

 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__208__CLK (.I(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__209__CLK (.I(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__210__CLK (.I(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__211__CLK (.I(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__212__CLK (.I(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__213__CLK (.I(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__214__CLK (.I(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__215__CLK (.I(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__216__CLK (.I(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__217__CLK (.I(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__218__CLK (.I(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__219__CLK (.I(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__220__CLK (.I(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__221__CLK (.I(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__222__CLK (.I(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__223__CLK (.I(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__224__CLK (.I(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__225__CLK (.I(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__226__CLK (.I(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__227__CLK (.I(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__228__CLK (.I(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__229__CLK (.I(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__230__CLK (.I(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__231__CLK (.I(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__232__CLK (.I(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__233__CLK (.I(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_0_clk_I (.I(clk));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_14_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_14_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_15_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_16_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_19_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_20_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_23_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_23_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_25_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_25_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_27_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_28_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_29_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_29_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_30_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_30_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_31_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_32_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_43_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_43_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Left_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Left_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Left_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Left_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Left_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Left_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Left_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Left_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Left_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Left_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Left_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Left_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Left_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Left_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Left_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Left_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Left_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Left_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Left_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Right_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Left_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Right_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Left_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Right_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Left_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Right_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Left_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Left_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Right_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Left_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Right_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Left_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Right_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Left_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Right_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Left_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Right_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Left_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Right_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Left_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Right_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Left_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Right_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Left_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Right_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Left_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Right_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Left_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Left_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Right_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Left_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Right_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Left_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Right_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Left_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Right_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Left_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Right_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Left_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Left_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Left_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Left_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Left_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Left_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_90 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_91 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_92 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_93 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_94 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_95 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_96 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_97 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_98 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_99 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_139 ();
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _104_ (.I(\dut17.count[0] ),
    .Z(_064_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _105_ (.I(_064_),
    .Z(_065_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _106_ (.I(\dut17.count[1] ),
    .Z(_066_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _107_ (.I(_066_),
    .Z(_067_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _108_ (.I(\dut17.count[2] ),
    .ZN(_068_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _109_ (.I(_068_),
    .Z(_069_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _110_ (.I(\dut17.count[3] ),
    .Z(_070_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _111_ (.I(_070_),
    .Z(_071_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _112_ (.A1(_069_),
    .A2(_071_),
    .ZN(_072_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _113_ (.I(\dut17.count[2] ),
    .Z(_073_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _114_ (.A1(_073_),
    .A2(_070_),
    .Z(_074_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _115_ (.I(_074_),
    .Z(_075_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _116_ (.A1(net23),
    .A2(_075_),
    .ZN(_076_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _117_ (.A1(_065_),
    .A2(_067_),
    .A3(_072_),
    .B(_076_),
    .ZN(_000_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _118_ (.I(\dut17.count[0] ),
    .ZN(_077_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _119_ (.I(\dut17.count[1] ),
    .Z(_078_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _120_ (.I(_078_),
    .Z(_079_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _121_ (.A1(_077_),
    .A2(_079_),
    .ZN(_080_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _122_ (.I(\dut17.count[2] ),
    .Z(_081_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _123_ (.I(_070_),
    .ZN(_082_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _124_ (.A1(_081_),
    .A2(_082_),
    .ZN(_083_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _125_ (.I(_083_),
    .Z(_084_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _126_ (.I(_074_),
    .Z(_085_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _127_ (.A1(net21),
    .A2(_085_),
    .ZN(_086_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _128_ (.A1(_080_),
    .A2(_084_),
    .B(_086_),
    .ZN(_001_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _129_ (.I(\dut17.count[0] ),
    .Z(_087_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _130_ (.I(_066_),
    .ZN(_088_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _131_ (.A1(_087_),
    .A2(_088_),
    .ZN(_089_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _132_ (.A1(net20),
    .A2(_075_),
    .ZN(_090_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _133_ (.A1(_084_),
    .A2(_089_),
    .B(_090_),
    .ZN(_002_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _134_ (.I(_070_),
    .Z(_091_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _135_ (.I(_091_),
    .Z(_092_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _136_ (.A1(_073_),
    .A2(_064_),
    .A3(_078_),
    .Z(_093_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _137_ (.A1(_092_),
    .A2(_093_),
    .ZN(_094_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _138_ (.I(_082_),
    .Z(_095_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _139_ (.A1(_081_),
    .A2(_095_),
    .A3(_088_),
    .B(net24),
    .ZN(_096_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _140_ (.A1(_072_),
    .A2(_089_),
    .B1(_094_),
    .B2(_096_),
    .ZN(_003_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _141_ (.I(_077_),
    .Z(_004_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _142_ (.A1(_080_),
    .A2(_089_),
    .ZN(_005_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _143_ (.I(_068_),
    .Z(_097_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _144_ (.A1(\dut17.count[0] ),
    .A2(_078_),
    .Z(_098_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _145_ (.I(_098_),
    .Z(_099_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _146_ (.I(_078_),
    .Z(_100_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _147_ (.A1(\dut17.count[2] ),
    .A2(\dut17.count[3] ),
    .ZN(_101_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _148_ (.I(_101_),
    .Z(_102_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _149_ (.A1(_065_),
    .A2(_100_),
    .A3(_102_),
    .ZN(_103_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _150_ (.A1(_097_),
    .A2(_099_),
    .B(_103_),
    .ZN(_006_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _151_ (.I(_091_),
    .Z(_026_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _152_ (.A1(_026_),
    .A2(_099_),
    .ZN(_027_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _153_ (.A1(_084_),
    .A2(_099_),
    .B(_027_),
    .ZN(_007_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _154_ (.A1(net19),
    .A2(_074_),
    .ZN(_028_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _155_ (.A1(_065_),
    .A2(_067_),
    .A3(_083_),
    .B(_028_),
    .ZN(_008_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _156_ (.A1(net8),
    .A2(_085_),
    .ZN(_029_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _157_ (.A1(_103_),
    .A2(_029_),
    .ZN(_009_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _158_ (.A1(net17),
    .A2(_085_),
    .ZN(_030_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _159_ (.A1(_004_),
    .A2(_079_),
    .A3(_102_),
    .ZN(_031_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _160_ (.A1(_030_),
    .A2(_031_),
    .ZN(_010_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _161_ (.A1(_087_),
    .A2(_088_),
    .A3(_101_),
    .ZN(_032_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _162_ (.A1(net16),
    .A2(_085_),
    .ZN(_033_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _163_ (.A1(_032_),
    .A2(_033_),
    .ZN(_011_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _164_ (.A1(net13),
    .A2(_075_),
    .ZN(_034_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _165_ (.A1(_092_),
    .A2(_093_),
    .B(_034_),
    .ZN(_012_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _166_ (.A1(_087_),
    .A2(_066_),
    .A3(_101_),
    .Z(_035_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _167_ (.A1(_091_),
    .A2(_064_),
    .ZN(_036_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _168_ (.A1(_102_),
    .A2(_036_),
    .ZN(_037_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _169_ (.I(_073_),
    .Z(_038_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _170_ (.A1(_038_),
    .A2(_067_),
    .B(_026_),
    .C(net3),
    .ZN(_039_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _171_ (.A1(_069_),
    .A2(_071_),
    .A3(_079_),
    .ZN(_040_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _172_ (.A1(_035_),
    .A2(_037_),
    .B(_039_),
    .C(_040_),
    .ZN(_013_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _173_ (.A1(_081_),
    .A2(_100_),
    .B(_026_),
    .C(net4),
    .ZN(_041_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _174_ (.A1(_038_),
    .A2(_095_),
    .A3(_004_),
    .ZN(_042_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _175_ (.A1(_040_),
    .A2(_032_),
    .A3(_041_),
    .A4(_042_),
    .ZN(_014_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _176_ (.A1(_087_),
    .A2(_079_),
    .ZN(_043_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _177_ (.A1(_038_),
    .A2(_043_),
    .B(_026_),
    .ZN(_044_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _178_ (.I(_073_),
    .Z(_045_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _179_ (.A1(net10),
    .A2(_045_),
    .ZN(_046_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _180_ (.A1(_071_),
    .A2(_093_),
    .Z(_047_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _181_ (.A1(_031_),
    .A2(_044_),
    .B1(_046_),
    .B2(_047_),
    .ZN(_015_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _182_ (.A1(net11),
    .A2(_045_),
    .ZN(_048_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _183_ (.A1(_047_),
    .A2(_048_),
    .B(_035_),
    .ZN(_016_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _184_ (.A1(net12),
    .A2(_045_),
    .ZN(_049_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _185_ (.A1(_067_),
    .A2(_102_),
    .B1(_049_),
    .B2(_047_),
    .ZN(_017_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _186_ (.A1(net1),
    .A2(_075_),
    .ZN(_050_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _187_ (.A1(_004_),
    .A2(_084_),
    .B(_050_),
    .ZN(_018_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _188_ (.A1(net22),
    .A2(_095_),
    .B(_038_),
    .ZN(_051_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _189_ (.A1(_027_),
    .A2(_051_),
    .ZN(_019_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _190_ (.A1(net14),
    .A2(_045_),
    .A3(_092_),
    .ZN(_052_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _191_ (.A1(_065_),
    .A2(_040_),
    .B(_052_),
    .ZN(_020_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _192_ (.A1(_081_),
    .A2(_098_),
    .B(_091_),
    .ZN(_053_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _193_ (.A1(net15),
    .A2(_097_),
    .ZN(_054_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _194_ (.A1(_053_),
    .A2(_054_),
    .ZN(_021_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _195_ (.A1(_064_),
    .A2(_066_),
    .ZN(_055_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _196_ (.A1(_069_),
    .A2(_055_),
    .B(_095_),
    .C(net7),
    .ZN(_056_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _197_ (.A1(_097_),
    .A2(_080_),
    .B(_036_),
    .C(_056_),
    .ZN(_022_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _198_ (.I(_068_),
    .Z(_057_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _199_ (.A1(net9),
    .A2(_057_),
    .ZN(_058_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _200_ (.A1(_097_),
    .A2(_088_),
    .B(_036_),
    .ZN(_059_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _201_ (.A1(_053_),
    .A2(_058_),
    .B(_059_),
    .ZN(_023_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _202_ (.A1(_069_),
    .A2(_100_),
    .ZN(_060_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _203_ (.A1(net2),
    .A2(_057_),
    .ZN(_061_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _204_ (.A1(_092_),
    .A2(_099_),
    .A3(_060_),
    .B1(_061_),
    .B2(_053_),
    .ZN(_024_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _205_ (.A1(net5),
    .A2(_057_),
    .ZN(_062_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _206_ (.A1(_057_),
    .A2(_100_),
    .B(_077_),
    .C(_071_),
    .ZN(_063_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _207_ (.A1(_053_),
    .A2(_062_),
    .B1(_063_),
    .B2(_047_),
    .ZN(_025_));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _208_ (.D(_000_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net23));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _209_ (.D(_001_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net21));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _210_ (.D(_002_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net20));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _211_ (.D(_003_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net24));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _212_ (.D(_004_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(\dut17.count[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _213_ (.D(_005_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(\dut17.count[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _214_ (.D(_006_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(\dut17.count[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _215_ (.D(_007_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(\dut17.count[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _216_ (.D(_008_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net19));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _217_ (.D(_009_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net8));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _218_ (.D(_010_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net17));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _219_ (.D(_011_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net16));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _220_ (.D(_012_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net13));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _221_ (.D(_013_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net3));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _222_ (.D(_014_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net4));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _223_ (.D(_015_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net10));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _224_ (.D(_016_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net11));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _225_ (.D(_017_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net12));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _226_ (.D(_018_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _227_ (.D(_019_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net22));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _228_ (.D(_020_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net14));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _229_ (.D(_021_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net15));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _230_ (.D(_022_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net7));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _231_ (.D(_023_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net9));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _232_ (.D(_024_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net2));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _233_ (.D(_025_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net5));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _236_ (.I(net8),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _237_ (.I(net8),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_clk (.I(clk),
    .Z(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_1_0__f_clk (.I(clknet_0_clk),
    .Z(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_1_1__f_clk (.I(clknet_0_clk),
    .Z(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__tiel ita17_25 (.ZN(net25));
 gf180mcu_fd_sc_mcu7t5v0__tiel ita17_26 (.ZN(net26));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output1 (.I(net1),
    .Z(segm[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output10 (.I(net10),
    .Z(segm[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output11 (.I(net11),
    .Z(segm[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output12 (.I(net12),
    .Z(segm[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output13 (.I(net13),
    .Z(sel[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output14 (.I(net14),
    .Z(sel[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output15 (.I(net15),
    .Z(sel[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output16 (.I(net16),
    .Z(sel[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output17 (.I(net17),
    .Z(sel[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output18 (.I(net18),
    .Z(sel[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output19 (.I(net19),
    .Z(sel[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output2 (.I(net2),
    .Z(segm[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output20 (.I(net20),
    .Z(sel[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output21 (.I(net21),
    .Z(sel[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output22 (.I(net22),
    .Z(sel[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output23 (.I(net23),
    .Z(sel[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output24 (.I(net24),
    .Z(sel[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output3 (.I(net3),
    .Z(segm[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output4 (.I(net4),
    .Z(segm[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output5 (.I(net5),
    .Z(segm[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output6 (.I(net6),
    .Z(segm[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output7 (.I(net7),
    .Z(segm[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output8 (.I(net8),
    .Z(segm[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output9 (.I(net9),
    .Z(segm[6]));
 assign segm[2] = net25;
 assign segm[5] = net26;
endmodule

