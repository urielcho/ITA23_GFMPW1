magic
tech gf180mcuD
magscale 1 5
timestamp 1699642985
<< obsm1 >>
rect 672 1538 20328 19305
<< metal2 >>
rect 8064 20600 8120 21000
rect 8400 20600 8456 21000
rect 9408 20600 9464 21000
rect 10080 20600 10136 21000
rect 11088 20600 11144 21000
rect 12432 20600 12488 21000
rect 12768 20600 12824 21000
rect 13104 20600 13160 21000
rect 8064 0 8120 400
rect 9408 0 9464 400
rect 10080 0 10136 400
rect 11760 0 11816 400
rect 12096 0 12152 400
rect 12432 0 12488 400
rect 12768 0 12824 400
<< obsm2 >>
rect 854 20570 8034 20600
rect 8150 20570 8370 20600
rect 8486 20570 9378 20600
rect 9494 20570 10050 20600
rect 10166 20570 11058 20600
rect 11174 20570 12402 20600
rect 12518 20570 12738 20600
rect 12854 20570 13074 20600
rect 13190 20570 20034 20600
rect 854 430 20034 20570
rect 854 400 8034 430
rect 8150 400 9378 430
rect 9494 400 10050 430
rect 10166 400 11730 430
rect 11846 400 12066 430
rect 12182 400 12402 430
rect 12518 400 12738 430
rect 12854 400 20034 430
<< metal3 >>
rect 0 18144 400 18200
rect 0 14112 400 14168
rect 0 12096 400 12152
rect 0 11760 400 11816
rect 20600 11760 21000 11816
rect 20600 11088 21000 11144
rect 20600 10416 21000 10472
rect 20600 9072 21000 9128
rect 0 8736 400 8792
rect 20600 8736 21000 8792
rect 0 8400 400 8456
rect 0 7728 400 7784
<< obsm3 >>
rect 400 18230 20600 19306
rect 430 18114 20600 18230
rect 400 14198 20600 18114
rect 430 14082 20600 14198
rect 400 12182 20600 14082
rect 430 12066 20600 12182
rect 400 11846 20600 12066
rect 430 11730 20570 11846
rect 400 11174 20600 11730
rect 400 11058 20570 11174
rect 400 10502 20600 11058
rect 400 10386 20570 10502
rect 400 9158 20600 10386
rect 400 9042 20570 9158
rect 400 8822 20600 9042
rect 430 8706 20570 8822
rect 400 8486 20600 8706
rect 430 8370 20600 8486
rect 400 7814 20600 8370
rect 430 7698 20600 7814
rect 400 1554 20600 7698
<< metal4 >>
rect 2224 1538 2384 19238
rect 9904 1538 10064 19238
rect 17584 1538 17744 19238
<< obsm4 >>
rect 9758 8633 9786 12087
<< labels >>
rlabel metal3 s 0 14112 400 14168 6 clk
port 1 nsew signal input
rlabel metal3 s 0 18144 400 18200 6 segm[0]
port 2 nsew signal output
rlabel metal3 s 20600 10416 21000 10472 6 segm[10]
port 3 nsew signal output
rlabel metal3 s 20600 9072 21000 9128 6 segm[11]
port 4 nsew signal output
rlabel metal3 s 0 11760 400 11816 6 segm[12]
port 5 nsew signal output
rlabel metal2 s 9408 0 9464 400 6 segm[13]
port 6 nsew signal output
rlabel metal2 s 12432 0 12488 400 6 segm[1]
port 7 nsew signal output
rlabel metal2 s 12432 20600 12488 21000 6 segm[2]
port 8 nsew signal output
rlabel metal2 s 12768 20600 12824 21000 6 segm[3]
port 9 nsew signal output
rlabel metal2 s 12096 0 12152 400 6 segm[4]
port 10 nsew signal output
rlabel metal2 s 9408 20600 9464 21000 6 segm[5]
port 11 nsew signal output
rlabel metal3 s 0 12096 400 12152 6 segm[6]
port 12 nsew signal output
rlabel metal3 s 0 7728 400 7784 6 segm[7]
port 13 nsew signal output
rlabel metal3 s 0 8736 400 8792 6 segm[8]
port 14 nsew signal output
rlabel metal3 s 20600 8736 21000 8792 6 segm[9]
port 15 nsew signal output
rlabel metal3 s 20600 11088 21000 11144 6 sel[0]
port 16 nsew signal output
rlabel metal3 s 0 8400 400 8456 6 sel[10]
port 17 nsew signal output
rlabel metal2 s 8064 0 8120 400 6 sel[11]
port 18 nsew signal output
rlabel metal2 s 8400 20600 8456 21000 6 sel[1]
port 19 nsew signal output
rlabel metal2 s 8064 20600 8120 21000 6 sel[2]
port 20 nsew signal output
rlabel metal2 s 10080 20600 10136 21000 6 sel[3]
port 21 nsew signal output
rlabel metal2 s 13104 20600 13160 21000 6 sel[4]
port 22 nsew signal output
rlabel metal2 s 12768 0 12824 400 6 sel[5]
port 23 nsew signal output
rlabel metal3 s 20600 11760 21000 11816 6 sel[6]
port 24 nsew signal output
rlabel metal2 s 11088 20600 11144 21000 6 sel[7]
port 25 nsew signal output
rlabel metal2 s 10080 0 10136 400 6 sel[8]
port 26 nsew signal output
rlabel metal2 s 11760 0 11816 400 6 sel[9]
port 27 nsew signal output
rlabel metal4 s 2224 1538 2384 19238 6 vdd
port 28 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 19238 6 vdd
port 28 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 19238 6 vss
port 29 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 21000 21000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 507360
string GDS_FILE /home/urielcho/Proyectos_caravel/ITA23_GFMPW1b/openlane/ita59/runs/23_11_10_13_01/results/signoff/ita59.magic.gds
string GDS_START 168648
<< end >>

