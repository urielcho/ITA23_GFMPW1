magic
tech gf180mcuD
magscale 1 5
timestamp 1699641240
<< metal1 >>
rect 672 19221 20328 19238
rect 672 19195 2239 19221
rect 2265 19195 2291 19221
rect 2317 19195 2343 19221
rect 2369 19195 17599 19221
rect 17625 19195 17651 19221
rect 17677 19195 17703 19221
rect 17729 19195 20328 19221
rect 672 19178 20328 19195
rect 9311 19137 9337 19143
rect 9311 19105 9337 19111
rect 11215 19137 11241 19143
rect 11215 19105 11241 19111
rect 12783 19137 12809 19143
rect 12783 19105 12809 19111
rect 9025 18999 9031 19025
rect 9057 18999 9063 19025
rect 10705 18999 10711 19025
rect 10737 18999 10743 19025
rect 12273 18999 12279 19025
rect 12305 18999 12311 19025
rect 10375 18969 10401 18975
rect 10375 18937 10401 18943
rect 672 18829 20328 18846
rect 672 18803 9919 18829
rect 9945 18803 9971 18829
rect 9997 18803 10023 18829
rect 10049 18803 20328 18829
rect 672 18786 20328 18803
rect 9199 18745 9225 18751
rect 9199 18713 9225 18719
rect 11047 18745 11073 18751
rect 11047 18713 11073 18719
rect 13119 18745 13145 18751
rect 13119 18713 13145 18719
rect 20119 18689 20145 18695
rect 20119 18657 20145 18663
rect 8689 18607 8695 18633
rect 8721 18607 8727 18633
rect 10537 18607 10543 18633
rect 10569 18607 10575 18633
rect 12609 18607 12615 18633
rect 12641 18607 12647 18633
rect 672 18437 20328 18454
rect 672 18411 2239 18437
rect 2265 18411 2291 18437
rect 2317 18411 2343 18437
rect 2369 18411 17599 18437
rect 17625 18411 17651 18437
rect 17677 18411 17703 18437
rect 17729 18411 20328 18437
rect 672 18394 20328 18411
rect 672 18045 20328 18062
rect 672 18019 9919 18045
rect 9945 18019 9971 18045
rect 9997 18019 10023 18045
rect 10049 18019 20328 18045
rect 672 18002 20328 18019
rect 672 17653 20328 17670
rect 672 17627 2239 17653
rect 2265 17627 2291 17653
rect 2317 17627 2343 17653
rect 2369 17627 17599 17653
rect 17625 17627 17651 17653
rect 17677 17627 17703 17653
rect 17729 17627 20328 17653
rect 672 17610 20328 17627
rect 672 17261 20328 17278
rect 672 17235 9919 17261
rect 9945 17235 9971 17261
rect 9997 17235 10023 17261
rect 10049 17235 20328 17261
rect 672 17218 20328 17235
rect 672 16869 20328 16886
rect 672 16843 2239 16869
rect 2265 16843 2291 16869
rect 2317 16843 2343 16869
rect 2369 16843 17599 16869
rect 17625 16843 17651 16869
rect 17677 16843 17703 16869
rect 17729 16843 20328 16869
rect 672 16826 20328 16843
rect 672 16477 20328 16494
rect 672 16451 9919 16477
rect 9945 16451 9971 16477
rect 9997 16451 10023 16477
rect 10049 16451 20328 16477
rect 672 16434 20328 16451
rect 672 16085 20328 16102
rect 672 16059 2239 16085
rect 2265 16059 2291 16085
rect 2317 16059 2343 16085
rect 2369 16059 17599 16085
rect 17625 16059 17651 16085
rect 17677 16059 17703 16085
rect 17729 16059 20328 16085
rect 672 16042 20328 16059
rect 672 15693 20328 15710
rect 672 15667 9919 15693
rect 9945 15667 9971 15693
rect 9997 15667 10023 15693
rect 10049 15667 20328 15693
rect 672 15650 20328 15667
rect 672 15301 20328 15318
rect 672 15275 2239 15301
rect 2265 15275 2291 15301
rect 2317 15275 2343 15301
rect 2369 15275 17599 15301
rect 17625 15275 17651 15301
rect 17677 15275 17703 15301
rect 17729 15275 20328 15301
rect 672 15258 20328 15275
rect 672 14909 20328 14926
rect 672 14883 9919 14909
rect 9945 14883 9971 14909
rect 9997 14883 10023 14909
rect 10049 14883 20328 14909
rect 672 14866 20328 14883
rect 672 14517 20328 14534
rect 672 14491 2239 14517
rect 2265 14491 2291 14517
rect 2317 14491 2343 14517
rect 2369 14491 17599 14517
rect 17625 14491 17651 14517
rect 17677 14491 17703 14517
rect 17729 14491 20328 14517
rect 672 14474 20328 14491
rect 672 14125 20328 14142
rect 672 14099 9919 14125
rect 9945 14099 9971 14125
rect 9997 14099 10023 14125
rect 10049 14099 20328 14125
rect 672 14082 20328 14099
rect 8969 13903 8975 13929
rect 9001 13903 9007 13929
rect 10761 13903 10767 13929
rect 10793 13903 10799 13929
rect 18937 13903 18943 13929
rect 18969 13903 18975 13929
rect 8863 13873 8889 13879
rect 12727 13873 12753 13879
rect 9361 13847 9367 13873
rect 9393 13847 9399 13873
rect 10425 13847 10431 13873
rect 10457 13847 10463 13873
rect 11153 13847 11159 13873
rect 11185 13847 11191 13873
rect 12217 13847 12223 13873
rect 12249 13847 12255 13873
rect 19945 13847 19951 13873
rect 19977 13847 19983 13873
rect 8863 13841 8889 13847
rect 12727 13841 12753 13847
rect 672 13733 20328 13750
rect 672 13707 2239 13733
rect 2265 13707 2291 13733
rect 2317 13707 2343 13733
rect 2369 13707 17599 13733
rect 17625 13707 17651 13733
rect 17677 13707 17703 13733
rect 17729 13707 20328 13733
rect 672 13690 20328 13707
rect 20007 13593 20033 13599
rect 8521 13567 8527 13593
rect 8553 13567 8559 13593
rect 20007 13561 20033 13567
rect 8751 13537 8777 13543
rect 7065 13511 7071 13537
rect 7097 13511 7103 13537
rect 8751 13505 8777 13511
rect 9367 13537 9393 13543
rect 9367 13505 9393 13511
rect 10151 13537 10177 13543
rect 10151 13505 10177 13511
rect 11271 13537 11297 13543
rect 11271 13505 11297 13511
rect 11831 13537 11857 13543
rect 13785 13511 13791 13537
rect 13817 13511 13823 13537
rect 18825 13511 18831 13537
rect 18857 13511 18863 13537
rect 11831 13505 11857 13511
rect 8695 13481 8721 13487
rect 7457 13455 7463 13481
rect 7489 13455 7495 13481
rect 8695 13449 8721 13455
rect 9087 13481 9113 13487
rect 9087 13449 9113 13455
rect 9479 13481 9505 13487
rect 9479 13449 9505 13455
rect 9535 13481 9561 13487
rect 9535 13449 9561 13455
rect 9983 13481 10009 13487
rect 9983 13449 10009 13455
rect 10095 13481 10121 13487
rect 10095 13449 10121 13455
rect 11383 13481 11409 13487
rect 11383 13449 11409 13455
rect 11439 13481 11465 13487
rect 11439 13449 11465 13455
rect 11663 13481 11689 13487
rect 11663 13449 11689 13455
rect 11775 13481 11801 13487
rect 11775 13449 11801 13455
rect 13175 13481 13201 13487
rect 13175 13449 13201 13455
rect 13231 13481 13257 13487
rect 13897 13455 13903 13481
rect 13929 13455 13935 13481
rect 13231 13449 13257 13455
rect 8807 13425 8833 13431
rect 8807 13393 8833 13399
rect 13063 13425 13089 13431
rect 13063 13393 13089 13399
rect 672 13341 20328 13358
rect 672 13315 9919 13341
rect 9945 13315 9971 13341
rect 9997 13315 10023 13341
rect 10049 13315 20328 13341
rect 672 13298 20328 13315
rect 8191 13257 8217 13263
rect 8191 13225 8217 13231
rect 8303 13201 8329 13207
rect 14401 13175 14407 13201
rect 14433 13175 14439 13201
rect 8303 13169 8329 13175
rect 8135 13145 8161 13151
rect 8135 13113 8161 13119
rect 8415 13145 8441 13151
rect 8415 13113 8441 13119
rect 8695 13145 8721 13151
rect 8695 13113 8721 13119
rect 8807 13145 8833 13151
rect 8807 13113 8833 13119
rect 8919 13145 8945 13151
rect 8919 13113 8945 13119
rect 9031 13145 9057 13151
rect 12609 13119 12615 13145
rect 12641 13119 12647 13145
rect 14289 13119 14295 13145
rect 14321 13119 14327 13145
rect 18825 13119 18831 13145
rect 18857 13119 18863 13145
rect 9031 13113 9057 13119
rect 6567 13089 6593 13095
rect 14631 13089 14657 13095
rect 13001 13063 13007 13089
rect 13033 13063 13039 13089
rect 14065 13063 14071 13089
rect 14097 13063 14103 13089
rect 19945 13063 19951 13089
rect 19977 13063 19983 13089
rect 6567 13057 6593 13063
rect 14631 13057 14657 13063
rect 672 12949 20328 12966
rect 672 12923 2239 12949
rect 2265 12923 2291 12949
rect 2317 12923 2343 12949
rect 2369 12923 17599 12949
rect 17625 12923 17651 12949
rect 17677 12923 17703 12949
rect 17729 12923 20328 12949
rect 672 12906 20328 12923
rect 967 12809 993 12815
rect 9479 12809 9505 12815
rect 20007 12809 20033 12815
rect 4993 12783 4999 12809
rect 5025 12783 5031 12809
rect 8185 12783 8191 12809
rect 8217 12783 8223 12809
rect 9249 12783 9255 12809
rect 9281 12783 9287 12809
rect 12161 12783 12167 12809
rect 12193 12783 12199 12809
rect 14009 12783 14015 12809
rect 14041 12783 14047 12809
rect 967 12777 993 12783
rect 9479 12777 9505 12783
rect 20007 12777 20033 12783
rect 2137 12727 2143 12753
rect 2169 12727 2175 12753
rect 6449 12727 6455 12753
rect 6481 12727 6487 12753
rect 7849 12727 7855 12753
rect 7881 12727 7887 12753
rect 10761 12727 10767 12753
rect 10793 12727 10799 12753
rect 12553 12727 12559 12753
rect 12585 12727 12591 12753
rect 18825 12727 18831 12753
rect 18857 12727 18863 12753
rect 6959 12697 6985 12703
rect 6057 12671 6063 12697
rect 6089 12671 6095 12697
rect 9977 12671 9983 12697
rect 10009 12671 10015 12697
rect 11097 12671 11103 12697
rect 11129 12671 11135 12697
rect 12945 12671 12951 12697
rect 12977 12671 12983 12697
rect 6959 12665 6985 12671
rect 6791 12641 6817 12647
rect 6791 12609 6817 12615
rect 6903 12641 6929 12647
rect 6903 12609 6929 12615
rect 7015 12641 7041 12647
rect 7015 12609 7041 12615
rect 9815 12641 9841 12647
rect 9815 12609 9841 12615
rect 12391 12641 12417 12647
rect 12391 12609 12417 12615
rect 14239 12641 14265 12647
rect 14239 12609 14265 12615
rect 672 12557 20328 12574
rect 672 12531 9919 12557
rect 9945 12531 9971 12557
rect 9997 12531 10023 12557
rect 10049 12531 20328 12557
rect 672 12514 20328 12531
rect 8807 12473 8833 12479
rect 8807 12441 8833 12447
rect 8863 12473 8889 12479
rect 8863 12441 8889 12447
rect 8919 12473 8945 12479
rect 8919 12441 8945 12447
rect 11775 12473 11801 12479
rect 11775 12441 11801 12447
rect 12783 12473 12809 12479
rect 12783 12441 12809 12447
rect 13231 12473 13257 12479
rect 13231 12441 13257 12447
rect 13511 12473 13537 12479
rect 13511 12441 13537 12447
rect 13623 12473 13649 12479
rect 13623 12441 13649 12447
rect 7631 12417 7657 12423
rect 7631 12385 7657 12391
rect 7687 12417 7713 12423
rect 7687 12385 7713 12391
rect 12895 12417 12921 12423
rect 12895 12385 12921 12391
rect 12951 12417 12977 12423
rect 12951 12385 12977 12391
rect 13455 12417 13481 12423
rect 13455 12385 13481 12391
rect 8751 12361 8777 12367
rect 11887 12361 11913 12367
rect 6001 12335 6007 12361
rect 6033 12335 6039 12361
rect 9025 12335 9031 12361
rect 9057 12335 9063 12361
rect 11265 12335 11271 12361
rect 11297 12335 11303 12361
rect 11489 12335 11495 12361
rect 11521 12335 11527 12361
rect 11657 12335 11663 12361
rect 11689 12335 11695 12361
rect 8751 12329 8777 12335
rect 11887 12329 11913 12335
rect 13175 12361 13201 12367
rect 13175 12329 13201 12335
rect 7911 12305 7937 12311
rect 6337 12279 6343 12305
rect 6369 12279 6375 12305
rect 7401 12279 7407 12305
rect 7433 12279 7439 12305
rect 9865 12279 9871 12305
rect 9897 12279 9903 12305
rect 10929 12279 10935 12305
rect 10961 12279 10967 12305
rect 11713 12279 11719 12305
rect 11745 12279 11751 12305
rect 7911 12273 7937 12279
rect 7631 12249 7657 12255
rect 7631 12217 7657 12223
rect 13231 12249 13257 12255
rect 13231 12217 13257 12223
rect 672 12165 20328 12182
rect 672 12139 2239 12165
rect 2265 12139 2291 12165
rect 2317 12139 2343 12165
rect 2369 12139 17599 12165
rect 17625 12139 17651 12165
rect 17677 12139 17703 12165
rect 17729 12139 20328 12165
rect 672 12122 20328 12139
rect 6399 12081 6425 12087
rect 6399 12049 6425 12055
rect 10655 12081 10681 12087
rect 10655 12049 10681 12055
rect 6791 12025 6817 12031
rect 6791 11993 6817 11999
rect 11719 12025 11745 12031
rect 11719 11993 11745 11999
rect 6847 11969 6873 11975
rect 6847 11937 6873 11943
rect 7071 11969 7097 11975
rect 7071 11937 7097 11943
rect 10711 11969 10737 11975
rect 10985 11943 10991 11969
rect 11017 11943 11023 11969
rect 10711 11937 10737 11943
rect 6399 11913 6425 11919
rect 6399 11881 6425 11887
rect 6455 11913 6481 11919
rect 6455 11881 6481 11887
rect 8135 11913 8161 11919
rect 8135 11881 8161 11887
rect 10823 11913 10849 11919
rect 10823 11881 10849 11887
rect 11103 11913 11129 11919
rect 11103 11881 11129 11887
rect 11439 11913 11465 11919
rect 11439 11881 11465 11887
rect 11495 11913 11521 11919
rect 11495 11881 11521 11887
rect 6735 11857 6761 11863
rect 6735 11825 6761 11831
rect 8191 11857 8217 11863
rect 8191 11825 8217 11831
rect 11047 11857 11073 11863
rect 11047 11825 11073 11831
rect 11383 11857 11409 11863
rect 11383 11825 11409 11831
rect 672 11773 20328 11790
rect 672 11747 9919 11773
rect 9945 11747 9971 11773
rect 9997 11747 10023 11773
rect 10049 11747 20328 11773
rect 672 11730 20328 11747
rect 9535 11689 9561 11695
rect 9535 11657 9561 11663
rect 10767 11689 10793 11695
rect 10767 11657 10793 11663
rect 7575 11633 7601 11639
rect 8807 11633 8833 11639
rect 7961 11607 7967 11633
rect 7993 11607 7999 11633
rect 7575 11601 7601 11607
rect 8807 11601 8833 11607
rect 9479 11633 9505 11639
rect 10823 11633 10849 11639
rect 9809 11607 9815 11633
rect 9841 11607 9847 11633
rect 9479 11601 9505 11607
rect 10823 11601 10849 11607
rect 7631 11577 7657 11583
rect 8135 11577 8161 11583
rect 7849 11551 7855 11577
rect 7881 11551 7887 11577
rect 7631 11545 7657 11551
rect 8135 11545 8161 11551
rect 8975 11577 9001 11583
rect 9199 11577 9225 11583
rect 9647 11577 9673 11583
rect 9081 11551 9087 11577
rect 9113 11551 9119 11577
rect 9361 11551 9367 11577
rect 9393 11551 9399 11577
rect 10649 11551 10655 11577
rect 10681 11551 10687 11577
rect 8975 11545 9001 11551
rect 9199 11545 9225 11551
rect 9647 11545 9673 11551
rect 6623 11521 6649 11527
rect 8353 11495 8359 11521
rect 8385 11495 8391 11521
rect 6623 11489 6649 11495
rect 7575 11465 7601 11471
rect 7575 11433 7601 11439
rect 8863 11465 8889 11471
rect 8863 11433 8889 11439
rect 672 11381 20328 11398
rect 672 11355 2239 11381
rect 2265 11355 2291 11381
rect 2317 11355 2343 11381
rect 2369 11355 17599 11381
rect 17625 11355 17651 11381
rect 17677 11355 17703 11381
rect 17729 11355 20328 11381
rect 672 11338 20328 11355
rect 12391 11297 12417 11303
rect 13567 11297 13593 11303
rect 12777 11271 12783 11297
rect 12809 11271 12815 11297
rect 12391 11265 12417 11271
rect 13567 11265 13593 11271
rect 13287 11241 13313 11247
rect 13287 11209 13313 11215
rect 20007 11241 20033 11247
rect 20007 11209 20033 11215
rect 7295 11185 7321 11191
rect 11159 11185 11185 11191
rect 9753 11159 9759 11185
rect 9785 11159 9791 11185
rect 7295 11153 7321 11159
rect 11159 11153 11185 11159
rect 11439 11185 11465 11191
rect 11439 11153 11465 11159
rect 12055 11185 12081 11191
rect 12671 11185 12697 11191
rect 12217 11159 12223 11185
rect 12249 11159 12255 11185
rect 12777 11159 12783 11185
rect 12809 11159 12815 11185
rect 13393 11159 13399 11185
rect 13425 11159 13431 11185
rect 13729 11159 13735 11185
rect 13761 11159 13767 11185
rect 18825 11159 18831 11185
rect 18857 11159 18863 11185
rect 12055 11153 12081 11159
rect 12671 11153 12697 11159
rect 6399 11129 6425 11135
rect 6399 11097 6425 11103
rect 6455 11129 6481 11135
rect 11327 11129 11353 11135
rect 7569 11103 7575 11129
rect 7601 11103 7607 11129
rect 6455 11097 6481 11103
rect 11327 11097 11353 11103
rect 12503 11129 12529 11135
rect 12503 11097 12529 11103
rect 13231 11129 13257 11135
rect 13231 11097 13257 11103
rect 6287 11073 6313 11079
rect 6287 11041 6313 11047
rect 6791 11073 6817 11079
rect 11215 11073 11241 11079
rect 6953 11047 6959 11073
rect 6985 11047 6991 11073
rect 7121 11047 7127 11073
rect 7153 11047 7159 11073
rect 6791 11041 6817 11047
rect 11215 11041 11241 11047
rect 12335 11073 12361 11079
rect 12335 11041 12361 11047
rect 12895 11073 12921 11079
rect 12895 11041 12921 11047
rect 13623 11073 13649 11079
rect 13623 11041 13649 11047
rect 672 10989 20328 11006
rect 672 10963 9919 10989
rect 9945 10963 9971 10989
rect 9997 10963 10023 10989
rect 10049 10963 20328 10989
rect 672 10946 20328 10963
rect 7631 10905 7657 10911
rect 7631 10873 7657 10879
rect 6113 10823 6119 10849
rect 6145 10823 6151 10849
rect 8297 10823 8303 10849
rect 8329 10823 8335 10849
rect 13001 10823 13007 10849
rect 13033 10823 13039 10849
rect 7127 10793 7153 10799
rect 7463 10793 7489 10799
rect 8807 10793 8833 10799
rect 2137 10767 2143 10793
rect 2169 10767 2175 10793
rect 6449 10767 6455 10793
rect 6481 10767 6487 10793
rect 7345 10767 7351 10793
rect 7377 10767 7383 10793
rect 8129 10767 8135 10793
rect 8161 10767 8167 10793
rect 8969 10767 8975 10793
rect 9001 10767 9007 10793
rect 12665 10767 12671 10793
rect 12697 10767 12703 10793
rect 18825 10767 18831 10793
rect 18857 10767 18863 10793
rect 7127 10761 7153 10767
rect 7463 10761 7489 10767
rect 8807 10761 8833 10767
rect 14295 10737 14321 10743
rect 5049 10711 5055 10737
rect 5081 10711 5087 10737
rect 6897 10711 6903 10737
rect 6929 10711 6935 10737
rect 8073 10711 8079 10737
rect 8105 10711 8111 10737
rect 10817 10711 10823 10737
rect 10849 10711 10855 10737
rect 14065 10711 14071 10737
rect 14097 10711 14103 10737
rect 19945 10711 19951 10737
rect 19977 10711 19983 10737
rect 14295 10705 14321 10711
rect 967 10681 993 10687
rect 967 10649 993 10655
rect 672 10597 20328 10614
rect 672 10571 2239 10597
rect 2265 10571 2291 10597
rect 2317 10571 2343 10597
rect 2369 10571 17599 10597
rect 17625 10571 17651 10597
rect 17677 10571 17703 10597
rect 17729 10571 20328 10597
rect 672 10554 20328 10571
rect 7127 10513 7153 10519
rect 9199 10513 9225 10519
rect 8521 10487 8527 10513
rect 8553 10487 8559 10513
rect 7127 10481 7153 10487
rect 9199 10481 9225 10487
rect 9311 10513 9337 10519
rect 9311 10481 9337 10487
rect 7351 10457 7377 10463
rect 20007 10457 20033 10463
rect 4825 10431 4831 10457
rect 4857 10431 4863 10457
rect 8409 10431 8415 10457
rect 8441 10431 8447 10457
rect 9697 10431 9703 10457
rect 9729 10431 9735 10457
rect 9809 10431 9815 10457
rect 9841 10431 9847 10457
rect 7351 10425 7377 10431
rect 20007 10425 20033 10431
rect 6791 10401 6817 10407
rect 6281 10375 6287 10401
rect 6313 10375 6319 10401
rect 6791 10369 6817 10375
rect 6903 10401 6929 10407
rect 6953 10375 6959 10401
rect 6985 10375 6991 10401
rect 7569 10375 7575 10401
rect 7601 10375 7607 10401
rect 8465 10375 8471 10401
rect 8497 10375 8503 10401
rect 8577 10375 8583 10401
rect 8609 10375 8615 10401
rect 9081 10375 9087 10401
rect 9113 10375 9119 10401
rect 9473 10375 9479 10401
rect 9505 10375 9511 10401
rect 9865 10375 9871 10401
rect 9897 10375 9903 10401
rect 10817 10375 10823 10401
rect 10849 10375 10855 10401
rect 18825 10375 18831 10401
rect 18857 10375 18863 10401
rect 6903 10369 6929 10375
rect 7295 10345 7321 10351
rect 9367 10345 9393 10351
rect 5889 10319 5895 10345
rect 5921 10319 5927 10345
rect 7737 10319 7743 10345
rect 7769 10319 7775 10345
rect 7905 10319 7911 10345
rect 7937 10319 7943 10345
rect 13225 10319 13231 10345
rect 13257 10319 13263 10345
rect 7295 10313 7321 10319
rect 9367 10313 9393 10319
rect 6847 10289 6873 10295
rect 7849 10263 7855 10289
rect 7881 10263 7887 10289
rect 6847 10257 6873 10263
rect 672 10205 20328 10222
rect 672 10179 9919 10205
rect 9945 10179 9971 10205
rect 9997 10179 10023 10205
rect 10049 10179 20328 10205
rect 672 10162 20328 10179
rect 6959 10121 6985 10127
rect 6959 10089 6985 10095
rect 6007 10065 6033 10071
rect 6007 10033 6033 10039
rect 6119 10065 6145 10071
rect 6119 10033 6145 10039
rect 6567 10065 6593 10071
rect 6567 10033 6593 10039
rect 6623 10065 6649 10071
rect 8191 10065 8217 10071
rect 7121 10039 7127 10065
rect 7153 10039 7159 10065
rect 7457 10039 7463 10065
rect 7489 10039 7495 10065
rect 6623 10033 6649 10039
rect 8191 10033 8217 10039
rect 8303 10065 8329 10071
rect 11271 10065 11297 10071
rect 14295 10065 14321 10071
rect 8913 10039 8919 10065
rect 8945 10039 8951 10065
rect 9641 10039 9647 10065
rect 9673 10039 9679 10065
rect 10145 10039 10151 10065
rect 10177 10039 10183 10065
rect 11825 10039 11831 10065
rect 11857 10039 11863 10065
rect 8303 10033 8329 10039
rect 11271 10033 11297 10039
rect 14295 10033 14321 10039
rect 11215 10009 11241 10015
rect 7345 9983 7351 10009
rect 7377 9983 7383 10009
rect 7681 9983 7687 10009
rect 7713 9983 7719 10009
rect 8073 9983 8079 10009
rect 8105 9983 8111 10009
rect 8409 9983 8415 10009
rect 8441 9983 8447 10009
rect 9025 9983 9031 10009
rect 9057 9983 9063 10009
rect 9249 9983 9255 10009
rect 9281 9983 9287 10009
rect 10089 9983 10095 10009
rect 10121 9983 10127 10009
rect 11215 9977 11241 9983
rect 11383 10009 11409 10015
rect 11383 9977 11409 9983
rect 11495 10009 11521 10015
rect 11495 9977 11521 9983
rect 11663 10009 11689 10015
rect 12665 9983 12671 10009
rect 12697 9983 12703 10009
rect 11663 9977 11689 9983
rect 6343 9953 6369 9959
rect 5945 9927 5951 9953
rect 5977 9927 5983 9953
rect 6343 9921 6369 9927
rect 7911 9953 7937 9959
rect 8297 9927 8303 9953
rect 8329 9927 8335 9953
rect 10705 9927 10711 9953
rect 10737 9927 10743 9953
rect 13001 9927 13007 9953
rect 13033 9927 13039 9953
rect 14065 9927 14071 9953
rect 14097 9927 14103 9953
rect 7911 9921 7937 9927
rect 6567 9897 6593 9903
rect 6567 9865 6593 9871
rect 672 9813 20328 9830
rect 672 9787 2239 9813
rect 2265 9787 2291 9813
rect 2317 9787 2343 9813
rect 2369 9787 17599 9813
rect 17625 9787 17651 9813
rect 17677 9787 17703 9813
rect 17729 9787 20328 9813
rect 672 9770 20328 9787
rect 7631 9729 7657 9735
rect 9977 9703 9983 9729
rect 10009 9703 10015 9729
rect 12889 9703 12895 9729
rect 12921 9703 12927 9729
rect 7631 9697 7657 9703
rect 8521 9647 8527 9673
rect 8553 9647 8559 9673
rect 9641 9647 9647 9673
rect 9673 9647 9679 9673
rect 11209 9647 11215 9673
rect 11241 9647 11247 9673
rect 12273 9647 12279 9673
rect 12305 9647 12311 9673
rect 7743 9617 7769 9623
rect 7743 9585 7769 9591
rect 7855 9617 7881 9623
rect 9087 9617 9113 9623
rect 10207 9617 10233 9623
rect 8241 9591 8247 9617
rect 8273 9591 8279 9617
rect 8689 9591 8695 9617
rect 8721 9591 8727 9617
rect 9585 9591 9591 9617
rect 9617 9591 9623 9617
rect 9753 9591 9759 9617
rect 9785 9591 9791 9617
rect 10873 9591 10879 9617
rect 10905 9591 10911 9617
rect 12889 9591 12895 9617
rect 12921 9591 12927 9617
rect 7855 9585 7881 9591
rect 9087 9585 9113 9591
rect 10207 9585 10233 9591
rect 8023 9561 8049 9567
rect 12615 9561 12641 9567
rect 8745 9535 8751 9561
rect 8777 9535 8783 9561
rect 12721 9535 12727 9561
rect 12753 9535 12759 9561
rect 8023 9529 8049 9535
rect 12615 9529 12641 9535
rect 7407 9505 7433 9511
rect 7407 9473 7433 9479
rect 9255 9505 9281 9511
rect 13007 9505 13033 9511
rect 10369 9479 10375 9505
rect 10401 9479 10407 9505
rect 9255 9473 9281 9479
rect 13007 9473 13033 9479
rect 13231 9505 13257 9511
rect 13231 9473 13257 9479
rect 672 9421 20328 9438
rect 672 9395 9919 9421
rect 9945 9395 9971 9421
rect 9997 9395 10023 9421
rect 10049 9395 20328 9421
rect 672 9378 20328 9395
rect 10599 9337 10625 9343
rect 7905 9311 7911 9337
rect 7937 9311 7943 9337
rect 10599 9305 10625 9311
rect 10823 9337 10849 9343
rect 10823 9305 10849 9311
rect 7631 9281 7657 9287
rect 6337 9255 6343 9281
rect 6369 9255 6375 9281
rect 7631 9249 7657 9255
rect 7687 9281 7713 9287
rect 7687 9249 7713 9255
rect 8247 9281 8273 9287
rect 8247 9249 8273 9255
rect 10711 9281 10737 9287
rect 10711 9249 10737 9255
rect 12727 9281 12753 9287
rect 12727 9249 12753 9255
rect 12839 9281 12865 9287
rect 12839 9249 12865 9255
rect 6511 9225 6537 9231
rect 2137 9199 2143 9225
rect 2169 9199 2175 9225
rect 6511 9193 6537 9199
rect 7799 9225 7825 9231
rect 7799 9193 7825 9199
rect 8079 9225 8105 9231
rect 8975 9225 9001 9231
rect 8409 9199 8415 9225
rect 8441 9199 8447 9225
rect 8079 9193 8105 9199
rect 8975 9193 9001 9199
rect 9143 9225 9169 9231
rect 9143 9193 9169 9199
rect 9255 9225 9281 9231
rect 9255 9193 9281 9199
rect 9479 9225 9505 9231
rect 9479 9193 9505 9199
rect 9535 9225 9561 9231
rect 9535 9193 9561 9199
rect 9759 9225 9785 9231
rect 10319 9225 10345 9231
rect 10089 9199 10095 9225
rect 10121 9199 10127 9225
rect 10201 9199 10207 9225
rect 10233 9199 10239 9225
rect 9759 9193 9785 9199
rect 10319 9193 10345 9199
rect 10543 9225 10569 9231
rect 10543 9193 10569 9199
rect 13063 9225 13089 9231
rect 13063 9193 13089 9199
rect 9031 9169 9057 9175
rect 9031 9137 9057 9143
rect 9647 9169 9673 9175
rect 9647 9137 9673 9143
rect 10431 9169 10457 9175
rect 10431 9137 10457 9143
rect 12783 9169 12809 9175
rect 12783 9137 12809 9143
rect 967 9113 993 9119
rect 967 9081 993 9087
rect 8415 9113 8441 9119
rect 8415 9081 8441 9087
rect 10879 9113 10905 9119
rect 10879 9081 10905 9087
rect 672 9029 20328 9046
rect 672 9003 2239 9029
rect 2265 9003 2291 9029
rect 2317 9003 2343 9029
rect 2369 9003 17599 9029
rect 17625 9003 17651 9029
rect 17677 9003 17703 9029
rect 17729 9003 20328 9029
rect 672 8986 20328 9003
rect 967 8889 993 8895
rect 9087 8889 9113 8895
rect 14295 8889 14321 8895
rect 8913 8863 8919 8889
rect 8945 8863 8951 8889
rect 13001 8863 13007 8889
rect 13033 8863 13039 8889
rect 14065 8863 14071 8889
rect 14097 8863 14103 8889
rect 967 8857 993 8863
rect 9087 8857 9113 8863
rect 14295 8857 14321 8863
rect 20007 8889 20033 8895
rect 20007 8857 20033 8863
rect 6007 8833 6033 8839
rect 2137 8807 2143 8833
rect 2169 8807 2175 8833
rect 5833 8807 5839 8833
rect 5865 8807 5871 8833
rect 6007 8801 6033 8807
rect 6231 8833 6257 8839
rect 6231 8801 6257 8807
rect 7127 8833 7153 8839
rect 7127 8801 7153 8807
rect 7575 8833 7601 8839
rect 7575 8801 7601 8807
rect 9759 8833 9785 8839
rect 9759 8801 9785 8807
rect 10207 8833 10233 8839
rect 10207 8801 10233 8807
rect 10375 8833 10401 8839
rect 12167 8833 12193 8839
rect 12049 8807 12055 8833
rect 12081 8807 12087 8833
rect 12665 8807 12671 8833
rect 12697 8807 12703 8833
rect 18825 8807 18831 8833
rect 18857 8807 18863 8833
rect 10375 8801 10401 8807
rect 12167 8801 12193 8807
rect 6287 8777 6313 8783
rect 6287 8745 6313 8751
rect 6399 8777 6425 8783
rect 6399 8745 6425 8751
rect 7015 8777 7041 8783
rect 7015 8745 7041 8751
rect 7295 8777 7321 8783
rect 7295 8745 7321 8751
rect 7407 8777 7433 8783
rect 7407 8745 7433 8751
rect 8023 8777 8049 8783
rect 8415 8777 8441 8783
rect 8241 8751 8247 8777
rect 8273 8751 8279 8777
rect 8023 8745 8049 8751
rect 8415 8745 8441 8751
rect 8751 8777 8777 8783
rect 8751 8745 8777 8751
rect 10263 8777 10289 8783
rect 10263 8745 10289 8751
rect 12335 8777 12361 8783
rect 12335 8745 12361 8751
rect 5951 8721 5977 8727
rect 5951 8689 5977 8695
rect 6175 8721 6201 8727
rect 6175 8689 6201 8695
rect 7183 8721 7209 8727
rect 7183 8689 7209 8695
rect 7519 8721 7545 8727
rect 7519 8689 7545 8695
rect 8079 8721 8105 8727
rect 8079 8689 8105 8695
rect 9367 8721 9393 8727
rect 12223 8721 12249 8727
rect 9921 8695 9927 8721
rect 9953 8695 9959 8721
rect 9367 8689 9393 8695
rect 12223 8689 12249 8695
rect 12279 8721 12305 8727
rect 12279 8689 12305 8695
rect 672 8637 20328 8654
rect 672 8611 9919 8637
rect 9945 8611 9971 8637
rect 9997 8611 10023 8637
rect 10049 8611 20328 8637
rect 672 8594 20328 8611
rect 13231 8553 13257 8559
rect 8689 8527 8695 8553
rect 8721 8527 8727 8553
rect 13231 8521 13257 8527
rect 12223 8497 12249 8503
rect 6841 8471 6847 8497
rect 6873 8471 6879 8497
rect 11041 8471 11047 8497
rect 11073 8471 11079 8497
rect 12223 8465 12249 8471
rect 8863 8441 8889 8447
rect 13175 8441 13201 8447
rect 2137 8415 2143 8441
rect 2169 8415 2175 8441
rect 7233 8415 7239 8441
rect 7265 8415 7271 8441
rect 11433 8415 11439 8441
rect 11465 8415 11471 8441
rect 18825 8415 18831 8441
rect 18857 8415 18863 8441
rect 8863 8409 8889 8415
rect 13175 8409 13201 8415
rect 967 8385 993 8391
rect 7463 8385 7489 8391
rect 11663 8385 11689 8391
rect 5777 8359 5783 8385
rect 5809 8359 5815 8385
rect 9977 8359 9983 8385
rect 10009 8359 10015 8385
rect 967 8353 993 8359
rect 7463 8353 7489 8359
rect 11663 8353 11689 8359
rect 20007 8385 20033 8391
rect 20007 8353 20033 8359
rect 12167 8329 12193 8335
rect 12167 8297 12193 8303
rect 13231 8329 13257 8335
rect 13231 8297 13257 8303
rect 672 8245 20328 8262
rect 672 8219 2239 8245
rect 2265 8219 2291 8245
rect 2317 8219 2343 8245
rect 2369 8219 17599 8245
rect 17625 8219 17651 8245
rect 17677 8219 17703 8245
rect 17729 8219 20328 8245
rect 672 8202 20328 8219
rect 10039 8161 10065 8167
rect 10039 8129 10065 8135
rect 4993 8079 4999 8105
rect 5025 8079 5031 8105
rect 6057 8079 6063 8105
rect 6089 8079 6095 8105
rect 12049 8079 12055 8105
rect 12081 8079 12087 8105
rect 13113 8079 13119 8105
rect 13145 8079 13151 8105
rect 10095 8049 10121 8055
rect 6449 8023 6455 8049
rect 6481 8023 6487 8049
rect 10095 8017 10121 8023
rect 10263 8049 10289 8055
rect 11713 8023 11719 8049
rect 11745 8023 11751 8049
rect 10263 8017 10289 8023
rect 8135 7993 8161 7999
rect 8135 7961 8161 7967
rect 8303 7993 8329 7999
rect 10873 7967 10879 7993
rect 10905 7967 10911 7993
rect 8303 7961 8329 7967
rect 6791 7937 6817 7943
rect 6791 7905 6817 7911
rect 10039 7937 10065 7943
rect 10039 7905 10065 7911
rect 10319 7937 10345 7943
rect 10319 7905 10345 7911
rect 10431 7937 10457 7943
rect 10431 7905 10457 7911
rect 10711 7937 10737 7943
rect 10711 7905 10737 7911
rect 13343 7937 13369 7943
rect 13343 7905 13369 7911
rect 672 7853 20328 7870
rect 672 7827 9919 7853
rect 9945 7827 9971 7853
rect 9997 7827 10023 7853
rect 10049 7827 20328 7853
rect 672 7810 20328 7827
rect 12727 7769 12753 7775
rect 12727 7737 12753 7743
rect 12615 7713 12641 7719
rect 7345 7687 7351 7713
rect 7377 7687 7383 7713
rect 10089 7687 10095 7713
rect 10121 7687 10127 7713
rect 12615 7681 12641 7687
rect 8751 7657 8777 7663
rect 10711 7657 10737 7663
rect 7009 7631 7015 7657
rect 7041 7631 7047 7657
rect 10425 7631 10431 7657
rect 10457 7631 10463 7657
rect 8751 7625 8777 7631
rect 10711 7625 10737 7631
rect 12783 7657 12809 7663
rect 12783 7625 12809 7631
rect 12839 7657 12865 7663
rect 12839 7625 12865 7631
rect 12895 7657 12921 7663
rect 12895 7625 12921 7631
rect 13175 7657 13201 7663
rect 13175 7625 13201 7631
rect 13119 7601 13145 7607
rect 8409 7575 8415 7601
rect 8441 7575 8447 7601
rect 9025 7575 9031 7601
rect 9057 7575 9063 7601
rect 13119 7569 13145 7575
rect 672 7461 20328 7478
rect 672 7435 2239 7461
rect 2265 7435 2291 7461
rect 2317 7435 2343 7461
rect 2369 7435 17599 7461
rect 17625 7435 17651 7461
rect 17677 7435 17703 7461
rect 17729 7435 20328 7461
rect 672 7418 20328 7435
rect 8079 7321 8105 7327
rect 13623 7321 13649 7327
rect 8465 7295 8471 7321
rect 8497 7295 8503 7321
rect 12329 7295 12335 7321
rect 12361 7295 12367 7321
rect 13393 7295 13399 7321
rect 13425 7295 13431 7321
rect 8079 7289 8105 7295
rect 13623 7289 13649 7295
rect 10767 7265 10793 7271
rect 8353 7239 8359 7265
rect 8385 7239 8391 7265
rect 10767 7233 10793 7239
rect 10935 7265 10961 7271
rect 11993 7239 11999 7265
rect 12025 7239 12031 7265
rect 10935 7233 10961 7239
rect 10879 7153 10905 7159
rect 10879 7121 10905 7127
rect 672 7069 20328 7086
rect 672 7043 9919 7069
rect 9945 7043 9971 7069
rect 9997 7043 10023 7069
rect 10049 7043 20328 7069
rect 672 7026 20328 7043
rect 11495 6985 11521 6991
rect 11495 6953 11521 6959
rect 10201 6903 10207 6929
rect 10233 6903 10239 6929
rect 9865 6847 9871 6873
rect 9897 6847 9903 6873
rect 11265 6791 11271 6817
rect 11297 6791 11303 6817
rect 672 6677 20328 6694
rect 672 6651 2239 6677
rect 2265 6651 2291 6677
rect 2317 6651 2343 6677
rect 2369 6651 17599 6677
rect 17625 6651 17651 6677
rect 17677 6651 17703 6677
rect 17729 6651 20328 6677
rect 672 6634 20328 6651
rect 672 6285 20328 6302
rect 672 6259 9919 6285
rect 9945 6259 9971 6285
rect 9997 6259 10023 6285
rect 10049 6259 20328 6285
rect 672 6242 20328 6259
rect 672 5893 20328 5910
rect 672 5867 2239 5893
rect 2265 5867 2291 5893
rect 2317 5867 2343 5893
rect 2369 5867 17599 5893
rect 17625 5867 17651 5893
rect 17677 5867 17703 5893
rect 17729 5867 20328 5893
rect 672 5850 20328 5867
rect 672 5501 20328 5518
rect 672 5475 9919 5501
rect 9945 5475 9971 5501
rect 9997 5475 10023 5501
rect 10049 5475 20328 5501
rect 672 5458 20328 5475
rect 672 5109 20328 5126
rect 672 5083 2239 5109
rect 2265 5083 2291 5109
rect 2317 5083 2343 5109
rect 2369 5083 17599 5109
rect 17625 5083 17651 5109
rect 17677 5083 17703 5109
rect 17729 5083 20328 5109
rect 672 5066 20328 5083
rect 672 4717 20328 4734
rect 672 4691 9919 4717
rect 9945 4691 9971 4717
rect 9997 4691 10023 4717
rect 10049 4691 20328 4717
rect 672 4674 20328 4691
rect 672 4325 20328 4342
rect 672 4299 2239 4325
rect 2265 4299 2291 4325
rect 2317 4299 2343 4325
rect 2369 4299 17599 4325
rect 17625 4299 17651 4325
rect 17677 4299 17703 4325
rect 17729 4299 20328 4325
rect 672 4282 20328 4299
rect 672 3933 20328 3950
rect 672 3907 9919 3933
rect 9945 3907 9971 3933
rect 9997 3907 10023 3933
rect 10049 3907 20328 3933
rect 672 3890 20328 3907
rect 672 3541 20328 3558
rect 672 3515 2239 3541
rect 2265 3515 2291 3541
rect 2317 3515 2343 3541
rect 2369 3515 17599 3541
rect 17625 3515 17651 3541
rect 17677 3515 17703 3541
rect 17729 3515 20328 3541
rect 672 3498 20328 3515
rect 672 3149 20328 3166
rect 672 3123 9919 3149
rect 9945 3123 9971 3149
rect 9997 3123 10023 3149
rect 10049 3123 20328 3149
rect 672 3106 20328 3123
rect 672 2757 20328 2774
rect 672 2731 2239 2757
rect 2265 2731 2291 2757
rect 2317 2731 2343 2757
rect 2369 2731 17599 2757
rect 17625 2731 17651 2757
rect 17677 2731 17703 2757
rect 17729 2731 20328 2757
rect 672 2714 20328 2731
rect 672 2365 20328 2382
rect 672 2339 9919 2365
rect 9945 2339 9971 2365
rect 9997 2339 10023 2365
rect 10049 2339 20328 2365
rect 672 2322 20328 2339
rect 10873 2143 10879 2169
rect 10905 2143 10911 2169
rect 11383 2057 11409 2063
rect 11383 2025 11409 2031
rect 672 1973 20328 1990
rect 672 1947 2239 1973
rect 2265 1947 2291 1973
rect 2317 1947 2343 1973
rect 2369 1947 17599 1973
rect 17625 1947 17651 1973
rect 17677 1947 17703 1973
rect 17729 1947 20328 1973
rect 672 1930 20328 1947
rect 12777 1807 12783 1833
rect 12809 1807 12815 1833
rect 10705 1751 10711 1777
rect 10737 1751 10743 1777
rect 13673 1751 13679 1777
rect 13705 1751 13711 1777
rect 3823 1665 3849 1671
rect 3823 1633 3849 1639
rect 11215 1665 11241 1671
rect 11215 1633 11241 1639
rect 672 1581 20328 1598
rect 672 1555 9919 1581
rect 9945 1555 9971 1581
rect 9997 1555 10023 1581
rect 10049 1555 20328 1581
rect 672 1538 20328 1555
<< via1 >>
rect 2239 19195 2265 19221
rect 2291 19195 2317 19221
rect 2343 19195 2369 19221
rect 17599 19195 17625 19221
rect 17651 19195 17677 19221
rect 17703 19195 17729 19221
rect 9311 19111 9337 19137
rect 11215 19111 11241 19137
rect 12783 19111 12809 19137
rect 9031 18999 9057 19025
rect 10711 18999 10737 19025
rect 12279 18999 12305 19025
rect 10375 18943 10401 18969
rect 9919 18803 9945 18829
rect 9971 18803 9997 18829
rect 10023 18803 10049 18829
rect 9199 18719 9225 18745
rect 11047 18719 11073 18745
rect 13119 18719 13145 18745
rect 20119 18663 20145 18689
rect 8695 18607 8721 18633
rect 10543 18607 10569 18633
rect 12615 18607 12641 18633
rect 2239 18411 2265 18437
rect 2291 18411 2317 18437
rect 2343 18411 2369 18437
rect 17599 18411 17625 18437
rect 17651 18411 17677 18437
rect 17703 18411 17729 18437
rect 9919 18019 9945 18045
rect 9971 18019 9997 18045
rect 10023 18019 10049 18045
rect 2239 17627 2265 17653
rect 2291 17627 2317 17653
rect 2343 17627 2369 17653
rect 17599 17627 17625 17653
rect 17651 17627 17677 17653
rect 17703 17627 17729 17653
rect 9919 17235 9945 17261
rect 9971 17235 9997 17261
rect 10023 17235 10049 17261
rect 2239 16843 2265 16869
rect 2291 16843 2317 16869
rect 2343 16843 2369 16869
rect 17599 16843 17625 16869
rect 17651 16843 17677 16869
rect 17703 16843 17729 16869
rect 9919 16451 9945 16477
rect 9971 16451 9997 16477
rect 10023 16451 10049 16477
rect 2239 16059 2265 16085
rect 2291 16059 2317 16085
rect 2343 16059 2369 16085
rect 17599 16059 17625 16085
rect 17651 16059 17677 16085
rect 17703 16059 17729 16085
rect 9919 15667 9945 15693
rect 9971 15667 9997 15693
rect 10023 15667 10049 15693
rect 2239 15275 2265 15301
rect 2291 15275 2317 15301
rect 2343 15275 2369 15301
rect 17599 15275 17625 15301
rect 17651 15275 17677 15301
rect 17703 15275 17729 15301
rect 9919 14883 9945 14909
rect 9971 14883 9997 14909
rect 10023 14883 10049 14909
rect 2239 14491 2265 14517
rect 2291 14491 2317 14517
rect 2343 14491 2369 14517
rect 17599 14491 17625 14517
rect 17651 14491 17677 14517
rect 17703 14491 17729 14517
rect 9919 14099 9945 14125
rect 9971 14099 9997 14125
rect 10023 14099 10049 14125
rect 8975 13903 9001 13929
rect 10767 13903 10793 13929
rect 18943 13903 18969 13929
rect 8863 13847 8889 13873
rect 9367 13847 9393 13873
rect 10431 13847 10457 13873
rect 11159 13847 11185 13873
rect 12223 13847 12249 13873
rect 12727 13847 12753 13873
rect 19951 13847 19977 13873
rect 2239 13707 2265 13733
rect 2291 13707 2317 13733
rect 2343 13707 2369 13733
rect 17599 13707 17625 13733
rect 17651 13707 17677 13733
rect 17703 13707 17729 13733
rect 8527 13567 8553 13593
rect 20007 13567 20033 13593
rect 7071 13511 7097 13537
rect 8751 13511 8777 13537
rect 9367 13511 9393 13537
rect 10151 13511 10177 13537
rect 11271 13511 11297 13537
rect 11831 13511 11857 13537
rect 13791 13511 13817 13537
rect 18831 13511 18857 13537
rect 7463 13455 7489 13481
rect 8695 13455 8721 13481
rect 9087 13455 9113 13481
rect 9479 13455 9505 13481
rect 9535 13455 9561 13481
rect 9983 13455 10009 13481
rect 10095 13455 10121 13481
rect 11383 13455 11409 13481
rect 11439 13455 11465 13481
rect 11663 13455 11689 13481
rect 11775 13455 11801 13481
rect 13175 13455 13201 13481
rect 13231 13455 13257 13481
rect 13903 13455 13929 13481
rect 8807 13399 8833 13425
rect 13063 13399 13089 13425
rect 9919 13315 9945 13341
rect 9971 13315 9997 13341
rect 10023 13315 10049 13341
rect 8191 13231 8217 13257
rect 8303 13175 8329 13201
rect 14407 13175 14433 13201
rect 8135 13119 8161 13145
rect 8415 13119 8441 13145
rect 8695 13119 8721 13145
rect 8807 13119 8833 13145
rect 8919 13119 8945 13145
rect 9031 13119 9057 13145
rect 12615 13119 12641 13145
rect 14295 13119 14321 13145
rect 18831 13119 18857 13145
rect 6567 13063 6593 13089
rect 13007 13063 13033 13089
rect 14071 13063 14097 13089
rect 14631 13063 14657 13089
rect 19951 13063 19977 13089
rect 2239 12923 2265 12949
rect 2291 12923 2317 12949
rect 2343 12923 2369 12949
rect 17599 12923 17625 12949
rect 17651 12923 17677 12949
rect 17703 12923 17729 12949
rect 967 12783 993 12809
rect 4999 12783 5025 12809
rect 8191 12783 8217 12809
rect 9255 12783 9281 12809
rect 9479 12783 9505 12809
rect 12167 12783 12193 12809
rect 14015 12783 14041 12809
rect 20007 12783 20033 12809
rect 2143 12727 2169 12753
rect 6455 12727 6481 12753
rect 7855 12727 7881 12753
rect 10767 12727 10793 12753
rect 12559 12727 12585 12753
rect 18831 12727 18857 12753
rect 6063 12671 6089 12697
rect 6959 12671 6985 12697
rect 9983 12671 10009 12697
rect 11103 12671 11129 12697
rect 12951 12671 12977 12697
rect 6791 12615 6817 12641
rect 6903 12615 6929 12641
rect 7015 12615 7041 12641
rect 9815 12615 9841 12641
rect 12391 12615 12417 12641
rect 14239 12615 14265 12641
rect 9919 12531 9945 12557
rect 9971 12531 9997 12557
rect 10023 12531 10049 12557
rect 8807 12447 8833 12473
rect 8863 12447 8889 12473
rect 8919 12447 8945 12473
rect 11775 12447 11801 12473
rect 12783 12447 12809 12473
rect 13231 12447 13257 12473
rect 13511 12447 13537 12473
rect 13623 12447 13649 12473
rect 7631 12391 7657 12417
rect 7687 12391 7713 12417
rect 12895 12391 12921 12417
rect 12951 12391 12977 12417
rect 13455 12391 13481 12417
rect 6007 12335 6033 12361
rect 8751 12335 8777 12361
rect 9031 12335 9057 12361
rect 11271 12335 11297 12361
rect 11495 12335 11521 12361
rect 11663 12335 11689 12361
rect 11887 12335 11913 12361
rect 13175 12335 13201 12361
rect 6343 12279 6369 12305
rect 7407 12279 7433 12305
rect 7911 12279 7937 12305
rect 9871 12279 9897 12305
rect 10935 12279 10961 12305
rect 11719 12279 11745 12305
rect 7631 12223 7657 12249
rect 13231 12223 13257 12249
rect 2239 12139 2265 12165
rect 2291 12139 2317 12165
rect 2343 12139 2369 12165
rect 17599 12139 17625 12165
rect 17651 12139 17677 12165
rect 17703 12139 17729 12165
rect 6399 12055 6425 12081
rect 10655 12055 10681 12081
rect 6791 11999 6817 12025
rect 11719 11999 11745 12025
rect 6847 11943 6873 11969
rect 7071 11943 7097 11969
rect 10711 11943 10737 11969
rect 10991 11943 11017 11969
rect 6399 11887 6425 11913
rect 6455 11887 6481 11913
rect 8135 11887 8161 11913
rect 10823 11887 10849 11913
rect 11103 11887 11129 11913
rect 11439 11887 11465 11913
rect 11495 11887 11521 11913
rect 6735 11831 6761 11857
rect 8191 11831 8217 11857
rect 11047 11831 11073 11857
rect 11383 11831 11409 11857
rect 9919 11747 9945 11773
rect 9971 11747 9997 11773
rect 10023 11747 10049 11773
rect 9535 11663 9561 11689
rect 10767 11663 10793 11689
rect 7575 11607 7601 11633
rect 7967 11607 7993 11633
rect 8807 11607 8833 11633
rect 9479 11607 9505 11633
rect 9815 11607 9841 11633
rect 10823 11607 10849 11633
rect 7631 11551 7657 11577
rect 7855 11551 7881 11577
rect 8135 11551 8161 11577
rect 8975 11551 9001 11577
rect 9087 11551 9113 11577
rect 9199 11551 9225 11577
rect 9367 11551 9393 11577
rect 9647 11551 9673 11577
rect 10655 11551 10681 11577
rect 6623 11495 6649 11521
rect 8359 11495 8385 11521
rect 7575 11439 7601 11465
rect 8863 11439 8889 11465
rect 2239 11355 2265 11381
rect 2291 11355 2317 11381
rect 2343 11355 2369 11381
rect 17599 11355 17625 11381
rect 17651 11355 17677 11381
rect 17703 11355 17729 11381
rect 12391 11271 12417 11297
rect 12783 11271 12809 11297
rect 13567 11271 13593 11297
rect 13287 11215 13313 11241
rect 20007 11215 20033 11241
rect 7295 11159 7321 11185
rect 9759 11159 9785 11185
rect 11159 11159 11185 11185
rect 11439 11159 11465 11185
rect 12055 11159 12081 11185
rect 12223 11159 12249 11185
rect 12671 11159 12697 11185
rect 12783 11159 12809 11185
rect 13399 11159 13425 11185
rect 13735 11159 13761 11185
rect 18831 11159 18857 11185
rect 6399 11103 6425 11129
rect 6455 11103 6481 11129
rect 7575 11103 7601 11129
rect 11327 11103 11353 11129
rect 12503 11103 12529 11129
rect 13231 11103 13257 11129
rect 6287 11047 6313 11073
rect 6791 11047 6817 11073
rect 6959 11047 6985 11073
rect 7127 11047 7153 11073
rect 11215 11047 11241 11073
rect 12335 11047 12361 11073
rect 12895 11047 12921 11073
rect 13623 11047 13649 11073
rect 9919 10963 9945 10989
rect 9971 10963 9997 10989
rect 10023 10963 10049 10989
rect 7631 10879 7657 10905
rect 6119 10823 6145 10849
rect 8303 10823 8329 10849
rect 13007 10823 13033 10849
rect 2143 10767 2169 10793
rect 6455 10767 6481 10793
rect 7127 10767 7153 10793
rect 7351 10767 7377 10793
rect 7463 10767 7489 10793
rect 8135 10767 8161 10793
rect 8807 10767 8833 10793
rect 8975 10767 9001 10793
rect 12671 10767 12697 10793
rect 18831 10767 18857 10793
rect 5055 10711 5081 10737
rect 6903 10711 6929 10737
rect 8079 10711 8105 10737
rect 10823 10711 10849 10737
rect 14071 10711 14097 10737
rect 14295 10711 14321 10737
rect 19951 10711 19977 10737
rect 967 10655 993 10681
rect 2239 10571 2265 10597
rect 2291 10571 2317 10597
rect 2343 10571 2369 10597
rect 17599 10571 17625 10597
rect 17651 10571 17677 10597
rect 17703 10571 17729 10597
rect 7127 10487 7153 10513
rect 8527 10487 8553 10513
rect 9199 10487 9225 10513
rect 9311 10487 9337 10513
rect 4831 10431 4857 10457
rect 7351 10431 7377 10457
rect 8415 10431 8441 10457
rect 9703 10431 9729 10457
rect 9815 10431 9841 10457
rect 20007 10431 20033 10457
rect 6287 10375 6313 10401
rect 6791 10375 6817 10401
rect 6903 10375 6929 10401
rect 6959 10375 6985 10401
rect 7575 10375 7601 10401
rect 8471 10375 8497 10401
rect 8583 10375 8609 10401
rect 9087 10375 9113 10401
rect 9479 10375 9505 10401
rect 9871 10375 9897 10401
rect 10823 10375 10849 10401
rect 18831 10375 18857 10401
rect 5895 10319 5921 10345
rect 7295 10319 7321 10345
rect 7743 10319 7769 10345
rect 7911 10319 7937 10345
rect 9367 10319 9393 10345
rect 13231 10319 13257 10345
rect 6847 10263 6873 10289
rect 7855 10263 7881 10289
rect 9919 10179 9945 10205
rect 9971 10179 9997 10205
rect 10023 10179 10049 10205
rect 6959 10095 6985 10121
rect 6007 10039 6033 10065
rect 6119 10039 6145 10065
rect 6567 10039 6593 10065
rect 6623 10039 6649 10065
rect 7127 10039 7153 10065
rect 7463 10039 7489 10065
rect 8191 10039 8217 10065
rect 8303 10039 8329 10065
rect 8919 10039 8945 10065
rect 9647 10039 9673 10065
rect 10151 10039 10177 10065
rect 11271 10039 11297 10065
rect 11831 10039 11857 10065
rect 14295 10039 14321 10065
rect 7351 9983 7377 10009
rect 7687 9983 7713 10009
rect 8079 9983 8105 10009
rect 8415 9983 8441 10009
rect 9031 9983 9057 10009
rect 9255 9983 9281 10009
rect 10095 9983 10121 10009
rect 11215 9983 11241 10009
rect 11383 9983 11409 10009
rect 11495 9983 11521 10009
rect 11663 9983 11689 10009
rect 12671 9983 12697 10009
rect 5951 9927 5977 9953
rect 6343 9927 6369 9953
rect 7911 9927 7937 9953
rect 8303 9927 8329 9953
rect 10711 9927 10737 9953
rect 13007 9927 13033 9953
rect 14071 9927 14097 9953
rect 6567 9871 6593 9897
rect 2239 9787 2265 9813
rect 2291 9787 2317 9813
rect 2343 9787 2369 9813
rect 17599 9787 17625 9813
rect 17651 9787 17677 9813
rect 17703 9787 17729 9813
rect 7631 9703 7657 9729
rect 9983 9703 10009 9729
rect 12895 9703 12921 9729
rect 8527 9647 8553 9673
rect 9647 9647 9673 9673
rect 11215 9647 11241 9673
rect 12279 9647 12305 9673
rect 7743 9591 7769 9617
rect 7855 9591 7881 9617
rect 8247 9591 8273 9617
rect 8695 9591 8721 9617
rect 9087 9591 9113 9617
rect 9591 9591 9617 9617
rect 9759 9591 9785 9617
rect 10207 9591 10233 9617
rect 10879 9591 10905 9617
rect 12895 9591 12921 9617
rect 8023 9535 8049 9561
rect 8751 9535 8777 9561
rect 12615 9535 12641 9561
rect 12727 9535 12753 9561
rect 7407 9479 7433 9505
rect 9255 9479 9281 9505
rect 10375 9479 10401 9505
rect 13007 9479 13033 9505
rect 13231 9479 13257 9505
rect 9919 9395 9945 9421
rect 9971 9395 9997 9421
rect 10023 9395 10049 9421
rect 7911 9311 7937 9337
rect 10599 9311 10625 9337
rect 10823 9311 10849 9337
rect 6343 9255 6369 9281
rect 7631 9255 7657 9281
rect 7687 9255 7713 9281
rect 8247 9255 8273 9281
rect 10711 9255 10737 9281
rect 12727 9255 12753 9281
rect 12839 9255 12865 9281
rect 2143 9199 2169 9225
rect 6511 9199 6537 9225
rect 7799 9199 7825 9225
rect 8079 9199 8105 9225
rect 8415 9199 8441 9225
rect 8975 9199 9001 9225
rect 9143 9199 9169 9225
rect 9255 9199 9281 9225
rect 9479 9199 9505 9225
rect 9535 9199 9561 9225
rect 9759 9199 9785 9225
rect 10095 9199 10121 9225
rect 10207 9199 10233 9225
rect 10319 9199 10345 9225
rect 10543 9199 10569 9225
rect 13063 9199 13089 9225
rect 9031 9143 9057 9169
rect 9647 9143 9673 9169
rect 10431 9143 10457 9169
rect 12783 9143 12809 9169
rect 967 9087 993 9113
rect 8415 9087 8441 9113
rect 10879 9087 10905 9113
rect 2239 9003 2265 9029
rect 2291 9003 2317 9029
rect 2343 9003 2369 9029
rect 17599 9003 17625 9029
rect 17651 9003 17677 9029
rect 17703 9003 17729 9029
rect 967 8863 993 8889
rect 8919 8863 8945 8889
rect 9087 8863 9113 8889
rect 13007 8863 13033 8889
rect 14071 8863 14097 8889
rect 14295 8863 14321 8889
rect 20007 8863 20033 8889
rect 2143 8807 2169 8833
rect 5839 8807 5865 8833
rect 6007 8807 6033 8833
rect 6231 8807 6257 8833
rect 7127 8807 7153 8833
rect 7575 8807 7601 8833
rect 9759 8807 9785 8833
rect 10207 8807 10233 8833
rect 10375 8807 10401 8833
rect 12055 8807 12081 8833
rect 12167 8807 12193 8833
rect 12671 8807 12697 8833
rect 18831 8807 18857 8833
rect 6287 8751 6313 8777
rect 6399 8751 6425 8777
rect 7015 8751 7041 8777
rect 7295 8751 7321 8777
rect 7407 8751 7433 8777
rect 8023 8751 8049 8777
rect 8247 8751 8273 8777
rect 8415 8751 8441 8777
rect 8751 8751 8777 8777
rect 10263 8751 10289 8777
rect 12335 8751 12361 8777
rect 5951 8695 5977 8721
rect 6175 8695 6201 8721
rect 7183 8695 7209 8721
rect 7519 8695 7545 8721
rect 8079 8695 8105 8721
rect 9367 8695 9393 8721
rect 9927 8695 9953 8721
rect 12223 8695 12249 8721
rect 12279 8695 12305 8721
rect 9919 8611 9945 8637
rect 9971 8611 9997 8637
rect 10023 8611 10049 8637
rect 8695 8527 8721 8553
rect 13231 8527 13257 8553
rect 6847 8471 6873 8497
rect 11047 8471 11073 8497
rect 12223 8471 12249 8497
rect 2143 8415 2169 8441
rect 7239 8415 7265 8441
rect 8863 8415 8889 8441
rect 11439 8415 11465 8441
rect 13175 8415 13201 8441
rect 18831 8415 18857 8441
rect 967 8359 993 8385
rect 5783 8359 5809 8385
rect 7463 8359 7489 8385
rect 9983 8359 10009 8385
rect 11663 8359 11689 8385
rect 20007 8359 20033 8385
rect 12167 8303 12193 8329
rect 13231 8303 13257 8329
rect 2239 8219 2265 8245
rect 2291 8219 2317 8245
rect 2343 8219 2369 8245
rect 17599 8219 17625 8245
rect 17651 8219 17677 8245
rect 17703 8219 17729 8245
rect 10039 8135 10065 8161
rect 4999 8079 5025 8105
rect 6063 8079 6089 8105
rect 12055 8079 12081 8105
rect 13119 8079 13145 8105
rect 6455 8023 6481 8049
rect 10095 8023 10121 8049
rect 10263 8023 10289 8049
rect 11719 8023 11745 8049
rect 8135 7967 8161 7993
rect 8303 7967 8329 7993
rect 10879 7967 10905 7993
rect 6791 7911 6817 7937
rect 10039 7911 10065 7937
rect 10319 7911 10345 7937
rect 10431 7911 10457 7937
rect 10711 7911 10737 7937
rect 13343 7911 13369 7937
rect 9919 7827 9945 7853
rect 9971 7827 9997 7853
rect 10023 7827 10049 7853
rect 12727 7743 12753 7769
rect 7351 7687 7377 7713
rect 10095 7687 10121 7713
rect 12615 7687 12641 7713
rect 7015 7631 7041 7657
rect 8751 7631 8777 7657
rect 10431 7631 10457 7657
rect 10711 7631 10737 7657
rect 12783 7631 12809 7657
rect 12839 7631 12865 7657
rect 12895 7631 12921 7657
rect 13175 7631 13201 7657
rect 8415 7575 8441 7601
rect 9031 7575 9057 7601
rect 13119 7575 13145 7601
rect 2239 7435 2265 7461
rect 2291 7435 2317 7461
rect 2343 7435 2369 7461
rect 17599 7435 17625 7461
rect 17651 7435 17677 7461
rect 17703 7435 17729 7461
rect 8079 7295 8105 7321
rect 8471 7295 8497 7321
rect 12335 7295 12361 7321
rect 13399 7295 13425 7321
rect 13623 7295 13649 7321
rect 8359 7239 8385 7265
rect 10767 7239 10793 7265
rect 10935 7239 10961 7265
rect 11999 7239 12025 7265
rect 10879 7127 10905 7153
rect 9919 7043 9945 7069
rect 9971 7043 9997 7069
rect 10023 7043 10049 7069
rect 11495 6959 11521 6985
rect 10207 6903 10233 6929
rect 9871 6847 9897 6873
rect 11271 6791 11297 6817
rect 2239 6651 2265 6677
rect 2291 6651 2317 6677
rect 2343 6651 2369 6677
rect 17599 6651 17625 6677
rect 17651 6651 17677 6677
rect 17703 6651 17729 6677
rect 9919 6259 9945 6285
rect 9971 6259 9997 6285
rect 10023 6259 10049 6285
rect 2239 5867 2265 5893
rect 2291 5867 2317 5893
rect 2343 5867 2369 5893
rect 17599 5867 17625 5893
rect 17651 5867 17677 5893
rect 17703 5867 17729 5893
rect 9919 5475 9945 5501
rect 9971 5475 9997 5501
rect 10023 5475 10049 5501
rect 2239 5083 2265 5109
rect 2291 5083 2317 5109
rect 2343 5083 2369 5109
rect 17599 5083 17625 5109
rect 17651 5083 17677 5109
rect 17703 5083 17729 5109
rect 9919 4691 9945 4717
rect 9971 4691 9997 4717
rect 10023 4691 10049 4717
rect 2239 4299 2265 4325
rect 2291 4299 2317 4325
rect 2343 4299 2369 4325
rect 17599 4299 17625 4325
rect 17651 4299 17677 4325
rect 17703 4299 17729 4325
rect 9919 3907 9945 3933
rect 9971 3907 9997 3933
rect 10023 3907 10049 3933
rect 2239 3515 2265 3541
rect 2291 3515 2317 3541
rect 2343 3515 2369 3541
rect 17599 3515 17625 3541
rect 17651 3515 17677 3541
rect 17703 3515 17729 3541
rect 9919 3123 9945 3149
rect 9971 3123 9997 3149
rect 10023 3123 10049 3149
rect 2239 2731 2265 2757
rect 2291 2731 2317 2757
rect 2343 2731 2369 2757
rect 17599 2731 17625 2757
rect 17651 2731 17677 2757
rect 17703 2731 17729 2757
rect 9919 2339 9945 2365
rect 9971 2339 9997 2365
rect 10023 2339 10049 2365
rect 10879 2143 10905 2169
rect 11383 2031 11409 2057
rect 2239 1947 2265 1973
rect 2291 1947 2317 1973
rect 2343 1947 2369 1973
rect 17599 1947 17625 1973
rect 17651 1947 17677 1973
rect 17703 1947 17729 1973
rect 12783 1807 12809 1833
rect 10711 1751 10737 1777
rect 13679 1751 13705 1777
rect 3823 1639 3849 1665
rect 11215 1639 11241 1665
rect 9919 1555 9945 1581
rect 9971 1555 9997 1581
rect 10023 1555 10049 1581
<< metal2 >>
rect 8400 20600 8456 21000
rect 9072 20600 9128 21000
rect 9408 20600 9464 21000
rect 10416 20600 10472 21000
rect 11088 20600 11144 21000
rect 11760 20600 11816 21000
rect 12096 20600 12152 21000
rect 2238 19222 2370 19227
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2238 19189 2370 19194
rect 8414 18746 8442 20600
rect 9086 19138 9114 20600
rect 9310 19138 9338 19143
rect 9086 19137 9338 19138
rect 9086 19111 9311 19137
rect 9337 19111 9338 19137
rect 9086 19110 9338 19111
rect 9310 19105 9338 19110
rect 8414 18713 8442 18718
rect 9030 19025 9058 19031
rect 9030 18999 9031 19025
rect 9057 18999 9058 19025
rect 8694 18633 8722 18639
rect 8694 18607 8695 18633
rect 8721 18607 8722 18633
rect 2238 18438 2370 18443
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2238 18405 2370 18410
rect 2238 17654 2370 17659
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2238 17621 2370 17626
rect 2238 16870 2370 16875
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2238 16837 2370 16842
rect 2238 16086 2370 16091
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2238 16053 2370 16058
rect 8694 15974 8722 18607
rect 8526 15946 8722 15974
rect 9030 15974 9058 18999
rect 9422 18970 9450 20600
rect 9422 18937 9450 18942
rect 10374 18970 10402 18975
rect 10374 18923 10402 18942
rect 9918 18830 10050 18835
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 9918 18797 10050 18802
rect 9198 18746 9226 18751
rect 9198 18699 9226 18718
rect 10430 18746 10458 20600
rect 11102 19138 11130 20600
rect 11214 19138 11242 19143
rect 11102 19137 11242 19138
rect 11102 19111 11215 19137
rect 11241 19111 11242 19137
rect 11102 19110 11242 19111
rect 11214 19105 11242 19110
rect 11774 19138 11802 20600
rect 11774 19105 11802 19110
rect 10430 18713 10458 18718
rect 10710 19025 10738 19031
rect 10710 18999 10711 19025
rect 10737 18999 10738 19025
rect 10542 18633 10570 18639
rect 10542 18607 10543 18633
rect 10569 18607 10570 18633
rect 9918 18046 10050 18051
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 9918 18013 10050 18018
rect 9918 17262 10050 17267
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 9918 17229 10050 17234
rect 9918 16478 10050 16483
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 9918 16445 10050 16450
rect 10542 15974 10570 18607
rect 10710 15974 10738 18999
rect 11046 18746 11074 18751
rect 11046 18699 11074 18718
rect 12110 18746 12138 20600
rect 17598 19222 17730 19227
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17598 19189 17730 19194
rect 12782 19138 12810 19143
rect 12782 19091 12810 19110
rect 12110 18713 12138 18718
rect 12278 19025 12306 19031
rect 12278 18999 12279 19025
rect 12305 18999 12306 19025
rect 12278 15974 12306 18999
rect 13118 18746 13146 18751
rect 13118 18699 13146 18718
rect 20118 18689 20146 18695
rect 20118 18663 20119 18689
rect 20145 18663 20146 18689
rect 9030 15946 9226 15974
rect 2238 15302 2370 15307
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2238 15269 2370 15274
rect 2238 14518 2370 14523
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2238 14485 2370 14490
rect 2086 13818 2114 13823
rect 966 12809 994 12815
rect 966 12783 967 12809
rect 993 12783 994 12809
rect 966 12474 994 12783
rect 966 12441 994 12446
rect 2086 10738 2114 13790
rect 2238 13734 2370 13739
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2238 13701 2370 13706
rect 8526 13593 8554 15946
rect 8974 13929 9002 13935
rect 8974 13903 8975 13929
rect 9001 13903 9002 13929
rect 8526 13567 8527 13593
rect 8553 13567 8554 13593
rect 7070 13537 7098 13543
rect 7070 13511 7071 13537
rect 7097 13511 7098 13537
rect 6566 13482 6594 13487
rect 6566 13089 6594 13454
rect 7070 13482 7098 13511
rect 8246 13538 8274 13543
rect 7070 13449 7098 13454
rect 7462 13481 7490 13487
rect 7462 13455 7463 13481
rect 7489 13455 7490 13481
rect 7462 13258 7490 13455
rect 7462 13225 7490 13230
rect 8190 13258 8218 13263
rect 8190 13211 8218 13230
rect 8134 13146 8162 13151
rect 8134 13099 8162 13118
rect 6566 13063 6567 13089
rect 6593 13063 6594 13089
rect 2238 12950 2370 12955
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2238 12917 2370 12922
rect 4998 12810 5026 12815
rect 4998 12763 5026 12782
rect 5950 12810 5978 12815
rect 2142 12754 2170 12759
rect 2142 12707 2170 12726
rect 2238 12166 2370 12171
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2238 12133 2370 12138
rect 5950 11914 5978 12782
rect 6454 12754 6482 12759
rect 6566 12754 6594 13063
rect 8190 12810 8218 12815
rect 8246 12810 8274 13510
rect 8526 13426 8554 13567
rect 8862 13874 8890 13879
rect 8974 13874 9002 13903
rect 8862 13873 9002 13874
rect 8862 13847 8863 13873
rect 8889 13847 9002 13873
rect 8862 13846 9002 13847
rect 8750 13538 8778 13543
rect 8750 13491 8778 13510
rect 8694 13482 8722 13487
rect 8526 13393 8554 13398
rect 8638 13481 8722 13482
rect 8638 13455 8695 13481
rect 8721 13455 8722 13481
rect 8638 13454 8722 13455
rect 8302 13202 8330 13207
rect 8302 13155 8330 13174
rect 8190 12809 8274 12810
rect 8190 12783 8191 12809
rect 8217 12783 8274 12809
rect 8190 12782 8274 12783
rect 8414 13146 8442 13151
rect 8638 13146 8666 13454
rect 8694 13449 8722 13454
rect 8862 13482 8890 13846
rect 8862 13449 8890 13454
rect 9086 13482 9114 13487
rect 9086 13435 9114 13454
rect 9198 13454 9226 15946
rect 10430 15946 10570 15974
rect 10654 15946 10738 15974
rect 12222 15946 12306 15974
rect 12614 18633 12642 18639
rect 12614 18607 12615 18633
rect 12641 18607 12642 18633
rect 9918 15694 10050 15699
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 9918 15661 10050 15666
rect 9918 14910 10050 14915
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 9918 14877 10050 14882
rect 9918 14126 10050 14131
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 9918 14093 10050 14098
rect 9366 13873 9394 13879
rect 10430 13874 10458 15946
rect 9366 13847 9367 13873
rect 9393 13847 9394 13873
rect 9366 13537 9394 13847
rect 9366 13511 9367 13537
rect 9393 13511 9394 13537
rect 9366 13505 9394 13511
rect 10094 13873 10458 13874
rect 10094 13847 10431 13873
rect 10457 13847 10458 13873
rect 10094 13846 10458 13847
rect 9478 13481 9506 13487
rect 9478 13455 9479 13481
rect 9505 13455 9506 13481
rect 8750 13426 8778 13431
rect 8414 13145 8666 13146
rect 8414 13119 8415 13145
rect 8441 13119 8666 13145
rect 8414 13118 8666 13119
rect 8694 13145 8722 13151
rect 8694 13119 8695 13145
rect 8721 13119 8722 13145
rect 8190 12777 8218 12782
rect 6118 12753 6594 12754
rect 6118 12727 6455 12753
rect 6481 12727 6594 12753
rect 6118 12726 6594 12727
rect 7854 12754 7882 12759
rect 7854 12753 7938 12754
rect 7854 12727 7855 12753
rect 7881 12727 7938 12753
rect 7854 12726 7938 12727
rect 6062 12698 6090 12703
rect 6062 12651 6090 12670
rect 6006 12362 6034 12367
rect 6118 12362 6146 12726
rect 6454 12721 6482 12726
rect 6006 12361 6146 12362
rect 6006 12335 6007 12361
rect 6033 12335 6146 12361
rect 6006 12334 6146 12335
rect 6454 12642 6482 12647
rect 6006 12329 6034 12334
rect 6342 12306 6370 12311
rect 6342 12259 6370 12278
rect 6398 12082 6426 12087
rect 6454 12082 6482 12614
rect 6398 12081 6482 12082
rect 6398 12055 6399 12081
rect 6425 12055 6482 12081
rect 6398 12054 6482 12055
rect 6398 12049 6426 12054
rect 6398 11914 6426 11919
rect 5950 11913 6426 11914
rect 5950 11887 6399 11913
rect 6425 11887 6426 11913
rect 5950 11886 6426 11887
rect 6398 11881 6426 11886
rect 6454 11913 6482 11919
rect 6454 11887 6455 11913
rect 6481 11887 6482 11913
rect 2238 11382 2370 11387
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2238 11349 2370 11354
rect 6454 11298 6482 11887
rect 6510 11522 6538 12726
rect 7854 12721 7882 12726
rect 6958 12698 6986 12703
rect 6958 12651 6986 12670
rect 6790 12642 6818 12647
rect 6790 12595 6818 12614
rect 6902 12641 6930 12647
rect 6902 12615 6903 12641
rect 6929 12615 6930 12641
rect 6790 12306 6818 12311
rect 6790 12025 6818 12278
rect 6790 11999 6791 12025
rect 6817 11999 6818 12025
rect 6790 11993 6818 11999
rect 6902 12026 6930 12615
rect 6846 11970 6874 11975
rect 6902 11970 6930 11998
rect 6846 11969 6930 11970
rect 6846 11943 6847 11969
rect 6873 11943 6930 11969
rect 6846 11942 6930 11943
rect 7014 12641 7042 12647
rect 7014 12615 7015 12641
rect 7041 12615 7042 12641
rect 7014 12418 7042 12615
rect 6846 11937 6874 11942
rect 6734 11858 6762 11863
rect 7014 11858 7042 12390
rect 7630 12417 7658 12423
rect 7630 12391 7631 12417
rect 7657 12391 7658 12417
rect 7630 12362 7658 12391
rect 7686 12418 7714 12423
rect 7686 12371 7714 12390
rect 7630 12329 7658 12334
rect 7406 12305 7434 12311
rect 7406 12279 7407 12305
rect 7433 12279 7434 12305
rect 7070 12250 7098 12255
rect 7070 11969 7098 12222
rect 7070 11943 7071 11969
rect 7097 11943 7098 11969
rect 7070 11937 7098 11943
rect 6734 11857 7042 11858
rect 6734 11831 6735 11857
rect 6761 11831 7042 11857
rect 6734 11830 7042 11831
rect 6734 11802 6762 11830
rect 6678 11774 6762 11802
rect 7406 11802 7434 12279
rect 7910 12305 7938 12726
rect 7910 12279 7911 12305
rect 7937 12279 7938 12305
rect 7630 12250 7658 12255
rect 7630 12203 7658 12222
rect 6622 11522 6650 11527
rect 6510 11521 6650 11522
rect 6510 11495 6623 11521
rect 6649 11495 6650 11521
rect 6510 11494 6650 11495
rect 6454 11270 6594 11298
rect 6398 11130 6426 11135
rect 6398 11083 6426 11102
rect 6454 11130 6482 11135
rect 6454 11129 6538 11130
rect 6454 11103 6455 11129
rect 6481 11103 6538 11129
rect 6454 11102 6538 11103
rect 6454 11097 6482 11102
rect 6286 11074 6314 11079
rect 6118 11073 6314 11074
rect 6118 11047 6287 11073
rect 6313 11047 6314 11073
rect 6118 11046 6314 11047
rect 6118 10849 6146 11046
rect 6286 11041 6314 11046
rect 6118 10823 6119 10849
rect 6145 10823 6146 10849
rect 6118 10817 6146 10823
rect 6454 11018 6482 11023
rect 2142 10794 2170 10799
rect 2142 10747 2170 10766
rect 4830 10794 4858 10799
rect 2086 10705 2114 10710
rect 966 10681 994 10687
rect 966 10655 967 10681
rect 993 10655 994 10681
rect 966 10458 994 10655
rect 2238 10598 2370 10603
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2238 10565 2370 10570
rect 966 10425 994 10430
rect 4830 10457 4858 10766
rect 6454 10793 6482 10990
rect 6454 10767 6455 10793
rect 6481 10767 6482 10793
rect 4830 10431 4831 10457
rect 4857 10431 4858 10457
rect 4830 10402 4858 10431
rect 4830 10369 4858 10374
rect 5054 10737 5082 10743
rect 5054 10711 5055 10737
rect 5081 10711 5082 10737
rect 5054 10122 5082 10711
rect 6286 10401 6314 10407
rect 6286 10375 6287 10401
rect 6313 10375 6314 10401
rect 5054 10089 5082 10094
rect 5894 10345 5922 10351
rect 5894 10319 5895 10345
rect 5921 10319 5922 10345
rect 5894 10094 5922 10319
rect 6118 10290 6146 10295
rect 5894 10066 5978 10094
rect 5950 9953 5978 10066
rect 5950 9927 5951 9953
rect 5977 9927 5978 9953
rect 5950 9921 5978 9927
rect 6006 10065 6034 10071
rect 6006 10039 6007 10065
rect 6033 10039 6034 10065
rect 2238 9814 2370 9819
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2238 9781 2370 9786
rect 2142 9226 2170 9231
rect 2142 9179 2170 9198
rect 4998 9226 5026 9231
rect 966 9114 994 9119
rect 966 9067 994 9086
rect 2238 9030 2370 9035
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2238 8997 2370 9002
rect 966 8890 994 8895
rect 966 8843 994 8862
rect 2142 8834 2170 8839
rect 2142 8787 2170 8806
rect 4998 8778 5026 9198
rect 5894 9002 5922 9007
rect 6006 9002 6034 10039
rect 6118 10065 6146 10262
rect 6118 10039 6119 10065
rect 6145 10039 6146 10065
rect 6118 10033 6146 10039
rect 6286 9954 6314 10375
rect 6342 9954 6370 9959
rect 6454 9954 6482 10767
rect 6286 9953 6482 9954
rect 6286 9927 6343 9953
rect 6369 9927 6482 9953
rect 6286 9926 6482 9927
rect 6342 9921 6370 9926
rect 6398 9842 6426 9847
rect 5922 8974 6034 9002
rect 6342 9281 6370 9287
rect 6342 9255 6343 9281
rect 6369 9255 6370 9281
rect 5838 8834 5866 8839
rect 5894 8834 5922 8974
rect 5838 8833 5922 8834
rect 5838 8807 5839 8833
rect 5865 8807 5922 8833
rect 5838 8806 5922 8807
rect 6006 8834 6034 8839
rect 6230 8834 6258 8839
rect 6006 8833 6258 8834
rect 6006 8807 6007 8833
rect 6033 8807 6231 8833
rect 6257 8807 6258 8833
rect 6006 8806 6258 8807
rect 5838 8801 5866 8806
rect 6006 8801 6034 8806
rect 6230 8801 6258 8806
rect 6342 8834 6370 9255
rect 6342 8801 6370 8806
rect 966 8442 994 8447
rect 966 8385 994 8414
rect 2142 8442 2170 8447
rect 2142 8395 2170 8414
rect 966 8359 967 8385
rect 993 8359 994 8385
rect 966 8353 994 8359
rect 2238 8246 2370 8251
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2238 8213 2370 8218
rect 4998 8105 5026 8750
rect 6286 8778 6314 8783
rect 6286 8731 6314 8750
rect 6398 8777 6426 9814
rect 6398 8751 6399 8777
rect 6425 8751 6426 8777
rect 6398 8745 6426 8751
rect 5782 8722 5810 8727
rect 5782 8442 5810 8694
rect 5782 8385 5810 8414
rect 5782 8359 5783 8385
rect 5809 8359 5810 8385
rect 5782 8353 5810 8359
rect 5950 8721 5978 8727
rect 5950 8695 5951 8721
rect 5977 8695 5978 8721
rect 4998 8079 4999 8105
rect 5025 8079 5026 8105
rect 4998 8073 5026 8079
rect 5950 8106 5978 8695
rect 6174 8721 6202 8727
rect 6174 8695 6175 8721
rect 6201 8695 6202 8721
rect 6174 8666 6202 8695
rect 6174 8633 6202 8638
rect 6062 8106 6090 8111
rect 5950 8105 6090 8106
rect 5950 8079 6063 8105
rect 6089 8079 6090 8105
rect 5950 8078 6090 8079
rect 6062 8073 6090 8078
rect 6454 8050 6482 9926
rect 6510 9898 6538 11102
rect 6566 10962 6594 11270
rect 6622 11018 6650 11494
rect 6622 10985 6650 10990
rect 6566 10929 6594 10934
rect 6678 10738 6706 11774
rect 7294 11186 7322 11191
rect 7294 11139 7322 11158
rect 6790 11073 6818 11079
rect 6790 11047 6791 11073
rect 6817 11047 6818 11073
rect 6790 10906 6818 11047
rect 6790 10873 6818 10878
rect 6958 11073 6986 11079
rect 6958 11047 6959 11073
rect 6985 11047 6986 11073
rect 6622 10710 6706 10738
rect 6902 10737 6930 10743
rect 6902 10711 6903 10737
rect 6929 10711 6930 10737
rect 6622 10682 6650 10710
rect 6566 10065 6594 10071
rect 6566 10039 6567 10065
rect 6593 10039 6594 10065
rect 6566 10010 6594 10039
rect 6622 10065 6650 10654
rect 6902 10626 6930 10711
rect 6902 10593 6930 10598
rect 6790 10458 6818 10463
rect 6790 10401 6818 10430
rect 6790 10375 6791 10401
rect 6817 10375 6818 10401
rect 6790 10369 6818 10375
rect 6902 10402 6930 10407
rect 6902 10355 6930 10374
rect 6958 10402 6986 11047
rect 7126 11074 7154 11079
rect 7126 11027 7154 11046
rect 7126 10962 7154 10967
rect 7070 10934 7126 10962
rect 7406 10962 7434 11774
rect 7518 12026 7546 12031
rect 7462 11634 7490 11639
rect 7462 11074 7490 11606
rect 7518 11466 7546 11998
rect 7854 11914 7882 11919
rect 7574 11634 7602 11639
rect 7574 11587 7602 11606
rect 7630 11578 7658 11583
rect 7630 11577 7770 11578
rect 7630 11551 7631 11577
rect 7657 11551 7770 11577
rect 7630 11550 7770 11551
rect 7630 11545 7658 11550
rect 7574 11466 7602 11471
rect 7518 11465 7602 11466
rect 7518 11439 7575 11465
rect 7601 11439 7602 11465
rect 7518 11438 7602 11439
rect 7574 11433 7602 11438
rect 7462 11041 7490 11046
rect 7574 11129 7602 11135
rect 7574 11103 7575 11129
rect 7601 11103 7602 11129
rect 7574 11018 7602 11103
rect 7574 10985 7602 10990
rect 7686 11074 7714 11079
rect 7406 10934 7490 10962
rect 7070 10514 7098 10934
rect 7126 10929 7154 10934
rect 7126 10794 7154 10799
rect 7350 10794 7378 10799
rect 7126 10793 7434 10794
rect 7126 10767 7127 10793
rect 7153 10767 7351 10793
rect 7377 10767 7434 10793
rect 7126 10766 7434 10767
rect 7126 10761 7154 10766
rect 7350 10761 7378 10766
rect 7126 10514 7154 10519
rect 7070 10513 7154 10514
rect 7070 10487 7127 10513
rect 7153 10487 7154 10513
rect 7070 10486 7154 10487
rect 7126 10481 7154 10486
rect 7350 10458 7378 10463
rect 7350 10411 7378 10430
rect 6958 10401 7042 10402
rect 6958 10375 6959 10401
rect 6985 10375 7042 10401
rect 6958 10374 7042 10375
rect 6958 10369 6986 10374
rect 6846 10290 6874 10295
rect 6846 10243 6874 10262
rect 6958 10122 6986 10141
rect 6958 10089 6986 10094
rect 6622 10039 6623 10065
rect 6649 10039 6650 10065
rect 6622 10033 6650 10039
rect 7014 10066 7042 10374
rect 7294 10346 7322 10351
rect 7294 10122 7322 10318
rect 7406 10094 7434 10766
rect 7462 10793 7490 10934
rect 7462 10767 7463 10793
rect 7489 10767 7490 10793
rect 7462 10761 7490 10767
rect 7630 10906 7658 10911
rect 7294 10089 7322 10094
rect 7014 10033 7042 10038
rect 7126 10065 7154 10071
rect 7126 10039 7127 10065
rect 7153 10039 7154 10065
rect 7126 10010 7154 10039
rect 7350 10066 7434 10094
rect 7574 10402 7602 10407
rect 7630 10402 7658 10878
rect 7574 10401 7658 10402
rect 7574 10375 7575 10401
rect 7601 10375 7658 10401
rect 7574 10374 7658 10375
rect 7350 10010 7378 10066
rect 7126 10009 7378 10010
rect 7126 9983 7351 10009
rect 7377 9983 7378 10009
rect 7126 9982 7378 9983
rect 6566 9977 6594 9982
rect 6566 9898 6594 9903
rect 6510 9897 6594 9898
rect 6510 9871 6567 9897
rect 6593 9871 6594 9897
rect 6510 9870 6594 9871
rect 6566 9865 6594 9870
rect 7350 9730 7378 9982
rect 7350 9697 7378 9702
rect 7462 10065 7490 10071
rect 7462 10039 7463 10065
rect 7489 10039 7490 10065
rect 7462 10010 7490 10039
rect 7462 9674 7490 9982
rect 7490 9646 7546 9674
rect 7462 9641 7490 9646
rect 7406 9505 7434 9511
rect 7406 9479 7407 9505
rect 7433 9479 7434 9505
rect 6510 9225 6538 9231
rect 6510 9199 6511 9225
rect 6537 9199 6538 9225
rect 6510 8778 6538 9199
rect 7126 9226 7154 9231
rect 6510 8745 6538 8750
rect 7014 9170 7042 9175
rect 7014 8777 7042 9142
rect 7126 8833 7154 9198
rect 7406 9226 7434 9479
rect 7518 9226 7546 9646
rect 7574 9282 7602 10374
rect 7686 10122 7714 11046
rect 7742 10626 7770 11550
rect 7854 11577 7882 11886
rect 7854 11551 7855 11577
rect 7881 11551 7882 11577
rect 7854 11545 7882 11551
rect 7742 10593 7770 10598
rect 7854 11130 7882 11135
rect 7630 10094 7714 10122
rect 7742 10345 7770 10351
rect 7742 10319 7743 10345
rect 7769 10319 7770 10345
rect 7630 9842 7658 10094
rect 7686 10010 7714 10015
rect 7742 10010 7770 10319
rect 7854 10289 7882 11102
rect 7910 11018 7938 12279
rect 8134 11914 8162 11919
rect 8134 11867 8162 11886
rect 8190 11857 8218 11863
rect 8190 11831 8191 11857
rect 8217 11831 8218 11857
rect 7910 10985 7938 10990
rect 7966 11633 7994 11639
rect 7966 11607 7967 11633
rect 7993 11607 7994 11633
rect 7966 10794 7994 11607
rect 8134 11578 8162 11583
rect 8190 11578 8218 11831
rect 8414 11634 8442 13118
rect 8694 12530 8722 13119
rect 8750 13146 8778 13398
rect 8806 13425 8834 13431
rect 9198 13426 9282 13454
rect 8806 13399 8807 13425
rect 8833 13399 8834 13425
rect 8806 13258 8834 13399
rect 8806 13230 8890 13258
rect 8806 13146 8834 13151
rect 8750 13145 8834 13146
rect 8750 13119 8807 13145
rect 8833 13119 8834 13145
rect 8750 13118 8834 13119
rect 8806 13113 8834 13118
rect 8526 12502 8834 12530
rect 8470 11634 8498 11639
rect 8414 11606 8470 11634
rect 8470 11601 8498 11606
rect 8134 11577 8218 11578
rect 8134 11551 8135 11577
rect 8161 11551 8218 11577
rect 8134 11550 8218 11551
rect 8134 11186 8162 11550
rect 8134 11153 8162 11158
rect 8358 11521 8386 11527
rect 8358 11495 8359 11521
rect 8385 11495 8386 11521
rect 8190 10962 8218 10967
rect 7966 10761 7994 10766
rect 8134 10793 8162 10799
rect 8134 10767 8135 10793
rect 8161 10767 8162 10793
rect 8078 10737 8106 10743
rect 8078 10711 8079 10737
rect 8105 10711 8106 10737
rect 8078 10682 8106 10711
rect 8078 10649 8106 10654
rect 7854 10263 7855 10289
rect 7881 10263 7882 10289
rect 7854 10257 7882 10263
rect 7910 10346 7938 10351
rect 7910 10066 7938 10318
rect 8134 10122 8162 10767
rect 7686 10009 7770 10010
rect 7686 9983 7687 10009
rect 7713 9983 7770 10009
rect 7686 9982 7770 9983
rect 7686 9977 7714 9982
rect 7630 9814 7714 9842
rect 7630 9730 7658 9735
rect 7630 9683 7658 9702
rect 7686 9562 7714 9814
rect 7686 9394 7714 9534
rect 7742 9617 7770 9982
rect 7742 9591 7743 9617
rect 7769 9591 7770 9617
rect 7742 9506 7770 9591
rect 7854 10038 7938 10066
rect 8022 10094 8162 10122
rect 7854 9618 7882 10038
rect 7910 9954 7938 9959
rect 8022 9954 8050 10094
rect 8190 10066 8218 10934
rect 8302 10850 8330 10855
rect 8302 10803 8330 10822
rect 8358 10682 8386 11495
rect 8414 10794 8442 10799
rect 8442 10766 8498 10794
rect 8414 10761 8442 10766
rect 8358 10649 8386 10654
rect 8470 10570 8498 10766
rect 8190 10019 8218 10038
rect 8246 10458 8274 10463
rect 7910 9953 8022 9954
rect 7910 9927 7911 9953
rect 7937 9927 8022 9953
rect 7910 9926 8022 9927
rect 7910 9921 7938 9926
rect 8022 9907 8050 9926
rect 8078 10009 8106 10015
rect 8078 9983 8079 10009
rect 8105 9983 8106 10009
rect 7854 9571 7882 9590
rect 8022 9562 8050 9567
rect 8022 9515 8050 9534
rect 7742 9473 7770 9478
rect 8078 9450 8106 9983
rect 8246 9730 8274 10430
rect 8414 10458 8442 10463
rect 8414 10411 8442 10430
rect 8470 10401 8498 10542
rect 8470 10375 8471 10401
rect 8497 10375 8498 10401
rect 8470 10369 8498 10375
rect 8526 10513 8554 12502
rect 8806 12473 8834 12502
rect 8806 12447 8807 12473
rect 8833 12447 8834 12473
rect 8806 12441 8834 12447
rect 8862 12473 8890 13230
rect 8918 13146 8946 13151
rect 8918 13099 8946 13118
rect 9030 13145 9058 13151
rect 9030 13119 9031 13145
rect 9057 13119 9058 13145
rect 8862 12447 8863 12473
rect 8889 12447 8890 12473
rect 8862 12441 8890 12447
rect 8918 12810 8946 12815
rect 8918 12473 8946 12782
rect 8918 12447 8919 12473
rect 8945 12447 8946 12473
rect 8918 12441 8946 12447
rect 8750 12361 8778 12367
rect 8750 12335 8751 12361
rect 8777 12335 8778 12361
rect 8582 11466 8610 11471
rect 8582 10962 8610 11438
rect 8582 10929 8610 10934
rect 8526 10487 8527 10513
rect 8553 10487 8554 10513
rect 8526 10290 8554 10487
rect 8582 10401 8610 10407
rect 8582 10375 8583 10401
rect 8609 10375 8610 10401
rect 8582 10346 8610 10375
rect 8582 10313 8610 10318
rect 8414 10262 8554 10290
rect 8302 10066 8330 10071
rect 8302 10019 8330 10038
rect 8414 10009 8442 10262
rect 8750 10066 8778 12335
rect 9030 12362 9058 13119
rect 9254 12810 9282 13426
rect 9422 13426 9450 13431
rect 9422 12810 9450 13398
rect 9478 13202 9506 13455
rect 9534 13482 9562 13487
rect 9982 13482 10010 13487
rect 9534 13481 10010 13482
rect 9534 13455 9535 13481
rect 9561 13455 9983 13481
rect 10009 13455 10010 13481
rect 9534 13454 10010 13455
rect 9534 13449 9562 13454
rect 9982 13449 10010 13454
rect 10094 13481 10122 13846
rect 10430 13841 10458 13846
rect 10094 13455 10095 13481
rect 10121 13455 10122 13481
rect 10094 13449 10122 13455
rect 10150 13538 10178 13543
rect 9918 13342 10050 13347
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 10150 13314 10178 13510
rect 9918 13309 10050 13314
rect 10094 13286 10178 13314
rect 10094 13258 10122 13286
rect 9982 13230 10122 13258
rect 9506 13174 9562 13202
rect 9478 13155 9506 13174
rect 9478 12810 9506 12815
rect 9422 12809 9506 12810
rect 9422 12783 9479 12809
rect 9505 12783 9506 12809
rect 9422 12782 9506 12783
rect 9254 12763 9282 12782
rect 9478 12777 9506 12782
rect 9030 12315 9058 12334
rect 8974 11746 9002 11751
rect 8806 11634 8834 11639
rect 8806 11587 8834 11606
rect 8974 11578 9002 11718
rect 9534 11689 9562 13174
rect 9982 12697 10010 13230
rect 9982 12671 9983 12697
rect 10009 12671 10010 12697
rect 9982 12665 10010 12671
rect 9814 12641 9842 12647
rect 9814 12615 9815 12641
rect 9841 12615 9842 12641
rect 9758 12362 9786 12367
rect 9534 11663 9535 11689
rect 9561 11663 9562 11689
rect 9534 11657 9562 11663
rect 9702 11970 9730 11975
rect 9478 11633 9506 11639
rect 9478 11607 9479 11633
rect 9505 11607 9506 11633
rect 9086 11578 9114 11583
rect 8974 11577 9058 11578
rect 8974 11551 8975 11577
rect 9001 11551 9058 11577
rect 8974 11550 9058 11551
rect 8974 11545 9002 11550
rect 8862 11466 8890 11471
rect 8862 11419 8890 11438
rect 9030 10962 9058 11550
rect 9086 11577 9170 11578
rect 9086 11551 9087 11577
rect 9113 11551 9170 11577
rect 9086 11550 9170 11551
rect 9086 11545 9114 11550
rect 8806 10794 8834 10799
rect 8974 10794 9002 10799
rect 8806 10793 9002 10794
rect 8806 10767 8807 10793
rect 8833 10767 8975 10793
rect 9001 10767 9002 10793
rect 8806 10766 9002 10767
rect 8806 10738 8834 10766
rect 8974 10761 9002 10766
rect 8806 10705 8834 10710
rect 9030 10682 9058 10934
rect 8694 10038 8750 10066
rect 8414 9983 8415 10009
rect 8441 9983 8442 10009
rect 8414 9977 8442 9983
rect 8470 10010 8498 10015
rect 8302 9953 8330 9959
rect 8302 9927 8303 9953
rect 8329 9927 8330 9953
rect 8302 9842 8330 9927
rect 8302 9809 8330 9814
rect 8190 9702 8274 9730
rect 8022 9422 8106 9450
rect 8134 9506 8162 9511
rect 7686 9366 7770 9394
rect 7630 9282 7658 9287
rect 7574 9281 7658 9282
rect 7574 9255 7631 9281
rect 7657 9255 7658 9281
rect 7574 9254 7658 9255
rect 7630 9249 7658 9254
rect 7686 9282 7714 9287
rect 7686 9235 7714 9254
rect 7518 9198 7602 9226
rect 7406 9193 7434 9198
rect 7126 8807 7127 8833
rect 7153 8807 7154 8833
rect 7126 8801 7154 8807
rect 7574 8833 7602 9198
rect 7742 9170 7770 9366
rect 7910 9338 7938 9343
rect 7910 9291 7938 9310
rect 7742 9137 7770 9142
rect 7798 9225 7826 9231
rect 7798 9199 7799 9225
rect 7825 9199 7826 9225
rect 7798 8946 7826 9199
rect 7798 8913 7826 8918
rect 8022 8890 8050 9422
rect 8078 9225 8106 9231
rect 8078 9199 8079 9225
rect 8105 9199 8106 9225
rect 8078 9170 8106 9199
rect 8134 9170 8162 9478
rect 8190 9282 8218 9702
rect 8246 9617 8274 9623
rect 8246 9591 8247 9617
rect 8273 9591 8274 9617
rect 8246 9394 8274 9591
rect 8246 9366 8386 9394
rect 8246 9282 8274 9287
rect 8190 9281 8274 9282
rect 8190 9255 8247 9281
rect 8273 9255 8274 9281
rect 8190 9254 8274 9255
rect 8246 9249 8274 9254
rect 8078 9142 8274 9170
rect 8022 8862 8162 8890
rect 7574 8807 7575 8833
rect 7601 8807 7602 8833
rect 7574 8801 7602 8807
rect 7014 8751 7015 8777
rect 7041 8751 7042 8777
rect 7014 8666 7042 8751
rect 7294 8778 7322 8783
rect 7406 8778 7434 8783
rect 7294 8777 7434 8778
rect 7294 8751 7295 8777
rect 7321 8751 7407 8777
rect 7433 8751 7434 8777
rect 7294 8750 7434 8751
rect 7294 8745 7322 8750
rect 7406 8745 7434 8750
rect 8022 8778 8050 8783
rect 7014 8633 7042 8638
rect 7182 8721 7210 8727
rect 7182 8695 7183 8721
rect 7209 8695 7210 8721
rect 7182 8554 7210 8695
rect 7518 8722 7546 8727
rect 7518 8675 7546 8694
rect 6846 8526 7210 8554
rect 8022 8554 8050 8750
rect 8078 8722 8106 8727
rect 8078 8675 8106 8694
rect 6846 8497 6874 8526
rect 8022 8521 8050 8526
rect 6846 8471 6847 8497
rect 6873 8471 6874 8497
rect 6846 8465 6874 8471
rect 7238 8441 7266 8447
rect 7238 8415 7239 8441
rect 7265 8415 7266 8441
rect 7238 8386 7266 8415
rect 7462 8386 7490 8391
rect 7238 8385 7490 8386
rect 7238 8359 7463 8385
rect 7489 8359 7490 8385
rect 7238 8358 7490 8359
rect 6454 8003 6482 8022
rect 6790 8050 6818 8055
rect 6790 7937 6818 8022
rect 6790 7911 6791 7937
rect 6817 7911 6818 7937
rect 6790 7658 6818 7911
rect 7350 7994 7378 7999
rect 7350 7713 7378 7966
rect 7350 7687 7351 7713
rect 7377 7687 7378 7713
rect 7350 7681 7378 7687
rect 7014 7658 7042 7663
rect 6790 7630 7014 7658
rect 7014 7611 7042 7630
rect 7462 7658 7490 8358
rect 8134 7994 8162 8862
rect 8246 8777 8274 9142
rect 8246 8751 8247 8777
rect 8273 8751 8274 8777
rect 8246 8745 8274 8751
rect 8302 8722 8330 8727
rect 8358 8722 8386 9366
rect 8414 9226 8442 9231
rect 8470 9226 8498 9982
rect 8526 9674 8554 9679
rect 8526 9627 8554 9646
rect 8694 9617 8722 10038
rect 8750 10033 8778 10038
rect 8918 10654 9058 10682
rect 8918 10065 8946 10654
rect 9086 10570 9114 10575
rect 9030 10542 9086 10570
rect 9030 10290 9058 10542
rect 9086 10537 9114 10542
rect 9086 10402 9114 10407
rect 9086 10355 9114 10374
rect 9030 10262 9114 10290
rect 8918 10039 8919 10065
rect 8945 10039 8946 10065
rect 8918 10033 8946 10039
rect 8974 10066 9002 10071
rect 8694 9591 8695 9617
rect 8721 9591 8722 9617
rect 8694 9338 8722 9591
rect 8750 9562 8778 9567
rect 8750 9515 8778 9534
rect 8694 9305 8722 9310
rect 8974 9226 9002 10038
rect 9030 10009 9058 10015
rect 9030 9983 9031 10009
rect 9057 9983 9058 10009
rect 9030 9282 9058 9983
rect 9086 9617 9114 10262
rect 9086 9591 9087 9617
rect 9113 9591 9114 9617
rect 9086 9585 9114 9591
rect 9142 9394 9170 11550
rect 9198 11577 9226 11583
rect 9198 11551 9199 11577
rect 9225 11551 9226 11577
rect 9198 11466 9226 11551
rect 9198 11433 9226 11438
rect 9366 11577 9394 11583
rect 9366 11551 9367 11577
rect 9393 11551 9394 11577
rect 9198 10682 9226 10687
rect 9198 10513 9226 10654
rect 9198 10487 9199 10513
rect 9225 10487 9226 10513
rect 9198 10010 9226 10487
rect 9310 10514 9338 10519
rect 9366 10514 9394 11551
rect 9478 10850 9506 11607
rect 9310 10513 9394 10514
rect 9310 10487 9311 10513
rect 9337 10487 9394 10513
rect 9310 10486 9394 10487
rect 9422 10822 9478 10850
rect 9310 10066 9338 10486
rect 9310 10033 9338 10038
rect 9366 10345 9394 10351
rect 9366 10319 9367 10345
rect 9393 10319 9394 10345
rect 9254 10010 9282 10015
rect 9226 10009 9282 10010
rect 9226 9983 9255 10009
rect 9281 9983 9282 10009
rect 9226 9982 9282 9983
rect 9198 9963 9226 9982
rect 9254 9977 9282 9982
rect 9366 9618 9394 10319
rect 9422 9898 9450 10822
rect 9478 10817 9506 10822
rect 9646 11577 9674 11583
rect 9646 11551 9647 11577
rect 9673 11551 9674 11577
rect 9478 10570 9506 10575
rect 9646 10570 9674 11551
rect 9506 10542 9674 10570
rect 9478 10401 9506 10542
rect 9478 10375 9479 10401
rect 9505 10375 9506 10401
rect 9478 10369 9506 10375
rect 9646 10458 9674 10463
rect 9646 10065 9674 10430
rect 9702 10457 9730 11942
rect 9758 11634 9786 12334
rect 9814 11746 9842 12615
rect 9918 12558 10050 12563
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 9918 12525 10050 12530
rect 9870 12306 9898 12311
rect 9870 12259 9898 12278
rect 10654 12306 10682 15946
rect 10766 13929 10794 13935
rect 10766 13903 10767 13929
rect 10793 13903 10794 13929
rect 10766 12754 10794 13903
rect 11158 13874 11186 13879
rect 12222 13874 12250 15946
rect 11158 13873 11298 13874
rect 11158 13847 11159 13873
rect 11185 13847 11298 13873
rect 11158 13846 11298 13847
rect 11158 13841 11186 13846
rect 11270 13537 11298 13846
rect 11270 13511 11271 13537
rect 11297 13511 11298 13537
rect 11270 13505 11298 13511
rect 11774 13873 12250 13874
rect 11774 13847 12223 13873
rect 12249 13847 12250 13873
rect 11774 13846 12250 13847
rect 11382 13481 11410 13487
rect 11382 13455 11383 13481
rect 11409 13455 11410 13481
rect 10766 12707 10794 12726
rect 11270 12754 11298 12759
rect 11102 12698 11130 12703
rect 11102 12697 11186 12698
rect 11102 12671 11103 12697
rect 11129 12671 11186 12697
rect 11102 12670 11186 12671
rect 11102 12665 11130 12670
rect 10934 12306 10962 12311
rect 10654 12081 10682 12278
rect 10654 12055 10655 12081
rect 10681 12055 10682 12081
rect 10654 12049 10682 12055
rect 10766 12305 10962 12306
rect 10766 12279 10935 12305
rect 10961 12279 10962 12305
rect 10766 12278 10962 12279
rect 10710 11970 10738 11975
rect 10710 11923 10738 11942
rect 10542 11858 10570 11863
rect 9918 11774 10050 11779
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 9918 11741 10050 11746
rect 9814 11713 9842 11718
rect 9814 11634 9842 11639
rect 9758 11633 9842 11634
rect 9758 11607 9815 11633
rect 9841 11607 9842 11633
rect 9758 11606 9842 11607
rect 9758 11185 9786 11191
rect 9758 11159 9759 11185
rect 9785 11159 9786 11185
rect 9758 10738 9786 11159
rect 9814 10906 9842 11606
rect 10542 11130 10570 11830
rect 10710 11802 10738 11807
rect 10542 11097 10570 11102
rect 10654 11577 10682 11583
rect 10654 11551 10655 11577
rect 10681 11551 10682 11577
rect 10654 11186 10682 11551
rect 9918 10990 10050 10995
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 9918 10957 10050 10962
rect 9814 10873 9842 10878
rect 9758 10705 9786 10710
rect 9702 10431 9703 10457
rect 9729 10431 9730 10457
rect 9702 10425 9730 10431
rect 9814 10626 9842 10631
rect 9814 10458 9842 10598
rect 9814 10411 9842 10430
rect 9870 10401 9898 10407
rect 9870 10375 9871 10401
rect 9897 10375 9898 10401
rect 9870 10346 9898 10375
rect 9646 10039 9647 10065
rect 9673 10039 9674 10065
rect 9590 10010 9618 10015
rect 9450 9870 9562 9898
rect 9422 9865 9450 9870
rect 9366 9585 9394 9590
rect 9254 9505 9282 9511
rect 9254 9479 9255 9505
rect 9281 9479 9282 9505
rect 9142 9366 9226 9394
rect 9030 9254 9114 9282
rect 8414 9225 8498 9226
rect 8414 9199 8415 9225
rect 8441 9199 8498 9225
rect 8414 9198 8498 9199
rect 8918 9225 9002 9226
rect 8918 9199 8975 9225
rect 9001 9199 9002 9225
rect 8918 9198 9002 9199
rect 8414 9193 8442 9198
rect 8414 9114 8442 9119
rect 8414 9067 8442 9086
rect 8918 8889 8946 9198
rect 8974 9193 9002 9198
rect 9030 9169 9058 9175
rect 9030 9143 9031 9169
rect 9057 9143 9058 9169
rect 9030 9002 9058 9143
rect 9086 9114 9114 9254
rect 9086 9081 9114 9086
rect 9142 9225 9170 9231
rect 9142 9199 9143 9225
rect 9169 9199 9170 9225
rect 9030 8969 9058 8974
rect 8918 8863 8919 8889
rect 8945 8863 8946 8889
rect 8918 8857 8946 8863
rect 9086 8890 9114 8895
rect 9086 8843 9114 8862
rect 8330 8694 8386 8722
rect 8414 8778 8442 8783
rect 8302 8689 8330 8694
rect 8134 7947 8162 7966
rect 8302 7993 8330 7999
rect 8302 7967 8303 7993
rect 8329 7967 8330 7993
rect 7462 7625 7490 7630
rect 8302 7574 8330 7967
rect 8190 7546 8330 7574
rect 8358 7602 8386 7607
rect 2238 7462 2370 7467
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2238 7429 2370 7434
rect 8078 7322 8106 7327
rect 8190 7322 8218 7546
rect 8078 7321 8218 7322
rect 8078 7295 8079 7321
rect 8105 7295 8218 7321
rect 8078 7294 8218 7295
rect 8078 7289 8106 7294
rect 8358 7265 8386 7574
rect 8414 7601 8442 8750
rect 8750 8778 8778 8783
rect 8750 8731 8778 8750
rect 9142 8722 9170 9199
rect 9198 9058 9226 9366
rect 9254 9226 9282 9479
rect 9478 9226 9506 9231
rect 9254 9225 9506 9226
rect 9254 9199 9255 9225
rect 9281 9199 9479 9225
rect 9505 9199 9506 9225
rect 9254 9198 9506 9199
rect 9254 9193 9282 9198
rect 9478 9170 9506 9198
rect 9478 9137 9506 9142
rect 9534 9225 9562 9870
rect 9590 9617 9618 9982
rect 9646 9673 9674 10039
rect 9646 9647 9647 9673
rect 9673 9647 9674 9673
rect 9646 9641 9674 9647
rect 9758 10318 9898 10346
rect 9758 9954 9786 10318
rect 9918 10206 10050 10211
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 9918 10173 10050 10178
rect 10094 10066 10122 10071
rect 10094 10009 10122 10038
rect 10094 9983 10095 10009
rect 10121 9983 10122 10009
rect 10094 9977 10122 9983
rect 10150 10065 10178 10071
rect 10150 10039 10151 10065
rect 10177 10039 10178 10065
rect 9590 9591 9591 9617
rect 9617 9591 9618 9617
rect 9590 9585 9618 9591
rect 9758 9617 9786 9926
rect 10150 9898 10178 10039
rect 10150 9865 10178 9870
rect 10318 10010 10346 10015
rect 9982 9730 10010 9735
rect 9982 9683 10010 9702
rect 10318 9730 10346 9982
rect 9758 9591 9759 9617
rect 9785 9591 9786 9617
rect 9534 9199 9535 9225
rect 9561 9199 9562 9225
rect 9198 9025 9226 9030
rect 9534 8890 9562 9199
rect 9758 9225 9786 9591
rect 10206 9618 10234 9623
rect 10206 9571 10234 9590
rect 9918 9422 10050 9427
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 9918 9389 10050 9394
rect 9758 9199 9759 9225
rect 9785 9199 9786 9225
rect 9758 9193 9786 9199
rect 10094 9226 10122 9231
rect 10122 9198 10178 9226
rect 10094 9179 10122 9198
rect 9646 9170 9674 9175
rect 9590 9169 9674 9170
rect 9590 9143 9647 9169
rect 9673 9143 9674 9169
rect 9590 9142 9674 9143
rect 9590 9058 9618 9142
rect 9646 9137 9674 9142
rect 9590 9025 9618 9030
rect 9758 9114 9786 9119
rect 9534 8857 9562 8862
rect 9758 8833 9786 9086
rect 9758 8807 9759 8833
rect 9785 8807 9786 8833
rect 9758 8801 9786 8807
rect 10150 8834 10178 9198
rect 10206 9225 10234 9231
rect 10206 9199 10207 9225
rect 10233 9199 10234 9225
rect 10206 9058 10234 9199
rect 10318 9225 10346 9702
rect 10374 9506 10402 9511
rect 10654 9506 10682 11158
rect 10710 9953 10738 11774
rect 10766 11689 10794 12278
rect 10934 12273 10962 12278
rect 10822 12138 10850 12143
rect 10822 11913 10850 12110
rect 10990 12026 11018 12031
rect 10990 11969 11018 11998
rect 10990 11943 10991 11969
rect 11017 11943 11018 11969
rect 10990 11937 11018 11943
rect 10822 11887 10823 11913
rect 10849 11887 10850 11913
rect 10822 11858 10850 11887
rect 11102 11913 11130 11919
rect 11102 11887 11103 11913
rect 11129 11887 11130 11913
rect 10822 11825 10850 11830
rect 11046 11857 11074 11863
rect 11046 11831 11047 11857
rect 11073 11831 11074 11857
rect 11046 11802 11074 11831
rect 11102 11858 11130 11887
rect 11158 11914 11186 12670
rect 11158 11881 11186 11886
rect 11270 12361 11298 12726
rect 11270 12335 11271 12361
rect 11297 12335 11298 12361
rect 11270 12026 11298 12335
rect 11382 12362 11410 13455
rect 11438 13482 11466 13487
rect 11662 13482 11690 13487
rect 11438 13481 11690 13482
rect 11438 13455 11439 13481
rect 11465 13455 11663 13481
rect 11689 13455 11690 13481
rect 11438 13454 11690 13455
rect 11438 13449 11466 13454
rect 11662 13449 11690 13454
rect 11774 13481 11802 13846
rect 12222 13841 12250 13846
rect 11830 13538 11858 13543
rect 11830 13491 11858 13510
rect 11774 13455 11775 13481
rect 11801 13455 11802 13481
rect 11774 13449 11802 13455
rect 12166 13258 12194 13263
rect 11774 12810 11802 12815
rect 11774 12473 11802 12782
rect 12166 12810 12194 13230
rect 12614 13258 12642 18607
rect 20118 18522 20146 18663
rect 20118 18489 20146 18494
rect 17598 18438 17730 18443
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17598 18405 17730 18410
rect 17598 17654 17730 17659
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17598 17621 17730 17626
rect 17598 16870 17730 16875
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17598 16837 17730 16842
rect 17598 16086 17730 16091
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17598 16053 17730 16058
rect 17598 15302 17730 15307
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17598 15269 17730 15274
rect 17598 14518 17730 14523
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17598 14485 17730 14490
rect 18942 13929 18970 13935
rect 18942 13903 18943 13929
rect 18969 13903 18970 13929
rect 12614 13225 12642 13230
rect 12726 13873 12754 13879
rect 12726 13847 12727 13873
rect 12753 13847 12754 13873
rect 12614 13146 12642 13151
rect 12726 13146 12754 13847
rect 17598 13734 17730 13739
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17598 13701 17730 13706
rect 13230 13538 13258 13543
rect 13174 13482 13202 13487
rect 13174 13435 13202 13454
rect 13230 13482 13258 13510
rect 13790 13537 13818 13543
rect 13790 13511 13791 13537
rect 13817 13511 13818 13537
rect 13790 13482 13818 13511
rect 18830 13537 18858 13543
rect 18830 13511 18831 13537
rect 18857 13511 18858 13537
rect 13230 13481 13482 13482
rect 13230 13455 13231 13481
rect 13257 13455 13482 13481
rect 13230 13454 13482 13455
rect 13230 13449 13258 13454
rect 12166 12763 12194 12782
rect 12558 13145 12754 13146
rect 12558 13119 12615 13145
rect 12641 13119 12754 13145
rect 12558 13118 12754 13119
rect 13062 13425 13090 13431
rect 13062 13399 13063 13425
rect 13089 13399 13090 13425
rect 12558 12753 12586 13118
rect 12614 13113 12642 13118
rect 13006 13090 13034 13095
rect 12558 12727 12559 12753
rect 12585 12727 12586 12753
rect 12390 12642 12418 12647
rect 12558 12642 12586 12727
rect 12418 12614 12586 12642
rect 12782 13089 13034 13090
rect 12782 13063 13007 13089
rect 13033 13063 13034 13089
rect 12782 13062 13034 13063
rect 12390 12595 12418 12614
rect 11774 12447 11775 12473
rect 11801 12447 11802 12473
rect 11774 12441 11802 12447
rect 12782 12473 12810 13062
rect 13006 13057 13034 13062
rect 13062 12922 13090 13399
rect 12894 12894 13090 12922
rect 12894 12586 12922 12894
rect 12950 12698 12978 12703
rect 12950 12697 13146 12698
rect 12950 12671 12951 12697
rect 12977 12671 13146 12697
rect 12950 12670 13146 12671
rect 12950 12665 12978 12670
rect 12894 12558 12978 12586
rect 12782 12447 12783 12473
rect 12809 12447 12810 12473
rect 12782 12441 12810 12447
rect 12894 12418 12922 12423
rect 12894 12371 12922 12390
rect 12950 12417 12978 12558
rect 12950 12391 12951 12417
rect 12977 12391 12978 12417
rect 12950 12385 12978 12391
rect 11494 12362 11522 12367
rect 11382 12361 11522 12362
rect 11382 12335 11495 12361
rect 11521 12335 11522 12361
rect 11382 12334 11522 12335
rect 11494 12138 11522 12334
rect 11662 12362 11690 12367
rect 11662 12315 11690 12334
rect 11774 12362 11802 12367
rect 11718 12305 11746 12311
rect 11718 12279 11719 12305
rect 11745 12279 11746 12305
rect 11718 12138 11746 12279
rect 11494 12105 11522 12110
rect 11662 12110 11746 12138
rect 11102 11825 11130 11830
rect 10934 11774 11074 11802
rect 11270 11774 11298 11998
rect 11662 11970 11690 12110
rect 11718 12026 11746 12031
rect 11718 11979 11746 11998
rect 11494 11942 11690 11970
rect 11438 11914 11466 11919
rect 11438 11867 11466 11886
rect 11494 11913 11522 11942
rect 11494 11887 11495 11913
rect 11521 11887 11522 11913
rect 11494 11881 11522 11887
rect 11382 11857 11410 11863
rect 11382 11831 11383 11857
rect 11409 11831 11410 11857
rect 10934 11746 10962 11774
rect 11270 11746 11354 11774
rect 10766 11663 10767 11689
rect 10793 11663 10794 11689
rect 10766 11657 10794 11663
rect 10822 11718 10962 11746
rect 10822 11633 10850 11718
rect 11326 11690 11354 11746
rect 10822 11607 10823 11633
rect 10849 11607 10850 11633
rect 10822 11601 10850 11607
rect 10990 11662 11354 11690
rect 10990 10794 11018 11662
rect 11158 11186 11186 11191
rect 11382 11186 11410 11831
rect 11606 11858 11634 11863
rect 11438 11186 11466 11191
rect 11158 11185 11298 11186
rect 11158 11159 11159 11185
rect 11185 11159 11298 11185
rect 11158 11158 11298 11159
rect 11382 11158 11438 11186
rect 11158 11153 11186 11158
rect 11214 11073 11242 11079
rect 11214 11047 11215 11073
rect 11241 11047 11242 11073
rect 10878 10766 11018 10794
rect 11046 10906 11074 10911
rect 10822 10738 10850 10743
rect 10822 10401 10850 10710
rect 10822 10375 10823 10401
rect 10849 10375 10850 10401
rect 10822 10369 10850 10375
rect 10710 9927 10711 9953
rect 10737 9927 10738 9953
rect 10710 9921 10738 9927
rect 10878 9617 10906 10766
rect 11046 9954 11074 10878
rect 11214 10122 11242 11047
rect 11046 9921 11074 9926
rect 11158 10094 11242 10122
rect 11158 9674 11186 10094
rect 11270 10065 11298 11158
rect 11438 11139 11466 11158
rect 11270 10039 11271 10065
rect 11297 10039 11298 10065
rect 11270 10033 11298 10039
rect 11326 11129 11354 11135
rect 11326 11103 11327 11129
rect 11353 11103 11354 11129
rect 11214 10009 11242 10015
rect 11214 9983 11215 10009
rect 11241 9983 11242 10009
rect 11214 9954 11242 9983
rect 11214 9921 11242 9926
rect 11214 9674 11242 9679
rect 11158 9673 11242 9674
rect 11158 9647 11215 9673
rect 11241 9647 11242 9673
rect 11158 9646 11242 9647
rect 11214 9641 11242 9646
rect 10878 9591 10879 9617
rect 10905 9591 10906 9617
rect 10374 9505 10850 9506
rect 10374 9479 10375 9505
rect 10401 9479 10850 9505
rect 10374 9478 10850 9479
rect 10374 9473 10402 9478
rect 10318 9199 10319 9225
rect 10345 9199 10346 9225
rect 10318 9193 10346 9199
rect 10486 9394 10514 9399
rect 10206 9025 10234 9030
rect 10430 9170 10458 9175
rect 10430 9002 10458 9142
rect 10262 8974 10458 9002
rect 10206 8834 10234 8839
rect 10150 8833 10234 8834
rect 10150 8807 10207 8833
rect 10233 8807 10234 8833
rect 10150 8806 10234 8807
rect 10206 8801 10234 8806
rect 10262 8777 10290 8974
rect 10374 8834 10402 8839
rect 10486 8834 10514 9366
rect 10598 9338 10626 9343
rect 10598 9337 10738 9338
rect 10598 9311 10599 9337
rect 10625 9311 10738 9337
rect 10598 9310 10738 9311
rect 10598 9305 10626 9310
rect 10710 9281 10738 9310
rect 10822 9337 10850 9478
rect 10822 9311 10823 9337
rect 10849 9311 10850 9337
rect 10822 9305 10850 9311
rect 10710 9255 10711 9281
rect 10737 9255 10738 9281
rect 10710 9249 10738 9255
rect 10878 9282 10906 9591
rect 11270 9562 11298 9567
rect 11326 9562 11354 11103
rect 11382 10009 11410 10015
rect 11382 9983 11383 10009
rect 11409 9983 11410 10009
rect 11382 9674 11410 9983
rect 11494 10010 11522 10015
rect 11494 9963 11522 9982
rect 11382 9641 11410 9646
rect 11298 9534 11354 9562
rect 11270 9529 11298 9534
rect 11606 9282 11634 11830
rect 11774 11802 11802 12334
rect 11886 12361 11914 12367
rect 11886 12335 11887 12361
rect 11913 12335 11914 12361
rect 11886 11970 11914 12335
rect 11886 11937 11914 11942
rect 12390 12362 12418 12367
rect 11774 11769 11802 11774
rect 12054 11802 12082 11807
rect 12054 11185 12082 11774
rect 12390 11297 12418 12334
rect 13118 12250 13146 12670
rect 13230 12474 13258 12479
rect 13230 12427 13258 12446
rect 13454 12417 13482 13454
rect 13790 13146 13818 13454
rect 13902 13482 13930 13487
rect 13902 13435 13930 13454
rect 18830 13258 18858 13511
rect 18942 13482 18970 13903
rect 18942 13449 18970 13454
rect 19950 13873 19978 13879
rect 19950 13847 19951 13873
rect 19977 13847 19978 13873
rect 19950 13482 19978 13847
rect 19950 13449 19978 13454
rect 20006 13593 20034 13599
rect 20006 13567 20007 13593
rect 20033 13567 20034 13593
rect 18830 13225 18858 13230
rect 14406 13202 14434 13207
rect 14406 13155 14434 13174
rect 13790 13113 13818 13118
rect 14070 13146 14098 13151
rect 14070 13089 14098 13118
rect 14294 13146 14322 13151
rect 14294 13099 14322 13118
rect 18830 13146 18858 13151
rect 18830 13099 18858 13118
rect 20006 13146 20034 13567
rect 20006 13113 20034 13118
rect 14070 13063 14071 13089
rect 14097 13063 14098 13089
rect 14070 13057 14098 13063
rect 14630 13089 14658 13095
rect 14630 13063 14631 13089
rect 14657 13063 14658 13089
rect 14014 12809 14042 12815
rect 14014 12783 14015 12809
rect 14041 12783 14042 12809
rect 13510 12754 13538 12759
rect 13510 12473 13538 12726
rect 14014 12754 14042 12783
rect 14014 12721 14042 12726
rect 14238 12642 14266 12647
rect 14238 12595 14266 12614
rect 14630 12642 14658 13063
rect 19950 13089 19978 13095
rect 19950 13063 19951 13089
rect 19977 13063 19978 13089
rect 17598 12950 17730 12955
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17598 12917 17730 12922
rect 19950 12810 19978 13063
rect 19950 12777 19978 12782
rect 20006 12809 20034 12815
rect 20006 12783 20007 12809
rect 20033 12783 20034 12809
rect 18830 12754 18858 12759
rect 18830 12707 18858 12726
rect 14630 12609 14658 12614
rect 13510 12447 13511 12473
rect 13537 12447 13538 12473
rect 13510 12441 13538 12447
rect 13622 12474 13650 12479
rect 13622 12427 13650 12446
rect 20006 12474 20034 12783
rect 20006 12441 20034 12446
rect 13454 12391 13455 12417
rect 13481 12391 13482 12417
rect 13454 12385 13482 12391
rect 13174 12362 13202 12367
rect 13174 12315 13202 12334
rect 13230 12250 13258 12255
rect 13118 12249 13258 12250
rect 13118 12223 13231 12249
rect 13257 12223 13258 12249
rect 13118 12222 13258 12223
rect 13230 12217 13258 12222
rect 17598 12166 17730 12171
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17598 12133 17730 12138
rect 13342 11970 13370 11975
rect 12390 11271 12391 11297
rect 12417 11271 12418 11297
rect 12390 11265 12418 11271
rect 12782 11298 12810 11303
rect 13342 11298 13370 11942
rect 17598 11382 17730 11387
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17598 11349 17730 11354
rect 13566 11298 13594 11303
rect 12782 11297 12866 11298
rect 12782 11271 12783 11297
rect 12809 11271 12866 11297
rect 12782 11270 12866 11271
rect 12782 11265 12810 11270
rect 12838 11242 12866 11270
rect 13342 11297 13594 11298
rect 13342 11271 13567 11297
rect 13593 11271 13594 11297
rect 13342 11270 13594 11271
rect 13286 11242 13314 11247
rect 12838 11241 13314 11242
rect 12838 11215 13287 11241
rect 13313 11215 13314 11241
rect 12838 11214 13314 11215
rect 13286 11209 13314 11214
rect 12054 11159 12055 11185
rect 12081 11159 12082 11185
rect 12054 11153 12082 11159
rect 12222 11186 12250 11191
rect 12222 11139 12250 11158
rect 12670 11186 12698 11191
rect 12782 11186 12810 11191
rect 12698 11158 12754 11186
rect 12670 11139 12698 11158
rect 12502 11129 12530 11135
rect 12502 11103 12503 11129
rect 12529 11103 12530 11129
rect 12334 11073 12362 11079
rect 12334 11047 12335 11073
rect 12361 11047 12362 11073
rect 11830 10066 11858 10071
rect 11830 10019 11858 10038
rect 11662 10009 11690 10015
rect 11662 9983 11663 10009
rect 11689 9983 11690 10009
rect 11662 9618 11690 9983
rect 11662 9585 11690 9590
rect 12166 10010 12194 10015
rect 10878 9254 10962 9282
rect 10374 8833 10514 8834
rect 10374 8807 10375 8833
rect 10401 8807 10514 8833
rect 10374 8806 10514 8807
rect 10542 9225 10570 9231
rect 10542 9199 10543 9225
rect 10569 9199 10570 9225
rect 10374 8801 10402 8806
rect 10262 8751 10263 8777
rect 10289 8751 10290 8777
rect 10262 8745 10290 8751
rect 9142 8610 9170 8694
rect 9366 8721 9394 8727
rect 9366 8695 9367 8721
rect 9393 8695 9394 8721
rect 9142 8582 9282 8610
rect 8694 8554 8722 8559
rect 8694 8507 8722 8526
rect 8862 8442 8890 8447
rect 8862 7938 8890 8414
rect 9254 8050 9282 8582
rect 9366 8442 9394 8695
rect 9926 8722 9954 8741
rect 9926 8689 9954 8694
rect 9918 8638 10050 8643
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 9918 8605 10050 8610
rect 9366 8409 9394 8414
rect 9982 8386 10010 8391
rect 9982 8339 10010 8358
rect 10542 8386 10570 9199
rect 10878 9114 10906 9119
rect 10878 9067 10906 9086
rect 10934 8442 10962 9254
rect 11606 9249 11634 9254
rect 12054 9282 12082 9287
rect 11046 9114 11074 9119
rect 11046 8497 11074 9086
rect 12054 8834 12082 9254
rect 11998 8833 12082 8834
rect 11998 8807 12055 8833
rect 12081 8807 12082 8833
rect 11998 8806 12082 8807
rect 11046 8471 11047 8497
rect 11073 8471 11074 8497
rect 11046 8465 11074 8471
rect 11102 8722 11130 8727
rect 10990 8442 11018 8447
rect 10934 8414 10990 8442
rect 10990 8409 11018 8414
rect 10038 8162 10066 8167
rect 10038 8161 10290 8162
rect 10038 8135 10039 8161
rect 10065 8135 10290 8161
rect 10038 8134 10290 8135
rect 10038 8129 10066 8134
rect 9254 8017 9282 8022
rect 10038 8050 10066 8055
rect 9030 7938 9058 7943
rect 8862 7910 9030 7938
rect 8750 7658 8778 7663
rect 8750 7611 8778 7630
rect 8414 7575 8415 7601
rect 8441 7575 8442 7601
rect 8414 7322 8442 7575
rect 9030 7602 9058 7910
rect 10038 7938 10066 8022
rect 10094 8050 10122 8055
rect 10094 8049 10178 8050
rect 10094 8023 10095 8049
rect 10121 8023 10178 8049
rect 10094 8022 10178 8023
rect 10094 8017 10122 8022
rect 10038 7937 10122 7938
rect 10038 7911 10039 7937
rect 10065 7911 10122 7937
rect 10038 7910 10122 7911
rect 10038 7905 10066 7910
rect 9918 7854 10050 7859
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 9918 7821 10050 7826
rect 10094 7713 10122 7910
rect 10150 7770 10178 8022
rect 10262 8049 10290 8134
rect 10262 8023 10263 8049
rect 10289 8023 10290 8049
rect 10262 8017 10290 8023
rect 10318 7937 10346 7943
rect 10430 7938 10458 7943
rect 10318 7911 10319 7937
rect 10345 7911 10346 7937
rect 10318 7826 10346 7911
rect 10318 7793 10346 7798
rect 10374 7937 10458 7938
rect 10374 7911 10431 7937
rect 10457 7911 10458 7937
rect 10374 7910 10458 7911
rect 10150 7737 10178 7742
rect 10094 7687 10095 7713
rect 10121 7687 10122 7713
rect 10094 7681 10122 7687
rect 9030 7569 9058 7574
rect 9814 7658 9842 7663
rect 8470 7322 8498 7327
rect 8414 7321 8498 7322
rect 8414 7295 8471 7321
rect 8497 7295 8498 7321
rect 8414 7294 8498 7295
rect 8470 7289 8498 7294
rect 8358 7239 8359 7265
rect 8385 7239 8386 7265
rect 8358 7233 8386 7239
rect 9814 6874 9842 7630
rect 10374 7378 10402 7910
rect 10430 7905 10458 7910
rect 10430 7658 10458 7677
rect 10430 7625 10458 7630
rect 10542 7574 10570 8358
rect 10878 7994 10906 7999
rect 10878 7947 10906 7966
rect 10710 7938 10738 7943
rect 10710 7891 10738 7910
rect 10598 7826 10626 7831
rect 10626 7798 10794 7826
rect 10598 7793 10626 7798
rect 10710 7658 10738 7663
rect 10710 7611 10738 7630
rect 10206 7350 10402 7378
rect 10430 7546 10570 7574
rect 9918 7070 10050 7075
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 9918 7037 10050 7042
rect 10206 6929 10234 7350
rect 10206 6903 10207 6929
rect 10233 6903 10234 6929
rect 10206 6897 10234 6903
rect 9870 6874 9898 6879
rect 9814 6873 9898 6874
rect 9814 6847 9871 6873
rect 9897 6847 9898 6873
rect 9814 6846 9898 6847
rect 9870 6841 9898 6846
rect 2238 6678 2370 6683
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2238 6645 2370 6650
rect 9918 6286 10050 6291
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 9918 6253 10050 6258
rect 2238 5894 2370 5899
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2238 5861 2370 5866
rect 9918 5502 10050 5507
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 9918 5469 10050 5474
rect 2238 5110 2370 5115
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2238 5077 2370 5082
rect 9918 4718 10050 4723
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 9918 4685 10050 4690
rect 2238 4326 2370 4331
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2238 4293 2370 4298
rect 10430 4214 10458 7546
rect 10766 7265 10794 7798
rect 11102 7574 11130 8694
rect 11438 8442 11466 8447
rect 11438 8386 11466 8414
rect 11662 8386 11690 8391
rect 11438 8385 11690 8386
rect 11438 8359 11663 8385
rect 11689 8359 11690 8385
rect 11438 8358 11690 8359
rect 11662 8050 11690 8358
rect 11718 8050 11746 8055
rect 11662 8049 11746 8050
rect 11662 8023 11719 8049
rect 11745 8023 11746 8049
rect 11662 8022 11746 8023
rect 10766 7239 10767 7265
rect 10793 7239 10794 7265
rect 10766 7233 10794 7239
rect 10934 7546 11130 7574
rect 11718 7658 11746 8022
rect 11998 7994 12026 8806
rect 12054 8801 12082 8806
rect 12166 8833 12194 9982
rect 12278 9674 12306 9679
rect 12278 9627 12306 9646
rect 12334 8946 12362 11047
rect 12502 9842 12530 11103
rect 12670 10793 12698 10799
rect 12670 10767 12671 10793
rect 12697 10767 12698 10793
rect 12670 10122 12698 10767
rect 12670 10009 12698 10094
rect 12670 9983 12671 10009
rect 12697 9983 12698 10009
rect 12670 9977 12698 9983
rect 12502 9809 12530 9814
rect 12614 9562 12642 9567
rect 12614 9515 12642 9534
rect 12726 9561 12754 11158
rect 12782 11185 12866 11186
rect 12782 11159 12783 11185
rect 12809 11159 12866 11185
rect 12782 11158 12866 11159
rect 12782 11153 12810 11158
rect 12838 10066 12866 11158
rect 13230 11130 13258 11135
rect 13342 11130 13370 11270
rect 13566 11265 13594 11270
rect 20006 11241 20034 11247
rect 20006 11215 20007 11241
rect 20033 11215 20034 11241
rect 13398 11186 13426 11191
rect 13398 11139 13426 11158
rect 13734 11185 13762 11191
rect 13734 11159 13735 11185
rect 13761 11159 13762 11185
rect 13230 11129 13370 11130
rect 13230 11103 13231 11129
rect 13257 11103 13370 11129
rect 13230 11102 13370 11103
rect 13230 11097 13258 11102
rect 12894 11074 12922 11079
rect 12894 11073 13034 11074
rect 12894 11047 12895 11073
rect 12921 11047 13034 11073
rect 12894 11046 13034 11047
rect 12894 11041 12922 11046
rect 13006 10849 13034 11046
rect 13006 10823 13007 10849
rect 13033 10823 13034 10849
rect 13006 10817 13034 10823
rect 13622 11073 13650 11079
rect 13622 11047 13623 11073
rect 13649 11047 13650 11073
rect 12838 9618 12866 10038
rect 12894 10570 12922 10575
rect 12894 9729 12922 10542
rect 13622 10570 13650 11047
rect 13734 10794 13762 11159
rect 13734 10761 13762 10766
rect 14070 11186 14098 11191
rect 14070 10737 14098 11158
rect 18830 11186 18858 11191
rect 18830 11139 18858 11158
rect 14070 10711 14071 10737
rect 14097 10711 14098 10737
rect 14070 10705 14098 10711
rect 14126 10794 14154 10799
rect 13622 10537 13650 10542
rect 13230 10345 13258 10351
rect 13230 10319 13231 10345
rect 13257 10319 13258 10345
rect 13230 10122 13258 10319
rect 14126 10094 14154 10766
rect 18830 10794 18858 10799
rect 18830 10747 18858 10766
rect 20006 10794 20034 11215
rect 20006 10761 20034 10766
rect 12894 9703 12895 9729
rect 12921 9703 12922 9729
rect 12894 9697 12922 9703
rect 13006 9953 13034 9959
rect 13006 9927 13007 9953
rect 13033 9927 13034 9953
rect 12894 9618 12922 9623
rect 12838 9617 12922 9618
rect 12838 9591 12895 9617
rect 12921 9591 12922 9617
rect 12838 9590 12922 9591
rect 12726 9535 12727 9561
rect 12753 9535 12754 9561
rect 12726 9450 12754 9535
rect 12726 9417 12754 9422
rect 12726 9282 12754 9287
rect 12334 8913 12362 8918
rect 12614 9281 12754 9282
rect 12614 9255 12727 9281
rect 12753 9255 12754 9281
rect 12614 9254 12754 9255
rect 12614 8946 12642 9254
rect 12726 9249 12754 9254
rect 12838 9282 12866 9287
rect 12838 9235 12866 9254
rect 12782 9170 12810 9175
rect 12782 9169 12866 9170
rect 12782 9143 12783 9169
rect 12809 9143 12866 9169
rect 12782 9142 12866 9143
rect 12782 9137 12810 9142
rect 12614 8913 12642 8918
rect 12726 9114 12754 9119
rect 12166 8807 12167 8833
rect 12193 8807 12194 8833
rect 12166 8801 12194 8807
rect 12670 8833 12698 8839
rect 12670 8807 12671 8833
rect 12697 8807 12698 8833
rect 12334 8778 12362 8783
rect 12222 8721 12250 8727
rect 12222 8695 12223 8721
rect 12249 8695 12250 8721
rect 12222 8497 12250 8695
rect 12278 8722 12306 8727
rect 12278 8675 12306 8694
rect 12222 8471 12223 8497
rect 12249 8471 12250 8497
rect 12222 8465 12250 8471
rect 12334 8442 12362 8750
rect 12670 8778 12698 8807
rect 12670 8745 12698 8750
rect 12334 8409 12362 8414
rect 12166 8330 12194 8335
rect 12054 8329 12194 8330
rect 12054 8303 12167 8329
rect 12193 8303 12194 8329
rect 12054 8302 12194 8303
rect 12054 8105 12082 8302
rect 12166 8297 12194 8302
rect 12054 8079 12055 8105
rect 12081 8079 12082 8105
rect 12054 8073 12082 8079
rect 11998 7961 12026 7966
rect 12614 7994 12642 7999
rect 12614 7713 12642 7966
rect 12726 7770 12754 9086
rect 12838 9002 12866 9142
rect 12894 9114 12922 9590
rect 13006 9505 13034 9927
rect 13006 9479 13007 9505
rect 13033 9479 13034 9505
rect 13006 9473 13034 9479
rect 13230 9505 13258 10094
rect 14070 10066 14154 10094
rect 14294 10737 14322 10743
rect 14294 10711 14295 10737
rect 14321 10711 14322 10737
rect 14294 10066 14322 10711
rect 19950 10737 19978 10743
rect 19950 10711 19951 10737
rect 19977 10711 19978 10737
rect 17598 10598 17730 10603
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17598 10565 17730 10570
rect 19950 10458 19978 10711
rect 19950 10425 19978 10430
rect 20006 10457 20034 10463
rect 20006 10431 20007 10457
rect 20033 10431 20034 10457
rect 14070 9953 14098 10066
rect 14070 9927 14071 9953
rect 14097 9927 14098 9953
rect 14070 9921 14098 9927
rect 13230 9479 13231 9505
rect 13257 9479 13258 9505
rect 13062 9226 13090 9231
rect 13062 9225 13146 9226
rect 13062 9199 13063 9225
rect 13089 9199 13146 9225
rect 13062 9198 13146 9199
rect 13062 9193 13090 9198
rect 12894 9081 12922 9086
rect 12838 8974 13034 9002
rect 13006 8889 13034 8974
rect 13006 8863 13007 8889
rect 13033 8863 13034 8889
rect 13006 8857 13034 8863
rect 13062 8722 13090 8727
rect 13062 8554 13090 8694
rect 12726 7723 12754 7742
rect 12894 8442 12922 8447
rect 12614 7687 12615 7713
rect 12641 7687 12642 7713
rect 12614 7681 12642 7687
rect 10934 7265 10962 7546
rect 10934 7239 10935 7265
rect 10961 7239 10962 7265
rect 10934 7233 10962 7239
rect 11494 7434 11522 7439
rect 10878 7153 10906 7159
rect 10878 7127 10879 7153
rect 10905 7127 10906 7153
rect 10878 6818 10906 7127
rect 11494 6985 11522 7406
rect 11718 7434 11746 7630
rect 12782 7658 12810 7663
rect 12782 7611 12810 7630
rect 12838 7657 12866 7663
rect 12838 7631 12839 7657
rect 12865 7631 12866 7657
rect 12334 7602 12362 7607
rect 11718 7401 11746 7406
rect 11998 7434 12026 7439
rect 11998 7265 12026 7406
rect 12334 7321 12362 7574
rect 12334 7295 12335 7321
rect 12361 7295 12362 7321
rect 12334 7289 12362 7295
rect 12838 7322 12866 7631
rect 12894 7657 12922 8414
rect 13062 8106 13090 8526
rect 13118 8330 13146 9198
rect 13174 8946 13202 8951
rect 13174 8554 13202 8918
rect 13230 8778 13258 9479
rect 14070 8946 14098 8951
rect 14070 8889 14098 8918
rect 14070 8863 14071 8889
rect 14097 8863 14098 8889
rect 14070 8857 14098 8863
rect 14294 8889 14322 10038
rect 18830 10401 18858 10407
rect 18830 10375 18831 10401
rect 18857 10375 18858 10401
rect 17598 9814 17730 9819
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17598 9781 17730 9786
rect 18830 9674 18858 10375
rect 20006 10122 20034 10431
rect 20006 10089 20034 10094
rect 18830 9641 18858 9646
rect 17598 9030 17730 9035
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17598 8997 17730 9002
rect 14294 8863 14295 8889
rect 14321 8863 14322 8889
rect 14294 8857 14322 8863
rect 20006 8889 20034 8895
rect 20006 8863 20007 8889
rect 20033 8863 20034 8889
rect 18830 8834 18858 8839
rect 18830 8787 18858 8806
rect 13342 8778 13370 8783
rect 13230 8750 13342 8778
rect 13230 8554 13258 8559
rect 13174 8553 13258 8554
rect 13174 8527 13231 8553
rect 13257 8527 13258 8553
rect 13174 8526 13258 8527
rect 13230 8521 13258 8526
rect 13174 8442 13202 8447
rect 13174 8395 13202 8414
rect 13230 8330 13258 8335
rect 13118 8329 13258 8330
rect 13118 8303 13231 8329
rect 13257 8303 13258 8329
rect 13118 8302 13258 8303
rect 13230 8297 13258 8302
rect 13118 8106 13146 8111
rect 13062 8105 13146 8106
rect 13062 8079 13119 8105
rect 13145 8079 13146 8105
rect 13062 8078 13146 8079
rect 13118 8073 13146 8078
rect 13342 7937 13370 8750
rect 20006 8778 20034 8863
rect 20006 8745 20034 8750
rect 18830 8442 18858 8447
rect 18830 8395 18858 8414
rect 20006 8442 20034 8447
rect 20006 8385 20034 8414
rect 20006 8359 20007 8385
rect 20033 8359 20034 8385
rect 20006 8353 20034 8359
rect 17598 8246 17730 8251
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17598 8213 17730 8218
rect 13342 7911 13343 7937
rect 13369 7911 13370 7937
rect 12894 7631 12895 7657
rect 12921 7631 12922 7657
rect 12894 7625 12922 7631
rect 13174 7658 13202 7663
rect 13118 7602 13146 7621
rect 13174 7611 13202 7630
rect 13118 7569 13146 7574
rect 13342 7434 13370 7911
rect 17598 7462 17730 7467
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 13370 7406 13650 7434
rect 17598 7429 17730 7434
rect 13342 7387 13370 7406
rect 13398 7322 13426 7327
rect 12838 7321 13426 7322
rect 12838 7295 13399 7321
rect 13425 7295 13426 7321
rect 12838 7294 13426 7295
rect 11998 7239 11999 7265
rect 12025 7239 12026 7265
rect 11998 7233 12026 7239
rect 11494 6959 11495 6985
rect 11521 6959 11522 6985
rect 11494 6953 11522 6959
rect 10878 4214 10906 6790
rect 11270 6818 11298 6823
rect 11270 6771 11298 6790
rect 13398 6426 13426 7294
rect 13622 7321 13650 7406
rect 13622 7295 13623 7321
rect 13649 7295 13650 7321
rect 13622 7289 13650 7295
rect 17598 6678 17730 6683
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17598 6645 17730 6650
rect 13398 6398 13482 6426
rect 10430 4186 10514 4214
rect 9918 3934 10050 3939
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 9918 3901 10050 3906
rect 2238 3542 2370 3547
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2238 3509 2370 3514
rect 9918 3150 10050 3155
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 9918 3117 10050 3122
rect 2238 2758 2370 2763
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2238 2725 2370 2730
rect 9918 2366 10050 2371
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 9918 2333 10050 2338
rect 10486 2170 10514 4186
rect 10486 2137 10514 2142
rect 10710 4186 10906 4214
rect 13454 4214 13482 6398
rect 17598 5894 17730 5899
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17598 5861 17730 5866
rect 17598 5110 17730 5115
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17598 5077 17730 5082
rect 17598 4326 17730 4331
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17598 4293 17730 4298
rect 13454 4186 13706 4214
rect 2238 1974 2370 1979
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2238 1941 2370 1946
rect 10710 1777 10738 4186
rect 10878 2170 10906 2175
rect 10878 2123 10906 2142
rect 10710 1751 10711 1777
rect 10737 1751 10738 1777
rect 10710 1745 10738 1751
rect 10766 2058 10794 2063
rect 3822 1666 3850 1671
rect 3710 1665 3850 1666
rect 3710 1639 3823 1665
rect 3849 1639 3850 1665
rect 3710 1638 3850 1639
rect 3710 400 3738 1638
rect 3822 1633 3850 1638
rect 9918 1582 10050 1587
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 9918 1549 10050 1554
rect 10766 400 10794 2030
rect 11382 2058 11410 2063
rect 11382 2011 11410 2030
rect 12782 1833 12810 1839
rect 12782 1807 12783 1833
rect 12809 1807 12810 1833
rect 11214 1666 11242 1671
rect 11102 1665 11242 1666
rect 11102 1639 11215 1665
rect 11241 1639 11242 1665
rect 11102 1638 11242 1639
rect 11102 400 11130 1638
rect 11214 1633 11242 1638
rect 12782 400 12810 1807
rect 13678 1777 13706 4186
rect 17598 3542 17730 3547
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17598 3509 17730 3514
rect 17598 2758 17730 2763
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17598 2725 17730 2730
rect 17598 1974 17730 1979
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17598 1941 17730 1946
rect 13678 1751 13679 1777
rect 13705 1751 13706 1777
rect 13678 1745 13706 1751
rect 3696 0 3752 400
rect 10752 0 10808 400
rect 11088 0 11144 400
rect 12768 0 12824 400
<< via2 >>
rect 2238 19221 2266 19222
rect 2238 19195 2239 19221
rect 2239 19195 2265 19221
rect 2265 19195 2266 19221
rect 2238 19194 2266 19195
rect 2290 19221 2318 19222
rect 2290 19195 2291 19221
rect 2291 19195 2317 19221
rect 2317 19195 2318 19221
rect 2290 19194 2318 19195
rect 2342 19221 2370 19222
rect 2342 19195 2343 19221
rect 2343 19195 2369 19221
rect 2369 19195 2370 19221
rect 2342 19194 2370 19195
rect 8414 18718 8442 18746
rect 2238 18437 2266 18438
rect 2238 18411 2239 18437
rect 2239 18411 2265 18437
rect 2265 18411 2266 18437
rect 2238 18410 2266 18411
rect 2290 18437 2318 18438
rect 2290 18411 2291 18437
rect 2291 18411 2317 18437
rect 2317 18411 2318 18437
rect 2290 18410 2318 18411
rect 2342 18437 2370 18438
rect 2342 18411 2343 18437
rect 2343 18411 2369 18437
rect 2369 18411 2370 18437
rect 2342 18410 2370 18411
rect 2238 17653 2266 17654
rect 2238 17627 2239 17653
rect 2239 17627 2265 17653
rect 2265 17627 2266 17653
rect 2238 17626 2266 17627
rect 2290 17653 2318 17654
rect 2290 17627 2291 17653
rect 2291 17627 2317 17653
rect 2317 17627 2318 17653
rect 2290 17626 2318 17627
rect 2342 17653 2370 17654
rect 2342 17627 2343 17653
rect 2343 17627 2369 17653
rect 2369 17627 2370 17653
rect 2342 17626 2370 17627
rect 2238 16869 2266 16870
rect 2238 16843 2239 16869
rect 2239 16843 2265 16869
rect 2265 16843 2266 16869
rect 2238 16842 2266 16843
rect 2290 16869 2318 16870
rect 2290 16843 2291 16869
rect 2291 16843 2317 16869
rect 2317 16843 2318 16869
rect 2290 16842 2318 16843
rect 2342 16869 2370 16870
rect 2342 16843 2343 16869
rect 2343 16843 2369 16869
rect 2369 16843 2370 16869
rect 2342 16842 2370 16843
rect 2238 16085 2266 16086
rect 2238 16059 2239 16085
rect 2239 16059 2265 16085
rect 2265 16059 2266 16085
rect 2238 16058 2266 16059
rect 2290 16085 2318 16086
rect 2290 16059 2291 16085
rect 2291 16059 2317 16085
rect 2317 16059 2318 16085
rect 2290 16058 2318 16059
rect 2342 16085 2370 16086
rect 2342 16059 2343 16085
rect 2343 16059 2369 16085
rect 2369 16059 2370 16085
rect 2342 16058 2370 16059
rect 9422 18942 9450 18970
rect 10374 18969 10402 18970
rect 10374 18943 10375 18969
rect 10375 18943 10401 18969
rect 10401 18943 10402 18969
rect 10374 18942 10402 18943
rect 9918 18829 9946 18830
rect 9918 18803 9919 18829
rect 9919 18803 9945 18829
rect 9945 18803 9946 18829
rect 9918 18802 9946 18803
rect 9970 18829 9998 18830
rect 9970 18803 9971 18829
rect 9971 18803 9997 18829
rect 9997 18803 9998 18829
rect 9970 18802 9998 18803
rect 10022 18829 10050 18830
rect 10022 18803 10023 18829
rect 10023 18803 10049 18829
rect 10049 18803 10050 18829
rect 10022 18802 10050 18803
rect 9198 18745 9226 18746
rect 9198 18719 9199 18745
rect 9199 18719 9225 18745
rect 9225 18719 9226 18745
rect 9198 18718 9226 18719
rect 11774 19110 11802 19138
rect 10430 18718 10458 18746
rect 9918 18045 9946 18046
rect 9918 18019 9919 18045
rect 9919 18019 9945 18045
rect 9945 18019 9946 18045
rect 9918 18018 9946 18019
rect 9970 18045 9998 18046
rect 9970 18019 9971 18045
rect 9971 18019 9997 18045
rect 9997 18019 9998 18045
rect 9970 18018 9998 18019
rect 10022 18045 10050 18046
rect 10022 18019 10023 18045
rect 10023 18019 10049 18045
rect 10049 18019 10050 18045
rect 10022 18018 10050 18019
rect 9918 17261 9946 17262
rect 9918 17235 9919 17261
rect 9919 17235 9945 17261
rect 9945 17235 9946 17261
rect 9918 17234 9946 17235
rect 9970 17261 9998 17262
rect 9970 17235 9971 17261
rect 9971 17235 9997 17261
rect 9997 17235 9998 17261
rect 9970 17234 9998 17235
rect 10022 17261 10050 17262
rect 10022 17235 10023 17261
rect 10023 17235 10049 17261
rect 10049 17235 10050 17261
rect 10022 17234 10050 17235
rect 9918 16477 9946 16478
rect 9918 16451 9919 16477
rect 9919 16451 9945 16477
rect 9945 16451 9946 16477
rect 9918 16450 9946 16451
rect 9970 16477 9998 16478
rect 9970 16451 9971 16477
rect 9971 16451 9997 16477
rect 9997 16451 9998 16477
rect 9970 16450 9998 16451
rect 10022 16477 10050 16478
rect 10022 16451 10023 16477
rect 10023 16451 10049 16477
rect 10049 16451 10050 16477
rect 10022 16450 10050 16451
rect 11046 18745 11074 18746
rect 11046 18719 11047 18745
rect 11047 18719 11073 18745
rect 11073 18719 11074 18745
rect 11046 18718 11074 18719
rect 17598 19221 17626 19222
rect 17598 19195 17599 19221
rect 17599 19195 17625 19221
rect 17625 19195 17626 19221
rect 17598 19194 17626 19195
rect 17650 19221 17678 19222
rect 17650 19195 17651 19221
rect 17651 19195 17677 19221
rect 17677 19195 17678 19221
rect 17650 19194 17678 19195
rect 17702 19221 17730 19222
rect 17702 19195 17703 19221
rect 17703 19195 17729 19221
rect 17729 19195 17730 19221
rect 17702 19194 17730 19195
rect 12782 19137 12810 19138
rect 12782 19111 12783 19137
rect 12783 19111 12809 19137
rect 12809 19111 12810 19137
rect 12782 19110 12810 19111
rect 12110 18718 12138 18746
rect 13118 18745 13146 18746
rect 13118 18719 13119 18745
rect 13119 18719 13145 18745
rect 13145 18719 13146 18745
rect 13118 18718 13146 18719
rect 2238 15301 2266 15302
rect 2238 15275 2239 15301
rect 2239 15275 2265 15301
rect 2265 15275 2266 15301
rect 2238 15274 2266 15275
rect 2290 15301 2318 15302
rect 2290 15275 2291 15301
rect 2291 15275 2317 15301
rect 2317 15275 2318 15301
rect 2290 15274 2318 15275
rect 2342 15301 2370 15302
rect 2342 15275 2343 15301
rect 2343 15275 2369 15301
rect 2369 15275 2370 15301
rect 2342 15274 2370 15275
rect 2238 14517 2266 14518
rect 2238 14491 2239 14517
rect 2239 14491 2265 14517
rect 2265 14491 2266 14517
rect 2238 14490 2266 14491
rect 2290 14517 2318 14518
rect 2290 14491 2291 14517
rect 2291 14491 2317 14517
rect 2317 14491 2318 14517
rect 2290 14490 2318 14491
rect 2342 14517 2370 14518
rect 2342 14491 2343 14517
rect 2343 14491 2369 14517
rect 2369 14491 2370 14517
rect 2342 14490 2370 14491
rect 2086 13790 2114 13818
rect 966 12446 994 12474
rect 2238 13733 2266 13734
rect 2238 13707 2239 13733
rect 2239 13707 2265 13733
rect 2265 13707 2266 13733
rect 2238 13706 2266 13707
rect 2290 13733 2318 13734
rect 2290 13707 2291 13733
rect 2291 13707 2317 13733
rect 2317 13707 2318 13733
rect 2290 13706 2318 13707
rect 2342 13733 2370 13734
rect 2342 13707 2343 13733
rect 2343 13707 2369 13733
rect 2369 13707 2370 13733
rect 2342 13706 2370 13707
rect 6566 13454 6594 13482
rect 8246 13510 8274 13538
rect 7070 13454 7098 13482
rect 7462 13230 7490 13258
rect 8190 13257 8218 13258
rect 8190 13231 8191 13257
rect 8191 13231 8217 13257
rect 8217 13231 8218 13257
rect 8190 13230 8218 13231
rect 8134 13145 8162 13146
rect 8134 13119 8135 13145
rect 8135 13119 8161 13145
rect 8161 13119 8162 13145
rect 8134 13118 8162 13119
rect 2238 12949 2266 12950
rect 2238 12923 2239 12949
rect 2239 12923 2265 12949
rect 2265 12923 2266 12949
rect 2238 12922 2266 12923
rect 2290 12949 2318 12950
rect 2290 12923 2291 12949
rect 2291 12923 2317 12949
rect 2317 12923 2318 12949
rect 2290 12922 2318 12923
rect 2342 12949 2370 12950
rect 2342 12923 2343 12949
rect 2343 12923 2369 12949
rect 2369 12923 2370 12949
rect 2342 12922 2370 12923
rect 4998 12809 5026 12810
rect 4998 12783 4999 12809
rect 4999 12783 5025 12809
rect 5025 12783 5026 12809
rect 4998 12782 5026 12783
rect 5950 12782 5978 12810
rect 2142 12753 2170 12754
rect 2142 12727 2143 12753
rect 2143 12727 2169 12753
rect 2169 12727 2170 12753
rect 2142 12726 2170 12727
rect 2238 12165 2266 12166
rect 2238 12139 2239 12165
rect 2239 12139 2265 12165
rect 2265 12139 2266 12165
rect 2238 12138 2266 12139
rect 2290 12165 2318 12166
rect 2290 12139 2291 12165
rect 2291 12139 2317 12165
rect 2317 12139 2318 12165
rect 2290 12138 2318 12139
rect 2342 12165 2370 12166
rect 2342 12139 2343 12165
rect 2343 12139 2369 12165
rect 2369 12139 2370 12165
rect 2342 12138 2370 12139
rect 8750 13537 8778 13538
rect 8750 13511 8751 13537
rect 8751 13511 8777 13537
rect 8777 13511 8778 13537
rect 8750 13510 8778 13511
rect 8526 13398 8554 13426
rect 8302 13201 8330 13202
rect 8302 13175 8303 13201
rect 8303 13175 8329 13201
rect 8329 13175 8330 13201
rect 8302 13174 8330 13175
rect 8862 13454 8890 13482
rect 9086 13481 9114 13482
rect 9086 13455 9087 13481
rect 9087 13455 9113 13481
rect 9113 13455 9114 13481
rect 9086 13454 9114 13455
rect 9918 15693 9946 15694
rect 9918 15667 9919 15693
rect 9919 15667 9945 15693
rect 9945 15667 9946 15693
rect 9918 15666 9946 15667
rect 9970 15693 9998 15694
rect 9970 15667 9971 15693
rect 9971 15667 9997 15693
rect 9997 15667 9998 15693
rect 9970 15666 9998 15667
rect 10022 15693 10050 15694
rect 10022 15667 10023 15693
rect 10023 15667 10049 15693
rect 10049 15667 10050 15693
rect 10022 15666 10050 15667
rect 9918 14909 9946 14910
rect 9918 14883 9919 14909
rect 9919 14883 9945 14909
rect 9945 14883 9946 14909
rect 9918 14882 9946 14883
rect 9970 14909 9998 14910
rect 9970 14883 9971 14909
rect 9971 14883 9997 14909
rect 9997 14883 9998 14909
rect 9970 14882 9998 14883
rect 10022 14909 10050 14910
rect 10022 14883 10023 14909
rect 10023 14883 10049 14909
rect 10049 14883 10050 14909
rect 10022 14882 10050 14883
rect 9918 14125 9946 14126
rect 9918 14099 9919 14125
rect 9919 14099 9945 14125
rect 9945 14099 9946 14125
rect 9918 14098 9946 14099
rect 9970 14125 9998 14126
rect 9970 14099 9971 14125
rect 9971 14099 9997 14125
rect 9997 14099 9998 14125
rect 9970 14098 9998 14099
rect 10022 14125 10050 14126
rect 10022 14099 10023 14125
rect 10023 14099 10049 14125
rect 10049 14099 10050 14125
rect 10022 14098 10050 14099
rect 8750 13398 8778 13426
rect 6062 12697 6090 12698
rect 6062 12671 6063 12697
rect 6063 12671 6089 12697
rect 6089 12671 6090 12697
rect 6062 12670 6090 12671
rect 6454 12614 6482 12642
rect 6342 12305 6370 12306
rect 6342 12279 6343 12305
rect 6343 12279 6369 12305
rect 6369 12279 6370 12305
rect 6342 12278 6370 12279
rect 2238 11381 2266 11382
rect 2238 11355 2239 11381
rect 2239 11355 2265 11381
rect 2265 11355 2266 11381
rect 2238 11354 2266 11355
rect 2290 11381 2318 11382
rect 2290 11355 2291 11381
rect 2291 11355 2317 11381
rect 2317 11355 2318 11381
rect 2290 11354 2318 11355
rect 2342 11381 2370 11382
rect 2342 11355 2343 11381
rect 2343 11355 2369 11381
rect 2369 11355 2370 11381
rect 2342 11354 2370 11355
rect 6958 12697 6986 12698
rect 6958 12671 6959 12697
rect 6959 12671 6985 12697
rect 6985 12671 6986 12697
rect 6958 12670 6986 12671
rect 6790 12641 6818 12642
rect 6790 12615 6791 12641
rect 6791 12615 6817 12641
rect 6817 12615 6818 12641
rect 6790 12614 6818 12615
rect 6790 12278 6818 12306
rect 6902 11998 6930 12026
rect 7014 12390 7042 12418
rect 7686 12417 7714 12418
rect 7686 12391 7687 12417
rect 7687 12391 7713 12417
rect 7713 12391 7714 12417
rect 7686 12390 7714 12391
rect 7630 12334 7658 12362
rect 7070 12222 7098 12250
rect 7630 12249 7658 12250
rect 7630 12223 7631 12249
rect 7631 12223 7657 12249
rect 7657 12223 7658 12249
rect 7630 12222 7658 12223
rect 7406 11774 7434 11802
rect 6398 11129 6426 11130
rect 6398 11103 6399 11129
rect 6399 11103 6425 11129
rect 6425 11103 6426 11129
rect 6398 11102 6426 11103
rect 6454 10990 6482 11018
rect 2142 10793 2170 10794
rect 2142 10767 2143 10793
rect 2143 10767 2169 10793
rect 2169 10767 2170 10793
rect 2142 10766 2170 10767
rect 4830 10766 4858 10794
rect 2086 10710 2114 10738
rect 2238 10597 2266 10598
rect 2238 10571 2239 10597
rect 2239 10571 2265 10597
rect 2265 10571 2266 10597
rect 2238 10570 2266 10571
rect 2290 10597 2318 10598
rect 2290 10571 2291 10597
rect 2291 10571 2317 10597
rect 2317 10571 2318 10597
rect 2290 10570 2318 10571
rect 2342 10597 2370 10598
rect 2342 10571 2343 10597
rect 2343 10571 2369 10597
rect 2369 10571 2370 10597
rect 2342 10570 2370 10571
rect 966 10430 994 10458
rect 4830 10374 4858 10402
rect 5054 10094 5082 10122
rect 6118 10262 6146 10290
rect 2238 9813 2266 9814
rect 2238 9787 2239 9813
rect 2239 9787 2265 9813
rect 2265 9787 2266 9813
rect 2238 9786 2266 9787
rect 2290 9813 2318 9814
rect 2290 9787 2291 9813
rect 2291 9787 2317 9813
rect 2317 9787 2318 9813
rect 2290 9786 2318 9787
rect 2342 9813 2370 9814
rect 2342 9787 2343 9813
rect 2343 9787 2369 9813
rect 2369 9787 2370 9813
rect 2342 9786 2370 9787
rect 2142 9225 2170 9226
rect 2142 9199 2143 9225
rect 2143 9199 2169 9225
rect 2169 9199 2170 9225
rect 2142 9198 2170 9199
rect 4998 9198 5026 9226
rect 966 9113 994 9114
rect 966 9087 967 9113
rect 967 9087 993 9113
rect 993 9087 994 9113
rect 966 9086 994 9087
rect 2238 9029 2266 9030
rect 2238 9003 2239 9029
rect 2239 9003 2265 9029
rect 2265 9003 2266 9029
rect 2238 9002 2266 9003
rect 2290 9029 2318 9030
rect 2290 9003 2291 9029
rect 2291 9003 2317 9029
rect 2317 9003 2318 9029
rect 2290 9002 2318 9003
rect 2342 9029 2370 9030
rect 2342 9003 2343 9029
rect 2343 9003 2369 9029
rect 2369 9003 2370 9029
rect 2342 9002 2370 9003
rect 966 8889 994 8890
rect 966 8863 967 8889
rect 967 8863 993 8889
rect 993 8863 994 8889
rect 966 8862 994 8863
rect 2142 8833 2170 8834
rect 2142 8807 2143 8833
rect 2143 8807 2169 8833
rect 2169 8807 2170 8833
rect 2142 8806 2170 8807
rect 6398 9814 6426 9842
rect 5894 8974 5922 9002
rect 6342 8806 6370 8834
rect 4998 8750 5026 8778
rect 966 8414 994 8442
rect 2142 8441 2170 8442
rect 2142 8415 2143 8441
rect 2143 8415 2169 8441
rect 2169 8415 2170 8441
rect 2142 8414 2170 8415
rect 2238 8245 2266 8246
rect 2238 8219 2239 8245
rect 2239 8219 2265 8245
rect 2265 8219 2266 8245
rect 2238 8218 2266 8219
rect 2290 8245 2318 8246
rect 2290 8219 2291 8245
rect 2291 8219 2317 8245
rect 2317 8219 2318 8245
rect 2290 8218 2318 8219
rect 2342 8245 2370 8246
rect 2342 8219 2343 8245
rect 2343 8219 2369 8245
rect 2369 8219 2370 8245
rect 2342 8218 2370 8219
rect 6286 8777 6314 8778
rect 6286 8751 6287 8777
rect 6287 8751 6313 8777
rect 6313 8751 6314 8777
rect 6286 8750 6314 8751
rect 5782 8694 5810 8722
rect 5782 8414 5810 8442
rect 6174 8638 6202 8666
rect 6622 10990 6650 11018
rect 6566 10934 6594 10962
rect 7294 11185 7322 11186
rect 7294 11159 7295 11185
rect 7295 11159 7321 11185
rect 7321 11159 7322 11185
rect 7294 11158 7322 11159
rect 6790 10878 6818 10906
rect 6622 10654 6650 10682
rect 6902 10598 6930 10626
rect 6790 10430 6818 10458
rect 6902 10401 6930 10402
rect 6902 10375 6903 10401
rect 6903 10375 6929 10401
rect 6929 10375 6930 10401
rect 6902 10374 6930 10375
rect 7126 11073 7154 11074
rect 7126 11047 7127 11073
rect 7127 11047 7153 11073
rect 7153 11047 7154 11073
rect 7126 11046 7154 11047
rect 7126 10934 7154 10962
rect 7518 11998 7546 12026
rect 7462 11606 7490 11634
rect 7854 11886 7882 11914
rect 7574 11633 7602 11634
rect 7574 11607 7575 11633
rect 7575 11607 7601 11633
rect 7601 11607 7602 11633
rect 7574 11606 7602 11607
rect 7462 11046 7490 11074
rect 7574 10990 7602 11018
rect 7686 11046 7714 11074
rect 7350 10457 7378 10458
rect 7350 10431 7351 10457
rect 7351 10431 7377 10457
rect 7377 10431 7378 10457
rect 7350 10430 7378 10431
rect 6846 10289 6874 10290
rect 6846 10263 6847 10289
rect 6847 10263 6873 10289
rect 6873 10263 6874 10289
rect 6846 10262 6874 10263
rect 6958 10121 6986 10122
rect 6958 10095 6959 10121
rect 6959 10095 6985 10121
rect 6985 10095 6986 10121
rect 6958 10094 6986 10095
rect 7294 10345 7322 10346
rect 7294 10319 7295 10345
rect 7295 10319 7321 10345
rect 7321 10319 7322 10345
rect 7294 10318 7322 10319
rect 7294 10094 7322 10122
rect 7630 10905 7658 10906
rect 7630 10879 7631 10905
rect 7631 10879 7657 10905
rect 7657 10879 7658 10905
rect 7630 10878 7658 10879
rect 7014 10038 7042 10066
rect 6566 9982 6594 10010
rect 7350 9702 7378 9730
rect 7462 9982 7490 10010
rect 7462 9646 7490 9674
rect 7126 9198 7154 9226
rect 6510 8750 6538 8778
rect 7014 9142 7042 9170
rect 7406 9198 7434 9226
rect 7742 10598 7770 10626
rect 7854 11102 7882 11130
rect 8134 11913 8162 11914
rect 8134 11887 8135 11913
rect 8135 11887 8161 11913
rect 8161 11887 8162 11913
rect 8134 11886 8162 11887
rect 7910 10990 7938 11018
rect 8470 11606 8498 11634
rect 8134 11158 8162 11186
rect 8190 10934 8218 10962
rect 7966 10766 7994 10794
rect 8078 10654 8106 10682
rect 7910 10345 7938 10346
rect 7910 10319 7911 10345
rect 7911 10319 7937 10345
rect 7937 10319 7938 10345
rect 7910 10318 7938 10319
rect 7630 9729 7658 9730
rect 7630 9703 7631 9729
rect 7631 9703 7657 9729
rect 7657 9703 7658 9729
rect 7630 9702 7658 9703
rect 7686 9534 7714 9562
rect 8302 10849 8330 10850
rect 8302 10823 8303 10849
rect 8303 10823 8329 10849
rect 8329 10823 8330 10849
rect 8302 10822 8330 10823
rect 8414 10766 8442 10794
rect 8358 10654 8386 10682
rect 8470 10542 8498 10570
rect 8190 10065 8218 10066
rect 8190 10039 8191 10065
rect 8191 10039 8217 10065
rect 8217 10039 8218 10065
rect 8190 10038 8218 10039
rect 8246 10430 8274 10458
rect 8022 9926 8050 9954
rect 7854 9617 7882 9618
rect 7854 9591 7855 9617
rect 7855 9591 7881 9617
rect 7881 9591 7882 9617
rect 7854 9590 7882 9591
rect 8022 9561 8050 9562
rect 8022 9535 8023 9561
rect 8023 9535 8049 9561
rect 8049 9535 8050 9561
rect 8022 9534 8050 9535
rect 7742 9478 7770 9506
rect 8414 10457 8442 10458
rect 8414 10431 8415 10457
rect 8415 10431 8441 10457
rect 8441 10431 8442 10457
rect 8414 10430 8442 10431
rect 8918 13145 8946 13146
rect 8918 13119 8919 13145
rect 8919 13119 8945 13145
rect 8945 13119 8946 13145
rect 8918 13118 8946 13119
rect 8918 12782 8946 12810
rect 8582 11438 8610 11466
rect 8582 10934 8610 10962
rect 8582 10318 8610 10346
rect 8302 10065 8330 10066
rect 8302 10039 8303 10065
rect 8303 10039 8329 10065
rect 8329 10039 8330 10065
rect 8302 10038 8330 10039
rect 9254 12809 9282 12810
rect 9254 12783 9255 12809
rect 9255 12783 9281 12809
rect 9281 12783 9282 12809
rect 9254 12782 9282 12783
rect 9422 13398 9450 13426
rect 10150 13537 10178 13538
rect 10150 13511 10151 13537
rect 10151 13511 10177 13537
rect 10177 13511 10178 13537
rect 10150 13510 10178 13511
rect 9918 13341 9946 13342
rect 9918 13315 9919 13341
rect 9919 13315 9945 13341
rect 9945 13315 9946 13341
rect 9918 13314 9946 13315
rect 9970 13341 9998 13342
rect 9970 13315 9971 13341
rect 9971 13315 9997 13341
rect 9997 13315 9998 13341
rect 9970 13314 9998 13315
rect 10022 13341 10050 13342
rect 10022 13315 10023 13341
rect 10023 13315 10049 13341
rect 10049 13315 10050 13341
rect 10022 13314 10050 13315
rect 9478 13174 9506 13202
rect 9030 12361 9058 12362
rect 9030 12335 9031 12361
rect 9031 12335 9057 12361
rect 9057 12335 9058 12361
rect 9030 12334 9058 12335
rect 8974 11718 9002 11746
rect 8806 11633 8834 11634
rect 8806 11607 8807 11633
rect 8807 11607 8833 11633
rect 8833 11607 8834 11633
rect 8806 11606 8834 11607
rect 9758 12334 9786 12362
rect 9702 11942 9730 11970
rect 8862 11465 8890 11466
rect 8862 11439 8863 11465
rect 8863 11439 8889 11465
rect 8889 11439 8890 11465
rect 8862 11438 8890 11439
rect 9030 10934 9058 10962
rect 8806 10710 8834 10738
rect 8750 10038 8778 10066
rect 8470 9982 8498 10010
rect 8302 9814 8330 9842
rect 8134 9478 8162 9506
rect 7686 9281 7714 9282
rect 7686 9255 7687 9281
rect 7687 9255 7713 9281
rect 7713 9255 7714 9281
rect 7686 9254 7714 9255
rect 7910 9337 7938 9338
rect 7910 9311 7911 9337
rect 7911 9311 7937 9337
rect 7937 9311 7938 9337
rect 7910 9310 7938 9311
rect 7742 9142 7770 9170
rect 7798 8918 7826 8946
rect 8022 8777 8050 8778
rect 8022 8751 8023 8777
rect 8023 8751 8049 8777
rect 8049 8751 8050 8777
rect 8022 8750 8050 8751
rect 7014 8638 7042 8666
rect 7518 8721 7546 8722
rect 7518 8695 7519 8721
rect 7519 8695 7545 8721
rect 7545 8695 7546 8721
rect 7518 8694 7546 8695
rect 8078 8721 8106 8722
rect 8078 8695 8079 8721
rect 8079 8695 8105 8721
rect 8105 8695 8106 8721
rect 8078 8694 8106 8695
rect 8022 8526 8050 8554
rect 6454 8049 6482 8050
rect 6454 8023 6455 8049
rect 6455 8023 6481 8049
rect 6481 8023 6482 8049
rect 6454 8022 6482 8023
rect 6790 8022 6818 8050
rect 7350 7966 7378 7994
rect 7014 7657 7042 7658
rect 7014 7631 7015 7657
rect 7015 7631 7041 7657
rect 7041 7631 7042 7657
rect 7014 7630 7042 7631
rect 8526 9673 8554 9674
rect 8526 9647 8527 9673
rect 8527 9647 8553 9673
rect 8553 9647 8554 9673
rect 8526 9646 8554 9647
rect 9086 10542 9114 10570
rect 9086 10401 9114 10402
rect 9086 10375 9087 10401
rect 9087 10375 9113 10401
rect 9113 10375 9114 10401
rect 9086 10374 9114 10375
rect 8974 10038 9002 10066
rect 8750 9561 8778 9562
rect 8750 9535 8751 9561
rect 8751 9535 8777 9561
rect 8777 9535 8778 9561
rect 8750 9534 8778 9535
rect 8694 9310 8722 9338
rect 9198 11438 9226 11466
rect 9198 10654 9226 10682
rect 9478 10822 9506 10850
rect 9310 10038 9338 10066
rect 9198 9982 9226 10010
rect 9478 10542 9506 10570
rect 9646 10430 9674 10458
rect 9918 12557 9946 12558
rect 9918 12531 9919 12557
rect 9919 12531 9945 12557
rect 9945 12531 9946 12557
rect 9918 12530 9946 12531
rect 9970 12557 9998 12558
rect 9970 12531 9971 12557
rect 9971 12531 9997 12557
rect 9997 12531 9998 12557
rect 9970 12530 9998 12531
rect 10022 12557 10050 12558
rect 10022 12531 10023 12557
rect 10023 12531 10049 12557
rect 10049 12531 10050 12557
rect 10022 12530 10050 12531
rect 9870 12305 9898 12306
rect 9870 12279 9871 12305
rect 9871 12279 9897 12305
rect 9897 12279 9898 12305
rect 9870 12278 9898 12279
rect 10766 12753 10794 12754
rect 10766 12727 10767 12753
rect 10767 12727 10793 12753
rect 10793 12727 10794 12753
rect 10766 12726 10794 12727
rect 11270 12726 11298 12754
rect 10654 12278 10682 12306
rect 10710 11969 10738 11970
rect 10710 11943 10711 11969
rect 10711 11943 10737 11969
rect 10737 11943 10738 11969
rect 10710 11942 10738 11943
rect 10542 11830 10570 11858
rect 9814 11718 9842 11746
rect 9918 11773 9946 11774
rect 9918 11747 9919 11773
rect 9919 11747 9945 11773
rect 9945 11747 9946 11773
rect 9918 11746 9946 11747
rect 9970 11773 9998 11774
rect 9970 11747 9971 11773
rect 9971 11747 9997 11773
rect 9997 11747 9998 11773
rect 9970 11746 9998 11747
rect 10022 11773 10050 11774
rect 10022 11747 10023 11773
rect 10023 11747 10049 11773
rect 10049 11747 10050 11773
rect 10022 11746 10050 11747
rect 10710 11774 10738 11802
rect 10542 11102 10570 11130
rect 10654 11158 10682 11186
rect 9918 10989 9946 10990
rect 9918 10963 9919 10989
rect 9919 10963 9945 10989
rect 9945 10963 9946 10989
rect 9918 10962 9946 10963
rect 9970 10989 9998 10990
rect 9970 10963 9971 10989
rect 9971 10963 9997 10989
rect 9997 10963 9998 10989
rect 9970 10962 9998 10963
rect 10022 10989 10050 10990
rect 10022 10963 10023 10989
rect 10023 10963 10049 10989
rect 10049 10963 10050 10989
rect 10022 10962 10050 10963
rect 9814 10878 9842 10906
rect 9758 10710 9786 10738
rect 9814 10598 9842 10626
rect 9814 10457 9842 10458
rect 9814 10431 9815 10457
rect 9815 10431 9841 10457
rect 9841 10431 9842 10457
rect 9814 10430 9842 10431
rect 9590 9982 9618 10010
rect 9422 9870 9450 9898
rect 9366 9590 9394 9618
rect 8414 9113 8442 9114
rect 8414 9087 8415 9113
rect 8415 9087 8441 9113
rect 8441 9087 8442 9113
rect 8414 9086 8442 9087
rect 9086 9086 9114 9114
rect 9030 8974 9058 9002
rect 9086 8889 9114 8890
rect 9086 8863 9087 8889
rect 9087 8863 9113 8889
rect 9113 8863 9114 8889
rect 9086 8862 9114 8863
rect 8302 8694 8330 8722
rect 8414 8777 8442 8778
rect 8414 8751 8415 8777
rect 8415 8751 8441 8777
rect 8441 8751 8442 8777
rect 8414 8750 8442 8751
rect 8134 7993 8162 7994
rect 8134 7967 8135 7993
rect 8135 7967 8161 7993
rect 8161 7967 8162 7993
rect 8134 7966 8162 7967
rect 7462 7630 7490 7658
rect 8358 7574 8386 7602
rect 2238 7461 2266 7462
rect 2238 7435 2239 7461
rect 2239 7435 2265 7461
rect 2265 7435 2266 7461
rect 2238 7434 2266 7435
rect 2290 7461 2318 7462
rect 2290 7435 2291 7461
rect 2291 7435 2317 7461
rect 2317 7435 2318 7461
rect 2290 7434 2318 7435
rect 2342 7461 2370 7462
rect 2342 7435 2343 7461
rect 2343 7435 2369 7461
rect 2369 7435 2370 7461
rect 2342 7434 2370 7435
rect 8750 8777 8778 8778
rect 8750 8751 8751 8777
rect 8751 8751 8777 8777
rect 8777 8751 8778 8777
rect 8750 8750 8778 8751
rect 9478 9142 9506 9170
rect 9918 10205 9946 10206
rect 9918 10179 9919 10205
rect 9919 10179 9945 10205
rect 9945 10179 9946 10205
rect 9918 10178 9946 10179
rect 9970 10205 9998 10206
rect 9970 10179 9971 10205
rect 9971 10179 9997 10205
rect 9997 10179 9998 10205
rect 9970 10178 9998 10179
rect 10022 10205 10050 10206
rect 10022 10179 10023 10205
rect 10023 10179 10049 10205
rect 10049 10179 10050 10205
rect 10022 10178 10050 10179
rect 10094 10038 10122 10066
rect 9758 9926 9786 9954
rect 10150 9870 10178 9898
rect 10318 9982 10346 10010
rect 9982 9729 10010 9730
rect 9982 9703 9983 9729
rect 9983 9703 10009 9729
rect 10009 9703 10010 9729
rect 9982 9702 10010 9703
rect 10318 9702 10346 9730
rect 9198 9030 9226 9058
rect 10206 9617 10234 9618
rect 10206 9591 10207 9617
rect 10207 9591 10233 9617
rect 10233 9591 10234 9617
rect 10206 9590 10234 9591
rect 9918 9421 9946 9422
rect 9918 9395 9919 9421
rect 9919 9395 9945 9421
rect 9945 9395 9946 9421
rect 9918 9394 9946 9395
rect 9970 9421 9998 9422
rect 9970 9395 9971 9421
rect 9971 9395 9997 9421
rect 9997 9395 9998 9421
rect 9970 9394 9998 9395
rect 10022 9421 10050 9422
rect 10022 9395 10023 9421
rect 10023 9395 10049 9421
rect 10049 9395 10050 9421
rect 10022 9394 10050 9395
rect 10094 9225 10122 9226
rect 10094 9199 10095 9225
rect 10095 9199 10121 9225
rect 10121 9199 10122 9225
rect 10094 9198 10122 9199
rect 9590 9030 9618 9058
rect 9758 9086 9786 9114
rect 9534 8862 9562 8890
rect 10822 12110 10850 12138
rect 10990 11998 11018 12026
rect 10822 11830 10850 11858
rect 11158 11886 11186 11914
rect 11830 13537 11858 13538
rect 11830 13511 11831 13537
rect 11831 13511 11857 13537
rect 11857 13511 11858 13537
rect 11830 13510 11858 13511
rect 12166 13230 12194 13258
rect 11774 12782 11802 12810
rect 20118 18494 20146 18522
rect 17598 18437 17626 18438
rect 17598 18411 17599 18437
rect 17599 18411 17625 18437
rect 17625 18411 17626 18437
rect 17598 18410 17626 18411
rect 17650 18437 17678 18438
rect 17650 18411 17651 18437
rect 17651 18411 17677 18437
rect 17677 18411 17678 18437
rect 17650 18410 17678 18411
rect 17702 18437 17730 18438
rect 17702 18411 17703 18437
rect 17703 18411 17729 18437
rect 17729 18411 17730 18437
rect 17702 18410 17730 18411
rect 17598 17653 17626 17654
rect 17598 17627 17599 17653
rect 17599 17627 17625 17653
rect 17625 17627 17626 17653
rect 17598 17626 17626 17627
rect 17650 17653 17678 17654
rect 17650 17627 17651 17653
rect 17651 17627 17677 17653
rect 17677 17627 17678 17653
rect 17650 17626 17678 17627
rect 17702 17653 17730 17654
rect 17702 17627 17703 17653
rect 17703 17627 17729 17653
rect 17729 17627 17730 17653
rect 17702 17626 17730 17627
rect 17598 16869 17626 16870
rect 17598 16843 17599 16869
rect 17599 16843 17625 16869
rect 17625 16843 17626 16869
rect 17598 16842 17626 16843
rect 17650 16869 17678 16870
rect 17650 16843 17651 16869
rect 17651 16843 17677 16869
rect 17677 16843 17678 16869
rect 17650 16842 17678 16843
rect 17702 16869 17730 16870
rect 17702 16843 17703 16869
rect 17703 16843 17729 16869
rect 17729 16843 17730 16869
rect 17702 16842 17730 16843
rect 17598 16085 17626 16086
rect 17598 16059 17599 16085
rect 17599 16059 17625 16085
rect 17625 16059 17626 16085
rect 17598 16058 17626 16059
rect 17650 16085 17678 16086
rect 17650 16059 17651 16085
rect 17651 16059 17677 16085
rect 17677 16059 17678 16085
rect 17650 16058 17678 16059
rect 17702 16085 17730 16086
rect 17702 16059 17703 16085
rect 17703 16059 17729 16085
rect 17729 16059 17730 16085
rect 17702 16058 17730 16059
rect 17598 15301 17626 15302
rect 17598 15275 17599 15301
rect 17599 15275 17625 15301
rect 17625 15275 17626 15301
rect 17598 15274 17626 15275
rect 17650 15301 17678 15302
rect 17650 15275 17651 15301
rect 17651 15275 17677 15301
rect 17677 15275 17678 15301
rect 17650 15274 17678 15275
rect 17702 15301 17730 15302
rect 17702 15275 17703 15301
rect 17703 15275 17729 15301
rect 17729 15275 17730 15301
rect 17702 15274 17730 15275
rect 17598 14517 17626 14518
rect 17598 14491 17599 14517
rect 17599 14491 17625 14517
rect 17625 14491 17626 14517
rect 17598 14490 17626 14491
rect 17650 14517 17678 14518
rect 17650 14491 17651 14517
rect 17651 14491 17677 14517
rect 17677 14491 17678 14517
rect 17650 14490 17678 14491
rect 17702 14517 17730 14518
rect 17702 14491 17703 14517
rect 17703 14491 17729 14517
rect 17729 14491 17730 14517
rect 17702 14490 17730 14491
rect 12614 13230 12642 13258
rect 17598 13733 17626 13734
rect 17598 13707 17599 13733
rect 17599 13707 17625 13733
rect 17625 13707 17626 13733
rect 17598 13706 17626 13707
rect 17650 13733 17678 13734
rect 17650 13707 17651 13733
rect 17651 13707 17677 13733
rect 17677 13707 17678 13733
rect 17650 13706 17678 13707
rect 17702 13733 17730 13734
rect 17702 13707 17703 13733
rect 17703 13707 17729 13733
rect 17729 13707 17730 13733
rect 17702 13706 17730 13707
rect 13230 13510 13258 13538
rect 13174 13481 13202 13482
rect 13174 13455 13175 13481
rect 13175 13455 13201 13481
rect 13201 13455 13202 13481
rect 13174 13454 13202 13455
rect 12166 12809 12194 12810
rect 12166 12783 12167 12809
rect 12167 12783 12193 12809
rect 12193 12783 12194 12809
rect 12166 12782 12194 12783
rect 12390 12641 12418 12642
rect 12390 12615 12391 12641
rect 12391 12615 12417 12641
rect 12417 12615 12418 12641
rect 12390 12614 12418 12615
rect 12894 12417 12922 12418
rect 12894 12391 12895 12417
rect 12895 12391 12921 12417
rect 12921 12391 12922 12417
rect 12894 12390 12922 12391
rect 11662 12361 11690 12362
rect 11662 12335 11663 12361
rect 11663 12335 11689 12361
rect 11689 12335 11690 12361
rect 11662 12334 11690 12335
rect 11774 12334 11802 12362
rect 11494 12110 11522 12138
rect 11270 11998 11298 12026
rect 11102 11830 11130 11858
rect 11718 12025 11746 12026
rect 11718 11999 11719 12025
rect 11719 11999 11745 12025
rect 11745 11999 11746 12025
rect 11718 11998 11746 11999
rect 11438 11913 11466 11914
rect 11438 11887 11439 11913
rect 11439 11887 11465 11913
rect 11465 11887 11466 11913
rect 11438 11886 11466 11887
rect 11606 11830 11634 11858
rect 11438 11185 11466 11186
rect 11438 11159 11439 11185
rect 11439 11159 11465 11185
rect 11465 11159 11466 11185
rect 11438 11158 11466 11159
rect 11046 10878 11074 10906
rect 10822 10737 10850 10738
rect 10822 10711 10823 10737
rect 10823 10711 10849 10737
rect 10849 10711 10850 10737
rect 10822 10710 10850 10711
rect 11046 9926 11074 9954
rect 11214 9926 11242 9954
rect 10486 9366 10514 9394
rect 10206 9030 10234 9058
rect 10430 9169 10458 9170
rect 10430 9143 10431 9169
rect 10431 9143 10457 9169
rect 10457 9143 10458 9169
rect 10430 9142 10458 9143
rect 11494 10009 11522 10010
rect 11494 9983 11495 10009
rect 11495 9983 11521 10009
rect 11521 9983 11522 10009
rect 11494 9982 11522 9983
rect 11382 9646 11410 9674
rect 11270 9534 11298 9562
rect 11886 11942 11914 11970
rect 12390 12334 12418 12362
rect 11774 11774 11802 11802
rect 12054 11774 12082 11802
rect 13230 12473 13258 12474
rect 13230 12447 13231 12473
rect 13231 12447 13257 12473
rect 13257 12447 13258 12473
rect 13230 12446 13258 12447
rect 13790 13454 13818 13482
rect 13902 13481 13930 13482
rect 13902 13455 13903 13481
rect 13903 13455 13929 13481
rect 13929 13455 13930 13481
rect 13902 13454 13930 13455
rect 18942 13454 18970 13482
rect 19950 13454 19978 13482
rect 18830 13230 18858 13258
rect 14406 13201 14434 13202
rect 14406 13175 14407 13201
rect 14407 13175 14433 13201
rect 14433 13175 14434 13201
rect 14406 13174 14434 13175
rect 13790 13118 13818 13146
rect 14070 13118 14098 13146
rect 14294 13145 14322 13146
rect 14294 13119 14295 13145
rect 14295 13119 14321 13145
rect 14321 13119 14322 13145
rect 14294 13118 14322 13119
rect 18830 13145 18858 13146
rect 18830 13119 18831 13145
rect 18831 13119 18857 13145
rect 18857 13119 18858 13145
rect 18830 13118 18858 13119
rect 20006 13118 20034 13146
rect 13510 12726 13538 12754
rect 14014 12726 14042 12754
rect 14238 12641 14266 12642
rect 14238 12615 14239 12641
rect 14239 12615 14265 12641
rect 14265 12615 14266 12641
rect 14238 12614 14266 12615
rect 17598 12949 17626 12950
rect 17598 12923 17599 12949
rect 17599 12923 17625 12949
rect 17625 12923 17626 12949
rect 17598 12922 17626 12923
rect 17650 12949 17678 12950
rect 17650 12923 17651 12949
rect 17651 12923 17677 12949
rect 17677 12923 17678 12949
rect 17650 12922 17678 12923
rect 17702 12949 17730 12950
rect 17702 12923 17703 12949
rect 17703 12923 17729 12949
rect 17729 12923 17730 12949
rect 17702 12922 17730 12923
rect 19950 12782 19978 12810
rect 18830 12753 18858 12754
rect 18830 12727 18831 12753
rect 18831 12727 18857 12753
rect 18857 12727 18858 12753
rect 18830 12726 18858 12727
rect 14630 12614 14658 12642
rect 13622 12473 13650 12474
rect 13622 12447 13623 12473
rect 13623 12447 13649 12473
rect 13649 12447 13650 12473
rect 13622 12446 13650 12447
rect 20006 12446 20034 12474
rect 13174 12361 13202 12362
rect 13174 12335 13175 12361
rect 13175 12335 13201 12361
rect 13201 12335 13202 12361
rect 13174 12334 13202 12335
rect 17598 12165 17626 12166
rect 17598 12139 17599 12165
rect 17599 12139 17625 12165
rect 17625 12139 17626 12165
rect 17598 12138 17626 12139
rect 17650 12165 17678 12166
rect 17650 12139 17651 12165
rect 17651 12139 17677 12165
rect 17677 12139 17678 12165
rect 17650 12138 17678 12139
rect 17702 12165 17730 12166
rect 17702 12139 17703 12165
rect 17703 12139 17729 12165
rect 17729 12139 17730 12165
rect 17702 12138 17730 12139
rect 13342 11942 13370 11970
rect 17598 11381 17626 11382
rect 17598 11355 17599 11381
rect 17599 11355 17625 11381
rect 17625 11355 17626 11381
rect 17598 11354 17626 11355
rect 17650 11381 17678 11382
rect 17650 11355 17651 11381
rect 17651 11355 17677 11381
rect 17677 11355 17678 11381
rect 17650 11354 17678 11355
rect 17702 11381 17730 11382
rect 17702 11355 17703 11381
rect 17703 11355 17729 11381
rect 17729 11355 17730 11381
rect 17702 11354 17730 11355
rect 12222 11185 12250 11186
rect 12222 11159 12223 11185
rect 12223 11159 12249 11185
rect 12249 11159 12250 11185
rect 12222 11158 12250 11159
rect 12670 11185 12698 11186
rect 12670 11159 12671 11185
rect 12671 11159 12697 11185
rect 12697 11159 12698 11185
rect 12670 11158 12698 11159
rect 11830 10065 11858 10066
rect 11830 10039 11831 10065
rect 11831 10039 11857 10065
rect 11857 10039 11858 10065
rect 11830 10038 11858 10039
rect 11662 9590 11690 9618
rect 12166 9982 12194 10010
rect 9142 8694 9170 8722
rect 8694 8553 8722 8554
rect 8694 8527 8695 8553
rect 8695 8527 8721 8553
rect 8721 8527 8722 8553
rect 8694 8526 8722 8527
rect 8862 8441 8890 8442
rect 8862 8415 8863 8441
rect 8863 8415 8889 8441
rect 8889 8415 8890 8441
rect 8862 8414 8890 8415
rect 9926 8721 9954 8722
rect 9926 8695 9927 8721
rect 9927 8695 9953 8721
rect 9953 8695 9954 8721
rect 9926 8694 9954 8695
rect 9918 8637 9946 8638
rect 9918 8611 9919 8637
rect 9919 8611 9945 8637
rect 9945 8611 9946 8637
rect 9918 8610 9946 8611
rect 9970 8637 9998 8638
rect 9970 8611 9971 8637
rect 9971 8611 9997 8637
rect 9997 8611 9998 8637
rect 9970 8610 9998 8611
rect 10022 8637 10050 8638
rect 10022 8611 10023 8637
rect 10023 8611 10049 8637
rect 10049 8611 10050 8637
rect 10022 8610 10050 8611
rect 9366 8414 9394 8442
rect 9982 8385 10010 8386
rect 9982 8359 9983 8385
rect 9983 8359 10009 8385
rect 10009 8359 10010 8385
rect 9982 8358 10010 8359
rect 10878 9113 10906 9114
rect 10878 9087 10879 9113
rect 10879 9087 10905 9113
rect 10905 9087 10906 9113
rect 10878 9086 10906 9087
rect 11606 9254 11634 9282
rect 12054 9254 12082 9282
rect 11046 9086 11074 9114
rect 11102 8694 11130 8722
rect 10990 8414 11018 8442
rect 10542 8358 10570 8386
rect 9254 8022 9282 8050
rect 10038 8022 10066 8050
rect 9030 7910 9058 7938
rect 8750 7657 8778 7658
rect 8750 7631 8751 7657
rect 8751 7631 8777 7657
rect 8777 7631 8778 7657
rect 8750 7630 8778 7631
rect 9918 7853 9946 7854
rect 9918 7827 9919 7853
rect 9919 7827 9945 7853
rect 9945 7827 9946 7853
rect 9918 7826 9946 7827
rect 9970 7853 9998 7854
rect 9970 7827 9971 7853
rect 9971 7827 9997 7853
rect 9997 7827 9998 7853
rect 9970 7826 9998 7827
rect 10022 7853 10050 7854
rect 10022 7827 10023 7853
rect 10023 7827 10049 7853
rect 10049 7827 10050 7853
rect 10022 7826 10050 7827
rect 10318 7798 10346 7826
rect 10150 7742 10178 7770
rect 9030 7601 9058 7602
rect 9030 7575 9031 7601
rect 9031 7575 9057 7601
rect 9057 7575 9058 7601
rect 9030 7574 9058 7575
rect 9814 7630 9842 7658
rect 10430 7657 10458 7658
rect 10430 7631 10431 7657
rect 10431 7631 10457 7657
rect 10457 7631 10458 7657
rect 10430 7630 10458 7631
rect 10878 7993 10906 7994
rect 10878 7967 10879 7993
rect 10879 7967 10905 7993
rect 10905 7967 10906 7993
rect 10878 7966 10906 7967
rect 10710 7937 10738 7938
rect 10710 7911 10711 7937
rect 10711 7911 10737 7937
rect 10737 7911 10738 7937
rect 10710 7910 10738 7911
rect 10598 7798 10626 7826
rect 10710 7657 10738 7658
rect 10710 7631 10711 7657
rect 10711 7631 10737 7657
rect 10737 7631 10738 7657
rect 10710 7630 10738 7631
rect 9918 7069 9946 7070
rect 9918 7043 9919 7069
rect 9919 7043 9945 7069
rect 9945 7043 9946 7069
rect 9918 7042 9946 7043
rect 9970 7069 9998 7070
rect 9970 7043 9971 7069
rect 9971 7043 9997 7069
rect 9997 7043 9998 7069
rect 9970 7042 9998 7043
rect 10022 7069 10050 7070
rect 10022 7043 10023 7069
rect 10023 7043 10049 7069
rect 10049 7043 10050 7069
rect 10022 7042 10050 7043
rect 2238 6677 2266 6678
rect 2238 6651 2239 6677
rect 2239 6651 2265 6677
rect 2265 6651 2266 6677
rect 2238 6650 2266 6651
rect 2290 6677 2318 6678
rect 2290 6651 2291 6677
rect 2291 6651 2317 6677
rect 2317 6651 2318 6677
rect 2290 6650 2318 6651
rect 2342 6677 2370 6678
rect 2342 6651 2343 6677
rect 2343 6651 2369 6677
rect 2369 6651 2370 6677
rect 2342 6650 2370 6651
rect 9918 6285 9946 6286
rect 9918 6259 9919 6285
rect 9919 6259 9945 6285
rect 9945 6259 9946 6285
rect 9918 6258 9946 6259
rect 9970 6285 9998 6286
rect 9970 6259 9971 6285
rect 9971 6259 9997 6285
rect 9997 6259 9998 6285
rect 9970 6258 9998 6259
rect 10022 6285 10050 6286
rect 10022 6259 10023 6285
rect 10023 6259 10049 6285
rect 10049 6259 10050 6285
rect 10022 6258 10050 6259
rect 2238 5893 2266 5894
rect 2238 5867 2239 5893
rect 2239 5867 2265 5893
rect 2265 5867 2266 5893
rect 2238 5866 2266 5867
rect 2290 5893 2318 5894
rect 2290 5867 2291 5893
rect 2291 5867 2317 5893
rect 2317 5867 2318 5893
rect 2290 5866 2318 5867
rect 2342 5893 2370 5894
rect 2342 5867 2343 5893
rect 2343 5867 2369 5893
rect 2369 5867 2370 5893
rect 2342 5866 2370 5867
rect 9918 5501 9946 5502
rect 9918 5475 9919 5501
rect 9919 5475 9945 5501
rect 9945 5475 9946 5501
rect 9918 5474 9946 5475
rect 9970 5501 9998 5502
rect 9970 5475 9971 5501
rect 9971 5475 9997 5501
rect 9997 5475 9998 5501
rect 9970 5474 9998 5475
rect 10022 5501 10050 5502
rect 10022 5475 10023 5501
rect 10023 5475 10049 5501
rect 10049 5475 10050 5501
rect 10022 5474 10050 5475
rect 2238 5109 2266 5110
rect 2238 5083 2239 5109
rect 2239 5083 2265 5109
rect 2265 5083 2266 5109
rect 2238 5082 2266 5083
rect 2290 5109 2318 5110
rect 2290 5083 2291 5109
rect 2291 5083 2317 5109
rect 2317 5083 2318 5109
rect 2290 5082 2318 5083
rect 2342 5109 2370 5110
rect 2342 5083 2343 5109
rect 2343 5083 2369 5109
rect 2369 5083 2370 5109
rect 2342 5082 2370 5083
rect 9918 4717 9946 4718
rect 9918 4691 9919 4717
rect 9919 4691 9945 4717
rect 9945 4691 9946 4717
rect 9918 4690 9946 4691
rect 9970 4717 9998 4718
rect 9970 4691 9971 4717
rect 9971 4691 9997 4717
rect 9997 4691 9998 4717
rect 9970 4690 9998 4691
rect 10022 4717 10050 4718
rect 10022 4691 10023 4717
rect 10023 4691 10049 4717
rect 10049 4691 10050 4717
rect 10022 4690 10050 4691
rect 2238 4325 2266 4326
rect 2238 4299 2239 4325
rect 2239 4299 2265 4325
rect 2265 4299 2266 4325
rect 2238 4298 2266 4299
rect 2290 4325 2318 4326
rect 2290 4299 2291 4325
rect 2291 4299 2317 4325
rect 2317 4299 2318 4325
rect 2290 4298 2318 4299
rect 2342 4325 2370 4326
rect 2342 4299 2343 4325
rect 2343 4299 2369 4325
rect 2369 4299 2370 4325
rect 2342 4298 2370 4299
rect 11438 8441 11466 8442
rect 11438 8415 11439 8441
rect 11439 8415 11465 8441
rect 11465 8415 11466 8441
rect 11438 8414 11466 8415
rect 12278 9673 12306 9674
rect 12278 9647 12279 9673
rect 12279 9647 12305 9673
rect 12305 9647 12306 9673
rect 12278 9646 12306 9647
rect 12670 10094 12698 10122
rect 12502 9814 12530 9842
rect 12614 9561 12642 9562
rect 12614 9535 12615 9561
rect 12615 9535 12641 9561
rect 12641 9535 12642 9561
rect 12614 9534 12642 9535
rect 13398 11185 13426 11186
rect 13398 11159 13399 11185
rect 13399 11159 13425 11185
rect 13425 11159 13426 11185
rect 13398 11158 13426 11159
rect 12838 10038 12866 10066
rect 12894 10542 12922 10570
rect 13734 10766 13762 10794
rect 14070 11158 14098 11186
rect 18830 11185 18858 11186
rect 18830 11159 18831 11185
rect 18831 11159 18857 11185
rect 18857 11159 18858 11185
rect 18830 11158 18858 11159
rect 14126 10766 14154 10794
rect 13622 10542 13650 10570
rect 13230 10094 13258 10122
rect 18830 10793 18858 10794
rect 18830 10767 18831 10793
rect 18831 10767 18857 10793
rect 18857 10767 18858 10793
rect 18830 10766 18858 10767
rect 20006 10766 20034 10794
rect 12726 9422 12754 9450
rect 12334 8918 12362 8946
rect 12838 9281 12866 9282
rect 12838 9255 12839 9281
rect 12839 9255 12865 9281
rect 12865 9255 12866 9281
rect 12838 9254 12866 9255
rect 12614 8918 12642 8946
rect 12726 9086 12754 9114
rect 12334 8777 12362 8778
rect 12334 8751 12335 8777
rect 12335 8751 12361 8777
rect 12361 8751 12362 8777
rect 12334 8750 12362 8751
rect 12278 8721 12306 8722
rect 12278 8695 12279 8721
rect 12279 8695 12305 8721
rect 12305 8695 12306 8721
rect 12278 8694 12306 8695
rect 12670 8750 12698 8778
rect 12334 8414 12362 8442
rect 11998 7966 12026 7994
rect 12614 7966 12642 7994
rect 17598 10597 17626 10598
rect 17598 10571 17599 10597
rect 17599 10571 17625 10597
rect 17625 10571 17626 10597
rect 17598 10570 17626 10571
rect 17650 10597 17678 10598
rect 17650 10571 17651 10597
rect 17651 10571 17677 10597
rect 17677 10571 17678 10597
rect 17650 10570 17678 10571
rect 17702 10597 17730 10598
rect 17702 10571 17703 10597
rect 17703 10571 17729 10597
rect 17729 10571 17730 10597
rect 17702 10570 17730 10571
rect 19950 10430 19978 10458
rect 14294 10065 14322 10066
rect 14294 10039 14295 10065
rect 14295 10039 14321 10065
rect 14321 10039 14322 10065
rect 14294 10038 14322 10039
rect 12894 9086 12922 9114
rect 13062 8694 13090 8722
rect 13062 8526 13090 8554
rect 12726 7769 12754 7770
rect 12726 7743 12727 7769
rect 12727 7743 12753 7769
rect 12753 7743 12754 7769
rect 12726 7742 12754 7743
rect 12894 8414 12922 8442
rect 11718 7630 11746 7658
rect 11494 7406 11522 7434
rect 12782 7657 12810 7658
rect 12782 7631 12783 7657
rect 12783 7631 12809 7657
rect 12809 7631 12810 7657
rect 12782 7630 12810 7631
rect 12334 7574 12362 7602
rect 11718 7406 11746 7434
rect 11998 7406 12026 7434
rect 13174 8918 13202 8946
rect 14070 8918 14098 8946
rect 17598 9813 17626 9814
rect 17598 9787 17599 9813
rect 17599 9787 17625 9813
rect 17625 9787 17626 9813
rect 17598 9786 17626 9787
rect 17650 9813 17678 9814
rect 17650 9787 17651 9813
rect 17651 9787 17677 9813
rect 17677 9787 17678 9813
rect 17650 9786 17678 9787
rect 17702 9813 17730 9814
rect 17702 9787 17703 9813
rect 17703 9787 17729 9813
rect 17729 9787 17730 9813
rect 17702 9786 17730 9787
rect 20006 10094 20034 10122
rect 18830 9646 18858 9674
rect 17598 9029 17626 9030
rect 17598 9003 17599 9029
rect 17599 9003 17625 9029
rect 17625 9003 17626 9029
rect 17598 9002 17626 9003
rect 17650 9029 17678 9030
rect 17650 9003 17651 9029
rect 17651 9003 17677 9029
rect 17677 9003 17678 9029
rect 17650 9002 17678 9003
rect 17702 9029 17730 9030
rect 17702 9003 17703 9029
rect 17703 9003 17729 9029
rect 17729 9003 17730 9029
rect 17702 9002 17730 9003
rect 18830 8833 18858 8834
rect 18830 8807 18831 8833
rect 18831 8807 18857 8833
rect 18857 8807 18858 8833
rect 18830 8806 18858 8807
rect 13342 8750 13370 8778
rect 13174 8441 13202 8442
rect 13174 8415 13175 8441
rect 13175 8415 13201 8441
rect 13201 8415 13202 8441
rect 13174 8414 13202 8415
rect 20006 8750 20034 8778
rect 18830 8441 18858 8442
rect 18830 8415 18831 8441
rect 18831 8415 18857 8441
rect 18857 8415 18858 8441
rect 18830 8414 18858 8415
rect 20006 8414 20034 8442
rect 17598 8245 17626 8246
rect 17598 8219 17599 8245
rect 17599 8219 17625 8245
rect 17625 8219 17626 8245
rect 17598 8218 17626 8219
rect 17650 8245 17678 8246
rect 17650 8219 17651 8245
rect 17651 8219 17677 8245
rect 17677 8219 17678 8245
rect 17650 8218 17678 8219
rect 17702 8245 17730 8246
rect 17702 8219 17703 8245
rect 17703 8219 17729 8245
rect 17729 8219 17730 8245
rect 17702 8218 17730 8219
rect 13174 7657 13202 7658
rect 13174 7631 13175 7657
rect 13175 7631 13201 7657
rect 13201 7631 13202 7657
rect 13174 7630 13202 7631
rect 13118 7601 13146 7602
rect 13118 7575 13119 7601
rect 13119 7575 13145 7601
rect 13145 7575 13146 7601
rect 13118 7574 13146 7575
rect 17598 7461 17626 7462
rect 17598 7435 17599 7461
rect 17599 7435 17625 7461
rect 17625 7435 17626 7461
rect 17598 7434 17626 7435
rect 17650 7461 17678 7462
rect 17650 7435 17651 7461
rect 17651 7435 17677 7461
rect 17677 7435 17678 7461
rect 17650 7434 17678 7435
rect 17702 7461 17730 7462
rect 17702 7435 17703 7461
rect 17703 7435 17729 7461
rect 17729 7435 17730 7461
rect 17702 7434 17730 7435
rect 13342 7406 13370 7434
rect 10878 6790 10906 6818
rect 11270 6817 11298 6818
rect 11270 6791 11271 6817
rect 11271 6791 11297 6817
rect 11297 6791 11298 6817
rect 11270 6790 11298 6791
rect 17598 6677 17626 6678
rect 17598 6651 17599 6677
rect 17599 6651 17625 6677
rect 17625 6651 17626 6677
rect 17598 6650 17626 6651
rect 17650 6677 17678 6678
rect 17650 6651 17651 6677
rect 17651 6651 17677 6677
rect 17677 6651 17678 6677
rect 17650 6650 17678 6651
rect 17702 6677 17730 6678
rect 17702 6651 17703 6677
rect 17703 6651 17729 6677
rect 17729 6651 17730 6677
rect 17702 6650 17730 6651
rect 9918 3933 9946 3934
rect 9918 3907 9919 3933
rect 9919 3907 9945 3933
rect 9945 3907 9946 3933
rect 9918 3906 9946 3907
rect 9970 3933 9998 3934
rect 9970 3907 9971 3933
rect 9971 3907 9997 3933
rect 9997 3907 9998 3933
rect 9970 3906 9998 3907
rect 10022 3933 10050 3934
rect 10022 3907 10023 3933
rect 10023 3907 10049 3933
rect 10049 3907 10050 3933
rect 10022 3906 10050 3907
rect 2238 3541 2266 3542
rect 2238 3515 2239 3541
rect 2239 3515 2265 3541
rect 2265 3515 2266 3541
rect 2238 3514 2266 3515
rect 2290 3541 2318 3542
rect 2290 3515 2291 3541
rect 2291 3515 2317 3541
rect 2317 3515 2318 3541
rect 2290 3514 2318 3515
rect 2342 3541 2370 3542
rect 2342 3515 2343 3541
rect 2343 3515 2369 3541
rect 2369 3515 2370 3541
rect 2342 3514 2370 3515
rect 9918 3149 9946 3150
rect 9918 3123 9919 3149
rect 9919 3123 9945 3149
rect 9945 3123 9946 3149
rect 9918 3122 9946 3123
rect 9970 3149 9998 3150
rect 9970 3123 9971 3149
rect 9971 3123 9997 3149
rect 9997 3123 9998 3149
rect 9970 3122 9998 3123
rect 10022 3149 10050 3150
rect 10022 3123 10023 3149
rect 10023 3123 10049 3149
rect 10049 3123 10050 3149
rect 10022 3122 10050 3123
rect 2238 2757 2266 2758
rect 2238 2731 2239 2757
rect 2239 2731 2265 2757
rect 2265 2731 2266 2757
rect 2238 2730 2266 2731
rect 2290 2757 2318 2758
rect 2290 2731 2291 2757
rect 2291 2731 2317 2757
rect 2317 2731 2318 2757
rect 2290 2730 2318 2731
rect 2342 2757 2370 2758
rect 2342 2731 2343 2757
rect 2343 2731 2369 2757
rect 2369 2731 2370 2757
rect 2342 2730 2370 2731
rect 9918 2365 9946 2366
rect 9918 2339 9919 2365
rect 9919 2339 9945 2365
rect 9945 2339 9946 2365
rect 9918 2338 9946 2339
rect 9970 2365 9998 2366
rect 9970 2339 9971 2365
rect 9971 2339 9997 2365
rect 9997 2339 9998 2365
rect 9970 2338 9998 2339
rect 10022 2365 10050 2366
rect 10022 2339 10023 2365
rect 10023 2339 10049 2365
rect 10049 2339 10050 2365
rect 10022 2338 10050 2339
rect 10486 2142 10514 2170
rect 17598 5893 17626 5894
rect 17598 5867 17599 5893
rect 17599 5867 17625 5893
rect 17625 5867 17626 5893
rect 17598 5866 17626 5867
rect 17650 5893 17678 5894
rect 17650 5867 17651 5893
rect 17651 5867 17677 5893
rect 17677 5867 17678 5893
rect 17650 5866 17678 5867
rect 17702 5893 17730 5894
rect 17702 5867 17703 5893
rect 17703 5867 17729 5893
rect 17729 5867 17730 5893
rect 17702 5866 17730 5867
rect 17598 5109 17626 5110
rect 17598 5083 17599 5109
rect 17599 5083 17625 5109
rect 17625 5083 17626 5109
rect 17598 5082 17626 5083
rect 17650 5109 17678 5110
rect 17650 5083 17651 5109
rect 17651 5083 17677 5109
rect 17677 5083 17678 5109
rect 17650 5082 17678 5083
rect 17702 5109 17730 5110
rect 17702 5083 17703 5109
rect 17703 5083 17729 5109
rect 17729 5083 17730 5109
rect 17702 5082 17730 5083
rect 17598 4325 17626 4326
rect 17598 4299 17599 4325
rect 17599 4299 17625 4325
rect 17625 4299 17626 4325
rect 17598 4298 17626 4299
rect 17650 4325 17678 4326
rect 17650 4299 17651 4325
rect 17651 4299 17677 4325
rect 17677 4299 17678 4325
rect 17650 4298 17678 4299
rect 17702 4325 17730 4326
rect 17702 4299 17703 4325
rect 17703 4299 17729 4325
rect 17729 4299 17730 4325
rect 17702 4298 17730 4299
rect 2238 1973 2266 1974
rect 2238 1947 2239 1973
rect 2239 1947 2265 1973
rect 2265 1947 2266 1973
rect 2238 1946 2266 1947
rect 2290 1973 2318 1974
rect 2290 1947 2291 1973
rect 2291 1947 2317 1973
rect 2317 1947 2318 1973
rect 2290 1946 2318 1947
rect 2342 1973 2370 1974
rect 2342 1947 2343 1973
rect 2343 1947 2369 1973
rect 2369 1947 2370 1973
rect 2342 1946 2370 1947
rect 10878 2169 10906 2170
rect 10878 2143 10879 2169
rect 10879 2143 10905 2169
rect 10905 2143 10906 2169
rect 10878 2142 10906 2143
rect 10766 2030 10794 2058
rect 9918 1581 9946 1582
rect 9918 1555 9919 1581
rect 9919 1555 9945 1581
rect 9945 1555 9946 1581
rect 9918 1554 9946 1555
rect 9970 1581 9998 1582
rect 9970 1555 9971 1581
rect 9971 1555 9997 1581
rect 9997 1555 9998 1581
rect 9970 1554 9998 1555
rect 10022 1581 10050 1582
rect 10022 1555 10023 1581
rect 10023 1555 10049 1581
rect 10049 1555 10050 1581
rect 10022 1554 10050 1555
rect 11382 2057 11410 2058
rect 11382 2031 11383 2057
rect 11383 2031 11409 2057
rect 11409 2031 11410 2057
rect 11382 2030 11410 2031
rect 17598 3541 17626 3542
rect 17598 3515 17599 3541
rect 17599 3515 17625 3541
rect 17625 3515 17626 3541
rect 17598 3514 17626 3515
rect 17650 3541 17678 3542
rect 17650 3515 17651 3541
rect 17651 3515 17677 3541
rect 17677 3515 17678 3541
rect 17650 3514 17678 3515
rect 17702 3541 17730 3542
rect 17702 3515 17703 3541
rect 17703 3515 17729 3541
rect 17729 3515 17730 3541
rect 17702 3514 17730 3515
rect 17598 2757 17626 2758
rect 17598 2731 17599 2757
rect 17599 2731 17625 2757
rect 17625 2731 17626 2757
rect 17598 2730 17626 2731
rect 17650 2757 17678 2758
rect 17650 2731 17651 2757
rect 17651 2731 17677 2757
rect 17677 2731 17678 2757
rect 17650 2730 17678 2731
rect 17702 2757 17730 2758
rect 17702 2731 17703 2757
rect 17703 2731 17729 2757
rect 17729 2731 17730 2757
rect 17702 2730 17730 2731
rect 17598 1973 17626 1974
rect 17598 1947 17599 1973
rect 17599 1947 17625 1973
rect 17625 1947 17626 1973
rect 17598 1946 17626 1947
rect 17650 1973 17678 1974
rect 17650 1947 17651 1973
rect 17651 1947 17677 1973
rect 17677 1947 17678 1973
rect 17650 1946 17678 1947
rect 17702 1973 17730 1974
rect 17702 1947 17703 1973
rect 17703 1947 17729 1973
rect 17729 1947 17730 1973
rect 17702 1946 17730 1947
<< metal3 >>
rect 2233 19194 2238 19222
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2370 19194 2375 19222
rect 17593 19194 17598 19222
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17730 19194 17735 19222
rect 11769 19110 11774 19138
rect 11802 19110 12782 19138
rect 12810 19110 12815 19138
rect 9417 18942 9422 18970
rect 9450 18942 10374 18970
rect 10402 18942 10407 18970
rect 9913 18802 9918 18830
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 10050 18802 10055 18830
rect 8409 18718 8414 18746
rect 8442 18718 9198 18746
rect 9226 18718 9231 18746
rect 10425 18718 10430 18746
rect 10458 18718 11046 18746
rect 11074 18718 11079 18746
rect 12105 18718 12110 18746
rect 12138 18718 13118 18746
rect 13146 18718 13151 18746
rect 20600 18522 21000 18536
rect 20113 18494 20118 18522
rect 20146 18494 21000 18522
rect 20600 18480 21000 18494
rect 2233 18410 2238 18438
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2370 18410 2375 18438
rect 17593 18410 17598 18438
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17730 18410 17735 18438
rect 9913 18018 9918 18046
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 10050 18018 10055 18046
rect 2233 17626 2238 17654
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2370 17626 2375 17654
rect 17593 17626 17598 17654
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17730 17626 17735 17654
rect 9913 17234 9918 17262
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 10050 17234 10055 17262
rect 2233 16842 2238 16870
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2370 16842 2375 16870
rect 17593 16842 17598 16870
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17730 16842 17735 16870
rect 9913 16450 9918 16478
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 10050 16450 10055 16478
rect 2233 16058 2238 16086
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2370 16058 2375 16086
rect 17593 16058 17598 16086
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17730 16058 17735 16086
rect 9913 15666 9918 15694
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 10050 15666 10055 15694
rect 2233 15274 2238 15302
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2370 15274 2375 15302
rect 17593 15274 17598 15302
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17730 15274 17735 15302
rect 9913 14882 9918 14910
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 10050 14882 10055 14910
rect 2233 14490 2238 14518
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2370 14490 2375 14518
rect 17593 14490 17598 14518
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17730 14490 17735 14518
rect 9913 14098 9918 14126
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 10050 14098 10055 14126
rect 0 13818 400 13832
rect 0 13790 2086 13818
rect 2114 13790 2119 13818
rect 0 13776 400 13790
rect 2233 13706 2238 13734
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2370 13706 2375 13734
rect 17593 13706 17598 13734
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17730 13706 17735 13734
rect 8241 13510 8246 13538
rect 8274 13510 8750 13538
rect 8778 13510 8783 13538
rect 10145 13510 10150 13538
rect 10178 13510 11830 13538
rect 11858 13510 13230 13538
rect 13258 13510 13263 13538
rect 20600 13482 21000 13496
rect 6561 13454 6566 13482
rect 6594 13454 7070 13482
rect 7098 13454 8862 13482
rect 8890 13454 9086 13482
rect 9114 13454 9119 13482
rect 13169 13454 13174 13482
rect 13202 13454 13790 13482
rect 13818 13454 13823 13482
rect 13897 13454 13902 13482
rect 13930 13454 18942 13482
rect 18970 13454 18975 13482
rect 19945 13454 19950 13482
rect 19978 13454 21000 13482
rect 9086 13426 9114 13454
rect 20600 13440 21000 13454
rect 8521 13398 8526 13426
rect 8554 13398 8750 13426
rect 8778 13398 8783 13426
rect 9086 13398 9422 13426
rect 9450 13398 9455 13426
rect 9913 13314 9918 13342
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 10050 13314 10055 13342
rect 7457 13230 7462 13258
rect 7490 13230 8190 13258
rect 8218 13230 8223 13258
rect 12161 13230 12166 13258
rect 12194 13230 12614 13258
rect 12642 13230 12647 13258
rect 15946 13230 18830 13258
rect 18858 13230 18863 13258
rect 15946 13202 15974 13230
rect 8297 13174 8302 13202
rect 8330 13174 9478 13202
rect 9506 13174 9511 13202
rect 14401 13174 14406 13202
rect 14434 13174 15974 13202
rect 20600 13146 21000 13160
rect 8129 13118 8134 13146
rect 8162 13118 8918 13146
rect 8946 13118 8951 13146
rect 13785 13118 13790 13146
rect 13818 13118 14070 13146
rect 14098 13118 14294 13146
rect 14322 13118 18830 13146
rect 18858 13118 18863 13146
rect 20001 13118 20006 13146
rect 20034 13118 21000 13146
rect 20600 13104 21000 13118
rect 2233 12922 2238 12950
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2370 12922 2375 12950
rect 17593 12922 17598 12950
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17730 12922 17735 12950
rect 20600 12810 21000 12824
rect 4186 12782 4998 12810
rect 5026 12782 5950 12810
rect 5978 12782 5983 12810
rect 8913 12782 8918 12810
rect 8946 12782 9254 12810
rect 9282 12782 9287 12810
rect 11769 12782 11774 12810
rect 11802 12782 12166 12810
rect 12194 12782 12199 12810
rect 19945 12782 19950 12810
rect 19978 12782 21000 12810
rect 4186 12754 4214 12782
rect 20600 12768 21000 12782
rect 2137 12726 2142 12754
rect 2170 12726 4214 12754
rect 10761 12726 10766 12754
rect 10794 12726 11270 12754
rect 11298 12726 11303 12754
rect 13505 12726 13510 12754
rect 13538 12726 14014 12754
rect 14042 12726 18830 12754
rect 18858 12726 18863 12754
rect 6057 12670 6062 12698
rect 6090 12670 6958 12698
rect 6986 12670 6991 12698
rect 11270 12642 11298 12726
rect 6449 12614 6454 12642
rect 6482 12614 6790 12642
rect 6818 12614 6823 12642
rect 11270 12614 12390 12642
rect 12418 12614 14238 12642
rect 14266 12614 14630 12642
rect 14658 12614 14663 12642
rect 9913 12530 9918 12558
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 10050 12530 10055 12558
rect 0 12474 400 12488
rect 20600 12474 21000 12488
rect 0 12446 966 12474
rect 994 12446 999 12474
rect 13225 12446 13230 12474
rect 13258 12446 13622 12474
rect 13650 12446 13655 12474
rect 20001 12446 20006 12474
rect 20034 12446 21000 12474
rect 0 12432 400 12446
rect 20600 12432 21000 12446
rect 7009 12390 7014 12418
rect 7042 12390 7686 12418
rect 7714 12390 7719 12418
rect 11774 12390 12894 12418
rect 12922 12390 12927 12418
rect 11774 12362 11802 12390
rect 7625 12334 7630 12362
rect 7658 12334 9030 12362
rect 9058 12334 9758 12362
rect 9786 12334 9791 12362
rect 11657 12334 11662 12362
rect 11690 12334 11774 12362
rect 11802 12334 11807 12362
rect 12385 12334 12390 12362
rect 12418 12334 13174 12362
rect 13202 12334 13207 12362
rect 6337 12278 6342 12306
rect 6370 12278 6790 12306
rect 6818 12278 6823 12306
rect 9865 12278 9870 12306
rect 9898 12278 10654 12306
rect 10682 12278 10687 12306
rect 7065 12222 7070 12250
rect 7098 12222 7630 12250
rect 7658 12222 7663 12250
rect 2233 12138 2238 12166
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2370 12138 2375 12166
rect 17593 12138 17598 12166
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17730 12138 17735 12166
rect 10817 12110 10822 12138
rect 10850 12110 11494 12138
rect 11522 12110 11527 12138
rect 6897 11998 6902 12026
rect 6930 11998 7518 12026
rect 7546 11998 10990 12026
rect 11018 11998 11023 12026
rect 11265 11998 11270 12026
rect 11298 11998 11718 12026
rect 11746 11998 11751 12026
rect 9697 11942 9702 11970
rect 9730 11942 10710 11970
rect 10738 11942 11886 11970
rect 11914 11942 13342 11970
rect 13370 11942 13375 11970
rect 7546 11886 7854 11914
rect 7882 11886 8134 11914
rect 8162 11886 8167 11914
rect 11153 11886 11158 11914
rect 11186 11886 11438 11914
rect 11466 11886 11471 11914
rect 7546 11802 7574 11886
rect 10537 11830 10542 11858
rect 10570 11830 10822 11858
rect 10850 11830 10855 11858
rect 11097 11830 11102 11858
rect 11130 11830 11606 11858
rect 11634 11830 11639 11858
rect 7401 11774 7406 11802
rect 7434 11774 7574 11802
rect 10705 11774 10710 11802
rect 10738 11774 11774 11802
rect 11802 11774 12054 11802
rect 12082 11774 12087 11802
rect 9913 11746 9918 11774
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 10050 11746 10055 11774
rect 8969 11718 8974 11746
rect 9002 11718 9814 11746
rect 9842 11718 9847 11746
rect 7457 11606 7462 11634
rect 7490 11606 7574 11634
rect 7602 11606 7607 11634
rect 8465 11606 8470 11634
rect 8498 11606 8806 11634
rect 8834 11606 8839 11634
rect 8577 11438 8582 11466
rect 8610 11438 8862 11466
rect 8890 11438 9198 11466
rect 9226 11438 9231 11466
rect 2233 11354 2238 11382
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2370 11354 2375 11382
rect 17593 11354 17598 11382
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17730 11354 17735 11382
rect 7289 11158 7294 11186
rect 7322 11158 8134 11186
rect 8162 11158 8167 11186
rect 10649 11158 10654 11186
rect 10682 11158 11438 11186
rect 11466 11158 11471 11186
rect 12217 11158 12222 11186
rect 12250 11158 12670 11186
rect 12698 11158 12703 11186
rect 13393 11158 13398 11186
rect 13426 11158 14070 11186
rect 14098 11158 18830 11186
rect 18858 11158 18863 11186
rect 6393 11102 6398 11130
rect 6426 11102 7854 11130
rect 7882 11102 10542 11130
rect 10570 11102 10575 11130
rect 7121 11046 7126 11074
rect 7154 11046 7462 11074
rect 7490 11046 7686 11074
rect 7714 11046 7719 11074
rect 6449 10990 6454 11018
rect 6482 10990 6622 11018
rect 6650 10990 7574 11018
rect 7602 10990 7910 11018
rect 7938 10990 7943 11018
rect 8078 10990 9058 11018
rect 8078 10962 8106 10990
rect 9030 10962 9058 10990
rect 9913 10962 9918 10990
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 10050 10962 10055 10990
rect 6561 10934 6566 10962
rect 6594 10934 7126 10962
rect 7154 10934 8106 10962
rect 8185 10934 8190 10962
rect 8218 10934 8582 10962
rect 8610 10934 8615 10962
rect 9025 10934 9030 10962
rect 9058 10934 9063 10962
rect 6785 10878 6790 10906
rect 6818 10878 7630 10906
rect 7658 10878 7663 10906
rect 9809 10878 9814 10906
rect 9842 10878 11046 10906
rect 11074 10878 11079 10906
rect 8297 10822 8302 10850
rect 8330 10822 9478 10850
rect 9506 10822 9511 10850
rect 20600 10794 21000 10808
rect 2137 10766 2142 10794
rect 2170 10766 4830 10794
rect 4858 10766 4863 10794
rect 7961 10766 7966 10794
rect 7994 10766 8414 10794
rect 8442 10766 8447 10794
rect 13729 10766 13734 10794
rect 13762 10766 14126 10794
rect 14154 10766 18830 10794
rect 18858 10766 18863 10794
rect 20001 10766 20006 10794
rect 20034 10766 21000 10794
rect 20600 10752 21000 10766
rect 2081 10710 2086 10738
rect 2114 10710 8806 10738
rect 8834 10710 8839 10738
rect 9753 10710 9758 10738
rect 9786 10710 10822 10738
rect 10850 10710 10855 10738
rect 6617 10654 6622 10682
rect 6650 10654 8078 10682
rect 8106 10654 8111 10682
rect 8353 10654 8358 10682
rect 8386 10654 9198 10682
rect 9226 10654 9231 10682
rect 6897 10598 6902 10626
rect 6930 10598 7742 10626
rect 7770 10598 9814 10626
rect 9842 10598 9847 10626
rect 2233 10570 2238 10598
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2370 10570 2375 10598
rect 17593 10570 17598 10598
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17730 10570 17735 10598
rect 8465 10542 8470 10570
rect 8498 10542 9086 10570
rect 9114 10542 9478 10570
rect 9506 10542 9511 10570
rect 12889 10542 12894 10570
rect 12922 10542 13622 10570
rect 13650 10542 13655 10570
rect 0 10458 400 10472
rect 20600 10458 21000 10472
rect 0 10430 966 10458
rect 994 10430 999 10458
rect 6785 10430 6790 10458
rect 6818 10430 7350 10458
rect 7378 10430 8246 10458
rect 8274 10430 8414 10458
rect 8442 10430 8447 10458
rect 9641 10430 9646 10458
rect 9674 10430 9814 10458
rect 9842 10430 9847 10458
rect 19945 10430 19950 10458
rect 19978 10430 21000 10458
rect 0 10416 400 10430
rect 20600 10416 21000 10430
rect 4825 10374 4830 10402
rect 4858 10374 6902 10402
rect 6930 10374 6935 10402
rect 7546 10374 9086 10402
rect 9114 10374 9119 10402
rect 7546 10346 7574 10374
rect 7289 10318 7294 10346
rect 7322 10318 7574 10346
rect 7905 10318 7910 10346
rect 7938 10318 8582 10346
rect 8610 10318 8615 10346
rect 6113 10262 6118 10290
rect 6146 10262 6846 10290
rect 6874 10262 6879 10290
rect 9913 10178 9918 10206
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 10050 10178 10055 10206
rect 20600 10122 21000 10136
rect 5049 10094 5054 10122
rect 5082 10094 6958 10122
rect 6986 10094 7294 10122
rect 7322 10094 7327 10122
rect 12665 10094 12670 10122
rect 12698 10094 13230 10122
rect 13258 10094 13454 10122
rect 20001 10094 20006 10122
rect 20034 10094 21000 10122
rect 13426 10066 13454 10094
rect 20600 10080 21000 10094
rect 7009 10038 7014 10066
rect 7042 10038 8190 10066
rect 8218 10038 8223 10066
rect 8297 10038 8302 10066
rect 8330 10038 8750 10066
rect 8778 10038 8783 10066
rect 8969 10038 8974 10066
rect 9002 10038 9310 10066
rect 9338 10038 10094 10066
rect 10122 10038 10127 10066
rect 11825 10038 11830 10066
rect 11858 10038 12838 10066
rect 12866 10038 12871 10066
rect 13426 10038 14294 10066
rect 14322 10038 14327 10066
rect 6398 9982 6566 10010
rect 6594 9982 7462 10010
rect 7490 9982 7495 10010
rect 8465 9982 8470 10010
rect 8498 9982 9198 10010
rect 9226 9982 9590 10010
rect 9618 9982 9623 10010
rect 10313 9982 10318 10010
rect 10346 9982 11494 10010
rect 11522 9982 12166 10010
rect 12194 9982 12199 10010
rect 6398 9842 6426 9982
rect 8017 9926 8022 9954
rect 8050 9926 9758 9954
rect 9786 9926 9791 9954
rect 11041 9926 11046 9954
rect 11074 9926 11214 9954
rect 11242 9926 11247 9954
rect 9417 9870 9422 9898
rect 9450 9870 10150 9898
rect 10178 9870 10183 9898
rect 6393 9814 6398 9842
rect 6426 9814 6431 9842
rect 8297 9814 8302 9842
rect 8330 9814 12502 9842
rect 12530 9814 12535 9842
rect 2233 9786 2238 9814
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2370 9786 2375 9814
rect 17593 9786 17598 9814
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17730 9786 17735 9814
rect 7345 9702 7350 9730
rect 7378 9702 7630 9730
rect 7658 9702 7663 9730
rect 9977 9702 9982 9730
rect 10010 9702 10318 9730
rect 10346 9702 10351 9730
rect 7457 9646 7462 9674
rect 7490 9646 8526 9674
rect 8554 9646 8559 9674
rect 11377 9646 11382 9674
rect 11410 9646 12278 9674
rect 12306 9646 18830 9674
rect 18858 9646 18863 9674
rect 7849 9590 7854 9618
rect 7882 9590 8022 9618
rect 8050 9590 8055 9618
rect 9361 9590 9366 9618
rect 9394 9590 10206 9618
rect 10234 9590 11662 9618
rect 11690 9590 11695 9618
rect 7681 9534 7686 9562
rect 7714 9534 8022 9562
rect 8050 9534 8055 9562
rect 8745 9534 8750 9562
rect 8778 9534 11270 9562
rect 11298 9534 12614 9562
rect 12642 9534 12647 9562
rect 7737 9478 7742 9506
rect 7770 9478 8134 9506
rect 8162 9478 8167 9506
rect 10486 9422 12726 9450
rect 12754 9422 12759 9450
rect 9913 9394 9918 9422
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 10050 9394 10055 9422
rect 10486 9394 10514 9422
rect 10481 9366 10486 9394
rect 10514 9366 10519 9394
rect 7905 9310 7910 9338
rect 7938 9310 8694 9338
rect 8722 9310 8727 9338
rect 7910 9282 7938 9310
rect 7681 9254 7686 9282
rect 7714 9254 7938 9282
rect 11601 9254 11606 9282
rect 11634 9254 12054 9282
rect 12082 9254 12838 9282
rect 12866 9254 12871 9282
rect 2137 9198 2142 9226
rect 2170 9198 4998 9226
rect 5026 9198 5031 9226
rect 7121 9198 7126 9226
rect 7154 9198 7406 9226
rect 7434 9198 10094 9226
rect 10122 9198 10127 9226
rect 7009 9142 7014 9170
rect 7042 9142 7742 9170
rect 7770 9142 7775 9170
rect 9473 9142 9478 9170
rect 9506 9142 10430 9170
rect 10458 9142 10463 9170
rect 0 9114 400 9128
rect 0 9086 966 9114
rect 994 9086 999 9114
rect 8409 9086 8414 9114
rect 8442 9086 9086 9114
rect 9114 9086 9758 9114
rect 9786 9086 9791 9114
rect 10873 9086 10878 9114
rect 10906 9086 11046 9114
rect 11074 9086 11079 9114
rect 12721 9086 12726 9114
rect 12754 9086 12894 9114
rect 12922 9086 12927 9114
rect 0 9072 400 9086
rect 9193 9030 9198 9058
rect 9226 9030 9590 9058
rect 9618 9030 10206 9058
rect 10234 9030 10239 9058
rect 2233 9002 2238 9030
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2370 9002 2375 9030
rect 17593 9002 17598 9030
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17730 9002 17735 9030
rect 5889 8974 5894 9002
rect 5922 8974 9030 9002
rect 9058 8974 9063 9002
rect 7793 8918 7798 8946
rect 7826 8918 12334 8946
rect 12362 8918 12614 8946
rect 12642 8918 12647 8946
rect 13169 8918 13174 8946
rect 13202 8918 14070 8946
rect 14098 8918 15974 8946
rect 961 8862 966 8890
rect 994 8862 999 8890
rect 9081 8862 9086 8890
rect 9114 8862 9534 8890
rect 9562 8862 9567 8890
rect 0 8778 400 8792
rect 966 8778 994 8862
rect 15946 8834 15974 8918
rect 2137 8806 2142 8834
rect 2170 8806 6342 8834
rect 6370 8806 6375 8834
rect 15946 8806 18830 8834
rect 18858 8806 18863 8834
rect 20600 8778 21000 8792
rect 0 8750 994 8778
rect 4993 8750 4998 8778
rect 5026 8750 6286 8778
rect 6314 8750 6510 8778
rect 6538 8750 6543 8778
rect 8003 8750 8022 8778
rect 8050 8750 8055 8778
rect 8409 8750 8414 8778
rect 8442 8750 8750 8778
rect 8778 8750 8783 8778
rect 11102 8750 12334 8778
rect 12362 8750 12367 8778
rect 12665 8750 12670 8778
rect 12698 8750 13342 8778
rect 13370 8750 13375 8778
rect 20001 8750 20006 8778
rect 20034 8750 21000 8778
rect 0 8736 400 8750
rect 11102 8722 11130 8750
rect 20600 8736 21000 8750
rect 5777 8694 5782 8722
rect 5810 8694 7518 8722
rect 7546 8694 7551 8722
rect 8073 8694 8078 8722
rect 8106 8694 8302 8722
rect 8330 8694 9142 8722
rect 9170 8694 9175 8722
rect 9921 8694 9926 8722
rect 9954 8694 11102 8722
rect 11130 8694 11135 8722
rect 12273 8694 12278 8722
rect 12306 8694 13062 8722
rect 13090 8694 13095 8722
rect 6169 8638 6174 8666
rect 6202 8638 7014 8666
rect 7042 8638 7047 8666
rect 9913 8610 9918 8638
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 10050 8610 10055 8638
rect 8017 8526 8022 8554
rect 8050 8526 8694 8554
rect 8722 8526 8727 8554
rect 13057 8526 13062 8554
rect 13090 8526 15974 8554
rect 0 8442 400 8456
rect 15946 8442 15974 8526
rect 20600 8442 21000 8456
rect 0 8414 966 8442
rect 994 8414 999 8442
rect 2137 8414 2142 8442
rect 2170 8414 5782 8442
rect 5810 8414 5815 8442
rect 8857 8414 8862 8442
rect 8890 8414 9366 8442
rect 9394 8414 9399 8442
rect 10985 8414 10990 8442
rect 11018 8414 11438 8442
rect 11466 8414 11471 8442
rect 12329 8414 12334 8442
rect 12362 8414 12894 8442
rect 12922 8414 13174 8442
rect 13202 8414 13207 8442
rect 15946 8414 18830 8442
rect 18858 8414 18863 8442
rect 20001 8414 20006 8442
rect 20034 8414 21000 8442
rect 0 8400 400 8414
rect 20600 8400 21000 8414
rect 9977 8358 9982 8386
rect 10010 8358 10542 8386
rect 10570 8358 10575 8386
rect 2233 8218 2238 8246
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2370 8218 2375 8246
rect 17593 8218 17598 8246
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17730 8218 17735 8246
rect 6449 8022 6454 8050
rect 6482 8022 6790 8050
rect 6818 8022 6823 8050
rect 9249 8022 9254 8050
rect 9282 8022 10038 8050
rect 10066 8022 10071 8050
rect 7345 7966 7350 7994
rect 7378 7966 8134 7994
rect 8162 7966 8167 7994
rect 10873 7966 10878 7994
rect 10906 7966 11998 7994
rect 12026 7966 12614 7994
rect 12642 7966 12647 7994
rect 9025 7910 9030 7938
rect 9058 7910 10710 7938
rect 10738 7910 10743 7938
rect 9913 7826 9918 7854
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 10050 7826 10055 7854
rect 10313 7798 10318 7826
rect 10346 7798 10598 7826
rect 10626 7798 10631 7826
rect 10145 7742 10150 7770
rect 10178 7742 12726 7770
rect 12754 7742 12759 7770
rect 7009 7630 7014 7658
rect 7042 7630 7462 7658
rect 7490 7630 8750 7658
rect 8778 7630 8783 7658
rect 9809 7630 9814 7658
rect 9842 7630 10430 7658
rect 10458 7630 10710 7658
rect 10738 7630 11718 7658
rect 11746 7630 11751 7658
rect 12777 7630 12782 7658
rect 12810 7630 13174 7658
rect 13202 7630 13207 7658
rect 8353 7574 8358 7602
rect 8386 7574 9030 7602
rect 9058 7574 9063 7602
rect 12329 7574 12334 7602
rect 12362 7574 13118 7602
rect 13146 7574 13151 7602
rect 2233 7434 2238 7462
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2370 7434 2375 7462
rect 17593 7434 17598 7462
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17730 7434 17735 7462
rect 11489 7406 11494 7434
rect 11522 7406 11718 7434
rect 11746 7406 11998 7434
rect 12026 7406 13342 7434
rect 13370 7406 13375 7434
rect 9913 7042 9918 7070
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 10050 7042 10055 7070
rect 10873 6790 10878 6818
rect 10906 6790 11270 6818
rect 11298 6790 11303 6818
rect 2233 6650 2238 6678
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2370 6650 2375 6678
rect 17593 6650 17598 6678
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17730 6650 17735 6678
rect 9913 6258 9918 6286
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 10050 6258 10055 6286
rect 2233 5866 2238 5894
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2370 5866 2375 5894
rect 17593 5866 17598 5894
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17730 5866 17735 5894
rect 9913 5474 9918 5502
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 10050 5474 10055 5502
rect 2233 5082 2238 5110
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2370 5082 2375 5110
rect 17593 5082 17598 5110
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17730 5082 17735 5110
rect 9913 4690 9918 4718
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 10050 4690 10055 4718
rect 2233 4298 2238 4326
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2370 4298 2375 4326
rect 17593 4298 17598 4326
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17730 4298 17735 4326
rect 9913 3906 9918 3934
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 10050 3906 10055 3934
rect 2233 3514 2238 3542
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2370 3514 2375 3542
rect 17593 3514 17598 3542
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17730 3514 17735 3542
rect 9913 3122 9918 3150
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 10050 3122 10055 3150
rect 2233 2730 2238 2758
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2370 2730 2375 2758
rect 17593 2730 17598 2758
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17730 2730 17735 2758
rect 9913 2338 9918 2366
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 10050 2338 10055 2366
rect 10481 2142 10486 2170
rect 10514 2142 10878 2170
rect 10906 2142 10911 2170
rect 10761 2030 10766 2058
rect 10794 2030 11382 2058
rect 11410 2030 11415 2058
rect 2233 1946 2238 1974
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2370 1946 2375 1974
rect 17593 1946 17598 1974
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17730 1946 17735 1974
rect 9913 1554 9918 1582
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 10050 1554 10055 1582
<< via3 >>
rect 2238 19194 2266 19222
rect 2290 19194 2318 19222
rect 2342 19194 2370 19222
rect 17598 19194 17626 19222
rect 17650 19194 17678 19222
rect 17702 19194 17730 19222
rect 9918 18802 9946 18830
rect 9970 18802 9998 18830
rect 10022 18802 10050 18830
rect 2238 18410 2266 18438
rect 2290 18410 2318 18438
rect 2342 18410 2370 18438
rect 17598 18410 17626 18438
rect 17650 18410 17678 18438
rect 17702 18410 17730 18438
rect 9918 18018 9946 18046
rect 9970 18018 9998 18046
rect 10022 18018 10050 18046
rect 2238 17626 2266 17654
rect 2290 17626 2318 17654
rect 2342 17626 2370 17654
rect 17598 17626 17626 17654
rect 17650 17626 17678 17654
rect 17702 17626 17730 17654
rect 9918 17234 9946 17262
rect 9970 17234 9998 17262
rect 10022 17234 10050 17262
rect 2238 16842 2266 16870
rect 2290 16842 2318 16870
rect 2342 16842 2370 16870
rect 17598 16842 17626 16870
rect 17650 16842 17678 16870
rect 17702 16842 17730 16870
rect 9918 16450 9946 16478
rect 9970 16450 9998 16478
rect 10022 16450 10050 16478
rect 2238 16058 2266 16086
rect 2290 16058 2318 16086
rect 2342 16058 2370 16086
rect 17598 16058 17626 16086
rect 17650 16058 17678 16086
rect 17702 16058 17730 16086
rect 9918 15666 9946 15694
rect 9970 15666 9998 15694
rect 10022 15666 10050 15694
rect 2238 15274 2266 15302
rect 2290 15274 2318 15302
rect 2342 15274 2370 15302
rect 17598 15274 17626 15302
rect 17650 15274 17678 15302
rect 17702 15274 17730 15302
rect 9918 14882 9946 14910
rect 9970 14882 9998 14910
rect 10022 14882 10050 14910
rect 2238 14490 2266 14518
rect 2290 14490 2318 14518
rect 2342 14490 2370 14518
rect 17598 14490 17626 14518
rect 17650 14490 17678 14518
rect 17702 14490 17730 14518
rect 9918 14098 9946 14126
rect 9970 14098 9998 14126
rect 10022 14098 10050 14126
rect 2238 13706 2266 13734
rect 2290 13706 2318 13734
rect 2342 13706 2370 13734
rect 17598 13706 17626 13734
rect 17650 13706 17678 13734
rect 17702 13706 17730 13734
rect 9918 13314 9946 13342
rect 9970 13314 9998 13342
rect 10022 13314 10050 13342
rect 2238 12922 2266 12950
rect 2290 12922 2318 12950
rect 2342 12922 2370 12950
rect 17598 12922 17626 12950
rect 17650 12922 17678 12950
rect 17702 12922 17730 12950
rect 9918 12530 9946 12558
rect 9970 12530 9998 12558
rect 10022 12530 10050 12558
rect 2238 12138 2266 12166
rect 2290 12138 2318 12166
rect 2342 12138 2370 12166
rect 17598 12138 17626 12166
rect 17650 12138 17678 12166
rect 17702 12138 17730 12166
rect 9918 11746 9946 11774
rect 9970 11746 9998 11774
rect 10022 11746 10050 11774
rect 2238 11354 2266 11382
rect 2290 11354 2318 11382
rect 2342 11354 2370 11382
rect 17598 11354 17626 11382
rect 17650 11354 17678 11382
rect 17702 11354 17730 11382
rect 9918 10962 9946 10990
rect 9970 10962 9998 10990
rect 10022 10962 10050 10990
rect 2238 10570 2266 10598
rect 2290 10570 2318 10598
rect 2342 10570 2370 10598
rect 17598 10570 17626 10598
rect 17650 10570 17678 10598
rect 17702 10570 17730 10598
rect 9918 10178 9946 10206
rect 9970 10178 9998 10206
rect 10022 10178 10050 10206
rect 2238 9786 2266 9814
rect 2290 9786 2318 9814
rect 2342 9786 2370 9814
rect 17598 9786 17626 9814
rect 17650 9786 17678 9814
rect 17702 9786 17730 9814
rect 8022 9590 8050 9618
rect 9918 9394 9946 9422
rect 9970 9394 9998 9422
rect 10022 9394 10050 9422
rect 2238 9002 2266 9030
rect 2290 9002 2318 9030
rect 2342 9002 2370 9030
rect 17598 9002 17626 9030
rect 17650 9002 17678 9030
rect 17702 9002 17730 9030
rect 8022 8750 8050 8778
rect 9918 8610 9946 8638
rect 9970 8610 9998 8638
rect 10022 8610 10050 8638
rect 2238 8218 2266 8246
rect 2290 8218 2318 8246
rect 2342 8218 2370 8246
rect 17598 8218 17626 8246
rect 17650 8218 17678 8246
rect 17702 8218 17730 8246
rect 9918 7826 9946 7854
rect 9970 7826 9998 7854
rect 10022 7826 10050 7854
rect 2238 7434 2266 7462
rect 2290 7434 2318 7462
rect 2342 7434 2370 7462
rect 17598 7434 17626 7462
rect 17650 7434 17678 7462
rect 17702 7434 17730 7462
rect 9918 7042 9946 7070
rect 9970 7042 9998 7070
rect 10022 7042 10050 7070
rect 2238 6650 2266 6678
rect 2290 6650 2318 6678
rect 2342 6650 2370 6678
rect 17598 6650 17626 6678
rect 17650 6650 17678 6678
rect 17702 6650 17730 6678
rect 9918 6258 9946 6286
rect 9970 6258 9998 6286
rect 10022 6258 10050 6286
rect 2238 5866 2266 5894
rect 2290 5866 2318 5894
rect 2342 5866 2370 5894
rect 17598 5866 17626 5894
rect 17650 5866 17678 5894
rect 17702 5866 17730 5894
rect 9918 5474 9946 5502
rect 9970 5474 9998 5502
rect 10022 5474 10050 5502
rect 2238 5082 2266 5110
rect 2290 5082 2318 5110
rect 2342 5082 2370 5110
rect 17598 5082 17626 5110
rect 17650 5082 17678 5110
rect 17702 5082 17730 5110
rect 9918 4690 9946 4718
rect 9970 4690 9998 4718
rect 10022 4690 10050 4718
rect 2238 4298 2266 4326
rect 2290 4298 2318 4326
rect 2342 4298 2370 4326
rect 17598 4298 17626 4326
rect 17650 4298 17678 4326
rect 17702 4298 17730 4326
rect 9918 3906 9946 3934
rect 9970 3906 9998 3934
rect 10022 3906 10050 3934
rect 2238 3514 2266 3542
rect 2290 3514 2318 3542
rect 2342 3514 2370 3542
rect 17598 3514 17626 3542
rect 17650 3514 17678 3542
rect 17702 3514 17730 3542
rect 9918 3122 9946 3150
rect 9970 3122 9998 3150
rect 10022 3122 10050 3150
rect 2238 2730 2266 2758
rect 2290 2730 2318 2758
rect 2342 2730 2370 2758
rect 17598 2730 17626 2758
rect 17650 2730 17678 2758
rect 17702 2730 17730 2758
rect 9918 2338 9946 2366
rect 9970 2338 9998 2366
rect 10022 2338 10050 2366
rect 2238 1946 2266 1974
rect 2290 1946 2318 1974
rect 2342 1946 2370 1974
rect 17598 1946 17626 1974
rect 17650 1946 17678 1974
rect 17702 1946 17730 1974
rect 9918 1554 9946 1582
rect 9970 1554 9998 1582
rect 10022 1554 10050 1582
<< metal4 >>
rect 2224 19222 2384 19238
rect 2224 19194 2238 19222
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2370 19194 2384 19222
rect 2224 18438 2384 19194
rect 2224 18410 2238 18438
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2370 18410 2384 18438
rect 2224 17654 2384 18410
rect 2224 17626 2238 17654
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2370 17626 2384 17654
rect 2224 16870 2384 17626
rect 2224 16842 2238 16870
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2370 16842 2384 16870
rect 2224 16086 2384 16842
rect 2224 16058 2238 16086
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2370 16058 2384 16086
rect 2224 15302 2384 16058
rect 2224 15274 2238 15302
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2370 15274 2384 15302
rect 2224 14518 2384 15274
rect 2224 14490 2238 14518
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2370 14490 2384 14518
rect 2224 13734 2384 14490
rect 2224 13706 2238 13734
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2370 13706 2384 13734
rect 2224 12950 2384 13706
rect 2224 12922 2238 12950
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2370 12922 2384 12950
rect 2224 12166 2384 12922
rect 2224 12138 2238 12166
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2370 12138 2384 12166
rect 2224 11382 2384 12138
rect 2224 11354 2238 11382
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2370 11354 2384 11382
rect 2224 10598 2384 11354
rect 2224 10570 2238 10598
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2370 10570 2384 10598
rect 2224 9814 2384 10570
rect 2224 9786 2238 9814
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2370 9786 2384 9814
rect 2224 9030 2384 9786
rect 9904 18830 10064 19238
rect 9904 18802 9918 18830
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 10050 18802 10064 18830
rect 9904 18046 10064 18802
rect 9904 18018 9918 18046
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 10050 18018 10064 18046
rect 9904 17262 10064 18018
rect 9904 17234 9918 17262
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 10050 17234 10064 17262
rect 9904 16478 10064 17234
rect 9904 16450 9918 16478
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 10050 16450 10064 16478
rect 9904 15694 10064 16450
rect 9904 15666 9918 15694
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 10050 15666 10064 15694
rect 9904 14910 10064 15666
rect 9904 14882 9918 14910
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 10050 14882 10064 14910
rect 9904 14126 10064 14882
rect 9904 14098 9918 14126
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 10050 14098 10064 14126
rect 9904 13342 10064 14098
rect 9904 13314 9918 13342
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 10050 13314 10064 13342
rect 9904 12558 10064 13314
rect 9904 12530 9918 12558
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 10050 12530 10064 12558
rect 9904 11774 10064 12530
rect 9904 11746 9918 11774
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 10050 11746 10064 11774
rect 9904 10990 10064 11746
rect 9904 10962 9918 10990
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 10050 10962 10064 10990
rect 9904 10206 10064 10962
rect 9904 10178 9918 10206
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 10050 10178 10064 10206
rect 2224 9002 2238 9030
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2370 9002 2384 9030
rect 2224 8246 2384 9002
rect 8022 9618 8050 9623
rect 8022 8778 8050 9590
rect 8022 8745 8050 8750
rect 9904 9422 10064 10178
rect 9904 9394 9918 9422
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 10050 9394 10064 9422
rect 2224 8218 2238 8246
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2370 8218 2384 8246
rect 2224 7462 2384 8218
rect 2224 7434 2238 7462
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2370 7434 2384 7462
rect 2224 6678 2384 7434
rect 2224 6650 2238 6678
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2370 6650 2384 6678
rect 2224 5894 2384 6650
rect 2224 5866 2238 5894
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2370 5866 2384 5894
rect 2224 5110 2384 5866
rect 2224 5082 2238 5110
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2370 5082 2384 5110
rect 2224 4326 2384 5082
rect 2224 4298 2238 4326
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2370 4298 2384 4326
rect 2224 3542 2384 4298
rect 2224 3514 2238 3542
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2370 3514 2384 3542
rect 2224 2758 2384 3514
rect 2224 2730 2238 2758
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2370 2730 2384 2758
rect 2224 1974 2384 2730
rect 2224 1946 2238 1974
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2370 1946 2384 1974
rect 2224 1538 2384 1946
rect 9904 8638 10064 9394
rect 9904 8610 9918 8638
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 10050 8610 10064 8638
rect 9904 7854 10064 8610
rect 9904 7826 9918 7854
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 10050 7826 10064 7854
rect 9904 7070 10064 7826
rect 9904 7042 9918 7070
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 10050 7042 10064 7070
rect 9904 6286 10064 7042
rect 9904 6258 9918 6286
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 10050 6258 10064 6286
rect 9904 5502 10064 6258
rect 9904 5474 9918 5502
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 10050 5474 10064 5502
rect 9904 4718 10064 5474
rect 9904 4690 9918 4718
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 10050 4690 10064 4718
rect 9904 3934 10064 4690
rect 9904 3906 9918 3934
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 10050 3906 10064 3934
rect 9904 3150 10064 3906
rect 9904 3122 9918 3150
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 10050 3122 10064 3150
rect 9904 2366 10064 3122
rect 9904 2338 9918 2366
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 10050 2338 10064 2366
rect 9904 1582 10064 2338
rect 9904 1554 9918 1582
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 10050 1554 10064 1582
rect 9904 1538 10064 1554
rect 17584 19222 17744 19238
rect 17584 19194 17598 19222
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17730 19194 17744 19222
rect 17584 18438 17744 19194
rect 17584 18410 17598 18438
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17730 18410 17744 18438
rect 17584 17654 17744 18410
rect 17584 17626 17598 17654
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17730 17626 17744 17654
rect 17584 16870 17744 17626
rect 17584 16842 17598 16870
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17730 16842 17744 16870
rect 17584 16086 17744 16842
rect 17584 16058 17598 16086
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17730 16058 17744 16086
rect 17584 15302 17744 16058
rect 17584 15274 17598 15302
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17730 15274 17744 15302
rect 17584 14518 17744 15274
rect 17584 14490 17598 14518
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17730 14490 17744 14518
rect 17584 13734 17744 14490
rect 17584 13706 17598 13734
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17730 13706 17744 13734
rect 17584 12950 17744 13706
rect 17584 12922 17598 12950
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17730 12922 17744 12950
rect 17584 12166 17744 12922
rect 17584 12138 17598 12166
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17730 12138 17744 12166
rect 17584 11382 17744 12138
rect 17584 11354 17598 11382
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17730 11354 17744 11382
rect 17584 10598 17744 11354
rect 17584 10570 17598 10598
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17730 10570 17744 10598
rect 17584 9814 17744 10570
rect 17584 9786 17598 9814
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17730 9786 17744 9814
rect 17584 9030 17744 9786
rect 17584 9002 17598 9030
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17730 9002 17744 9030
rect 17584 8246 17744 9002
rect 17584 8218 17598 8246
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17730 8218 17744 8246
rect 17584 7462 17744 8218
rect 17584 7434 17598 7462
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17730 7434 17744 7462
rect 17584 6678 17744 7434
rect 17584 6650 17598 6678
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17730 6650 17744 6678
rect 17584 5894 17744 6650
rect 17584 5866 17598 5894
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17730 5866 17744 5894
rect 17584 5110 17744 5866
rect 17584 5082 17598 5110
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17730 5082 17744 5110
rect 17584 4326 17744 5082
rect 17584 4298 17598 4326
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17730 4298 17744 4326
rect 17584 3542 17744 4298
rect 17584 3514 17598 3542
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17730 3514 17744 3542
rect 17584 2758 17744 3514
rect 17584 2730 17598 2758
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17730 2730 17744 2758
rect 17584 1974 17744 2730
rect 17584 1946 17598 1974
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17730 1946 17744 1974
rect 17584 1538 17744 1946
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _091_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 7728 0 -1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _092_
timestamp 1698175906
transform 1 0 9576 0 -1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _093_
timestamp 1698175906
transform -1 0 8960 0 -1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _094_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 7224 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _095_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8232 0 1 10192
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _096_
timestamp 1698175906
transform -1 0 8512 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _097_
timestamp 1698175906
transform -1 0 8176 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _098_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8624 0 -1 12544
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _099_
timestamp 1698175906
transform 1 0 6888 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _100_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 7784 0 -1 10976
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _101_
timestamp 1698175906
transform 1 0 6720 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _102_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8064 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _103_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8064 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _104_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8176 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _105_
timestamp 1698175906
transform -1 0 9184 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _106_
timestamp 1698175906
transform -1 0 9464 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _107_
timestamp 1698175906
transform 1 0 7560 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _108_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9016 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _109_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 9800 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _110_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 9184 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _111_
timestamp 1698175906
transform 1 0 8624 0 1 13328
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _112_
timestamp 1698175906
transform 1 0 7952 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _113_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8680 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _114_
timestamp 1698175906
transform 1 0 8904 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _115_
timestamp 1698175906
transform -1 0 7392 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _116_
timestamp 1698175906
transform 1 0 7224 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _117_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 6104 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _118_
timestamp 1698175906
transform -1 0 6104 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _119_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 8680 0 1 7056
box -43 -43 715 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _120_
timestamp 1698175906
transform -1 0 8400 0 1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _121_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 8232 0 1 10192
box -43 -43 771 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _122_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 8512 0 -1 10976
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _123_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 6720 0 -1 10192
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _124_
timestamp 1698175906
transform -1 0 6552 0 1 10976
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _125_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 7224 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _126_
timestamp 1698175906
transform -1 0 7728 0 -1 11760
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _127_
timestamp 1698175906
transform -1 0 7784 0 -1 12544
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _128_
timestamp 1698175906
transform 1 0 6664 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _129_
timestamp 1698175906
transform 1 0 10640 0 1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _130_
timestamp 1698175906
transform 1 0 7560 0 -1 9408
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _131_
timestamp 1698175906
transform 1 0 9688 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _132_
timestamp 1698175906
transform 1 0 13104 0 -1 8624
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _133_
timestamp 1698175906
transform 1 0 12656 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _134_
timestamp 1698175906
transform -1 0 6552 0 1 11760
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _135_
timestamp 1698175906
transform -1 0 7112 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _136_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9184 0 -1 11760
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _137_
timestamp 1698175906
transform 1 0 9744 0 1 12544
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _138_
timestamp 1698175906
transform -1 0 10248 0 1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _139_
timestamp 1698175906
transform -1 0 9632 0 1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _140_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 7224 0 1 10192
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _141_
timestamp 1698175906
transform -1 0 6216 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _142_
timestamp 1698175906
transform 1 0 13384 0 -1 12544
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _143_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 7952 0 1 9408
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _144_
timestamp 1698175906
transform 1 0 10136 0 1 8624
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _145_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9184 0 -1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _146_
timestamp 1698175906
transform 1 0 12040 0 1 10976
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _147_
timestamp 1698175906
transform 1 0 13104 0 -1 12544
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _148_
timestamp 1698175906
transform -1 0 9072 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _149_
timestamp 1698175906
transform 1 0 8064 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _150_
timestamp 1698175906
transform -1 0 11928 0 1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _151_
timestamp 1698175906
transform -1 0 11536 0 1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _152_
timestamp 1698175906
transform -1 0 11032 0 1 7056
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _153_
timestamp 1698175906
transform 1 0 9016 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _154_
timestamp 1698175906
transform 1 0 11592 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _155_
timestamp 1698175906
transform -1 0 10192 0 1 7840
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _156_
timestamp 1698175906
transform 1 0 10192 0 1 7840
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _157_
timestamp 1698175906
transform 1 0 12544 0 -1 7840
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _158_
timestamp 1698175906
transform -1 0 13272 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _159_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 8960 0 1 9408
box -43 -43 1051 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _160_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9464 0 1 10192
box -43 -43 883 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _161_
timestamp 1698175906
transform 1 0 13496 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _162_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 12544 0 1 9408
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _163_
timestamp 1698175906
transform -1 0 10136 0 1 9408
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _164_
timestamp 1698175906
transform 1 0 11144 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _165_
timestamp 1698175906
transform 1 0 10136 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _166_
timestamp 1698175906
transform 1 0 11088 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _167_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 11984 0 -1 12544
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _168_
timestamp 1698175906
transform -1 0 11592 0 1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _169_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10584 0 1 11760
box -43 -43 715 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _170_
timestamp 1698175906
transform -1 0 10920 0 -1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _171_
timestamp 1698175906
transform 1 0 8008 0 -1 10192
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _172_
timestamp 1698175906
transform 1 0 13160 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _173_
timestamp 1698175906
transform 1 0 12432 0 1 10976
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _174_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10024 0 -1 9408
box -43 -43 659 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _175_
timestamp 1698175906
transform 1 0 10640 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _176_
timestamp 1698175906
transform -1 0 13328 0 1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _177_
timestamp 1698175906
transform -1 0 13048 0 -1 12544
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _178_
timestamp 1698175906
transform -1 0 7672 0 1 8624
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _179_
timestamp 1698175906
transform -1 0 7392 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _180_
timestamp 1698175906
transform 1 0 11984 0 1 8624
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _181_
timestamp 1698175906
transform -1 0 12320 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _182_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 7728 0 1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _183_
timestamp 1698175906
transform -1 0 6552 0 1 7840
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _184_
timestamp 1698175906
transform -1 0 10584 0 -1 7840
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _185_
timestamp 1698175906
transform 1 0 6888 0 -1 7840
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _186_
timestamp 1698175906
transform -1 0 6608 0 -1 10976
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _187_
timestamp 1698175906
transform 1 0 5880 0 -1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _188_
timestamp 1698175906
transform 1 0 12544 0 1 8624
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _189_
timestamp 1698175906
transform -1 0 6552 0 1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _190_
timestamp 1698175906
transform 1 0 8904 0 -1 14112
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _191_
timestamp 1698175906
transform -1 0 6384 0 1 10192
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _192_
timestamp 1698175906
transform 1 0 12488 0 1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _193_
timestamp 1698175906
transform 1 0 7000 0 1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _194_
timestamp 1698175906
transform 1 0 10696 0 -1 14112
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _195_
timestamp 1698175906
transform 1 0 9744 0 -1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _196_
timestamp 1698175906
transform 1 0 11872 0 1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _197_
timestamp 1698175906
transform 1 0 12544 0 -1 10192
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _198_
timestamp 1698175906
transform 1 0 10752 0 1 9408
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _199_
timestamp 1698175906
transform 1 0 10640 0 1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _200_
timestamp 1698175906
transform -1 0 11424 0 -1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _201_
timestamp 1698175906
transform 1 0 12544 0 -1 10976
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _202_
timestamp 1698175906
transform -1 0 11536 0 -1 8624
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _203_
timestamp 1698175906
transform 1 0 12544 0 -1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _204_
timestamp 1698175906
transform -1 0 7336 0 -1 8624
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _205_
timestamp 1698175906
transform 1 0 11592 0 1 7840
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _209_
timestamp 1698175906
transform 1 0 13664 0 1 13328
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _210_
timestamp 1698175906
transform -1 0 6608 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _211_
timestamp 1698175906
transform 1 0 14168 0 -1 13328
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__182__CLK dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9464 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__183__CLK
timestamp 1698175906
transform 1 0 6776 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__184__CLK
timestamp 1698175906
transform 1 0 10696 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__185__CLK
timestamp 1698175906
transform 1 0 8736 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__186__CLK
timestamp 1698175906
transform 1 0 6608 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__187__CLK
timestamp 1698175906
transform 1 0 7896 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__188__CLK
timestamp 1698175906
transform 1 0 14280 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__189__CLK
timestamp 1698175906
transform 1 0 6552 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__190__CLK
timestamp 1698175906
transform -1 0 8904 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__191__CLK
timestamp 1698175906
transform 1 0 6328 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__192__CLK
timestamp 1698175906
transform 1 0 14224 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__193__CLK
timestamp 1698175906
transform 1 0 9072 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__194__CLK
timestamp 1698175906
transform -1 0 12768 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__195__CLK
timestamp 1698175906
transform 1 0 11480 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__196__CLK
timestamp 1698175906
transform 1 0 13608 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__197__CLK
timestamp 1698175906
transform 1 0 14280 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__198__CLK
timestamp 1698175906
transform 1 0 13216 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__199__CLK
timestamp 1698175906
transform 1 0 12376 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__200__CLK
timestamp 1698175906
transform 1 0 11704 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__201__CLK
timestamp 1698175906
transform 1 0 14280 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__202__CLK
timestamp 1698175906
transform 1 0 11648 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__203__CLK
timestamp 1698175906
transform 1 0 14616 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__204__CLK
timestamp 1698175906
transform 1 0 7448 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__205__CLK
timestamp 1698175906
transform 1 0 13328 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1698175906
transform 1 0 8792 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8904 0 -1 10976
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1698175906
transform -1 0 10192 0 1 10976
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1698175906
transform 1 0 10752 0 1 10192
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 784 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_36 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 2688 0 1 1568
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_52 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 3584 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_54 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 3696 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_59 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 3976 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_67
timestamp 1698175906
transform 1 0 4424 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698175906
transform 1 0 4592 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698175906
transform 1 0 6496 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_138
timestamp 1698175906
transform 1 0 8400 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_172 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10304 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_176
timestamp 1698175906
transform 1 0 10528 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_206
timestamp 1698175906
transform 1 0 12208 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_210
timestamp 1698175906
transform 1 0 12432 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_240
timestamp 1698175906
transform 1 0 14112 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_274
timestamp 1698175906
transform 1 0 16016 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_308
timestamp 1698175906
transform 1 0 17920 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_342
timestamp 1698175906
transform 1 0 19824 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_346
timestamp 1698175906
transform 1 0 20048 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_348
timestamp 1698175906
transform 1 0 20160 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 784 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698175906
transform 1 0 4368 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698175906
transform 1 0 4704 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698175906
transform 1 0 8288 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_142
timestamp 1698175906
transform 1 0 8624 0 -1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_174
timestamp 1698175906
transform 1 0 10416 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_178
timestamp 1698175906
transform 1 0 10640 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_180
timestamp 1698175906
transform 1 0 10752 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_207
timestamp 1698175906
transform 1 0 12264 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_209
timestamp 1698175906
transform 1 0 12376 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_212
timestamp 1698175906
transform 1 0 12544 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_276
timestamp 1698175906
transform 1 0 16128 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_282
timestamp 1698175906
transform 1 0 16464 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_346
timestamp 1698175906
transform 1 0 20048 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_348
timestamp 1698175906
transform 1 0 20160 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698175906
transform 1 0 784 0 1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698175906
transform 1 0 2576 0 1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698175906
transform 1 0 2744 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698175906
transform 1 0 6328 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_107
timestamp 1698175906
transform 1 0 6664 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_171
timestamp 1698175906
transform 1 0 10248 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_177
timestamp 1698175906
transform 1 0 10584 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_241
timestamp 1698175906
transform 1 0 14168 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698175906
transform 1 0 14504 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698175906
transform 1 0 18088 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_317
timestamp 1698175906
transform 1 0 18424 0 1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698175906
transform 1 0 784 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698175906
transform 1 0 4368 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698175906
transform 1 0 4704 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698175906
transform 1 0 8288 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_142
timestamp 1698175906
transform 1 0 8624 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_206
timestamp 1698175906
transform 1 0 12208 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_212
timestamp 1698175906
transform 1 0 12544 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_276
timestamp 1698175906
transform 1 0 16128 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_282
timestamp 1698175906
transform 1 0 16464 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_346
timestamp 1698175906
transform 1 0 20048 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_348
timestamp 1698175906
transform 1 0 20160 0 -1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698175906
transform 1 0 784 0 1 3136
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698175906
transform 1 0 2576 0 1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698175906
transform 1 0 2744 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698175906
transform 1 0 6328 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_107
timestamp 1698175906
transform 1 0 6664 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698175906
transform 1 0 10248 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_177
timestamp 1698175906
transform 1 0 10584 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_241
timestamp 1698175906
transform 1 0 14168 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698175906
transform 1 0 14504 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698175906
transform 1 0 18088 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_317
timestamp 1698175906
transform 1 0 18424 0 1 3136
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698175906
transform 1 0 784 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698175906
transform 1 0 4368 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698175906
transform 1 0 4704 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698175906
transform 1 0 8288 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_142
timestamp 1698175906
transform 1 0 8624 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_206
timestamp 1698175906
transform 1 0 12208 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_212
timestamp 1698175906
transform 1 0 12544 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698175906
transform 1 0 16128 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_282
timestamp 1698175906
transform 1 0 16464 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_346
timestamp 1698175906
transform 1 0 20048 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_348
timestamp 1698175906
transform 1 0 20160 0 -1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698175906
transform 1 0 784 0 1 3920
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698175906
transform 1 0 2576 0 1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698175906
transform 1 0 2744 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698175906
transform 1 0 6328 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_107
timestamp 1698175906
transform 1 0 6664 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_171
timestamp 1698175906
transform 1 0 10248 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_177
timestamp 1698175906
transform 1 0 10584 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_241
timestamp 1698175906
transform 1 0 14168 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_247
timestamp 1698175906
transform 1 0 14504 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_311
timestamp 1698175906
transform 1 0 18088 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_317
timestamp 1698175906
transform 1 0 18424 0 1 3920
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698175906
transform 1 0 784 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698175906
transform 1 0 4368 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_72
timestamp 1698175906
transform 1 0 4704 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698175906
transform 1 0 8288 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_142
timestamp 1698175906
transform 1 0 8624 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_206
timestamp 1698175906
transform 1 0 12208 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_212
timestamp 1698175906
transform 1 0 12544 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_276
timestamp 1698175906
transform 1 0 16128 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_282
timestamp 1698175906
transform 1 0 16464 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_346
timestamp 1698175906
transform 1 0 20048 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_348
timestamp 1698175906
transform 1 0 20160 0 -1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698175906
transform 1 0 784 0 1 4704
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698175906
transform 1 0 2576 0 1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_37
timestamp 1698175906
transform 1 0 2744 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_101
timestamp 1698175906
transform 1 0 6328 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_107
timestamp 1698175906
transform 1 0 6664 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_171
timestamp 1698175906
transform 1 0 10248 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_177
timestamp 1698175906
transform 1 0 10584 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_241
timestamp 1698175906
transform 1 0 14168 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_247
timestamp 1698175906
transform 1 0 14504 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_311
timestamp 1698175906
transform 1 0 18088 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_317
timestamp 1698175906
transform 1 0 18424 0 1 4704
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698175906
transform 1 0 784 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698175906
transform 1 0 4368 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_72
timestamp 1698175906
transform 1 0 4704 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_136
timestamp 1698175906
transform 1 0 8288 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_142
timestamp 1698175906
transform 1 0 8624 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_206
timestamp 1698175906
transform 1 0 12208 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_212
timestamp 1698175906
transform 1 0 12544 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_276
timestamp 1698175906
transform 1 0 16128 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_282
timestamp 1698175906
transform 1 0 16464 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_346
timestamp 1698175906
transform 1 0 20048 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_348
timestamp 1698175906
transform 1 0 20160 0 -1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698175906
transform 1 0 784 0 1 5488
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698175906
transform 1 0 2576 0 1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_37
timestamp 1698175906
transform 1 0 2744 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698175906
transform 1 0 6328 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_107
timestamp 1698175906
transform 1 0 6664 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_171
timestamp 1698175906
transform 1 0 10248 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_177
timestamp 1698175906
transform 1 0 10584 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_241
timestamp 1698175906
transform 1 0 14168 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_247
timestamp 1698175906
transform 1 0 14504 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_311
timestamp 1698175906
transform 1 0 18088 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_317
timestamp 1698175906
transform 1 0 18424 0 1 5488
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2
timestamp 1698175906
transform 1 0 784 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698175906
transform 1 0 4368 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_72
timestamp 1698175906
transform 1 0 4704 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698175906
transform 1 0 8288 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_142
timestamp 1698175906
transform 1 0 8624 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_206
timestamp 1698175906
transform 1 0 12208 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_212
timestamp 1698175906
transform 1 0 12544 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_276
timestamp 1698175906
transform 1 0 16128 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_282
timestamp 1698175906
transform 1 0 16464 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_346
timestamp 1698175906
transform 1 0 20048 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_348
timestamp 1698175906
transform 1 0 20160 0 -1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698175906
transform 1 0 784 0 1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698175906
transform 1 0 2576 0 1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_37
timestamp 1698175906
transform 1 0 2744 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698175906
transform 1 0 6328 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_107
timestamp 1698175906
transform 1 0 6664 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_171
timestamp 1698175906
transform 1 0 10248 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_177
timestamp 1698175906
transform 1 0 10584 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_241
timestamp 1698175906
transform 1 0 14168 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_247
timestamp 1698175906
transform 1 0 14504 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_311
timestamp 1698175906
transform 1 0 18088 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_317
timestamp 1698175906
transform 1 0 18424 0 1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_2
timestamp 1698175906
transform 1 0 784 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_66
timestamp 1698175906
transform 1 0 4368 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_72
timestamp 1698175906
transform 1 0 4704 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_136
timestamp 1698175906
transform 1 0 8288 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_142
timestamp 1698175906
transform 1 0 8624 0 -1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_158
timestamp 1698175906
transform 1 0 9520 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_191
timestamp 1698175906
transform 1 0 11368 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_195
timestamp 1698175906
transform 1 0 11592 0 -1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_203
timestamp 1698175906
transform 1 0 12040 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_207
timestamp 1698175906
transform 1 0 12264 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_209
timestamp 1698175906
transform 1 0 12376 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_212
timestamp 1698175906
transform 1 0 12544 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_276
timestamp 1698175906
transform 1 0 16128 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_282
timestamp 1698175906
transform 1 0 16464 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_346
timestamp 1698175906
transform 1 0 20048 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_348
timestamp 1698175906
transform 1 0 20160 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698175906
transform 1 0 784 0 1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698175906
transform 1 0 2576 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_37
timestamp 1698175906
transform 1 0 2744 0 1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_101
timestamp 1698175906
transform 1 0 6328 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_107
timestamp 1698175906
transform 1 0 6664 0 1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_123
timestamp 1698175906
transform 1 0 7560 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_143
timestamp 1698175906
transform 1 0 8680 0 1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_177
timestamp 1698175906
transform 1 0 10584 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_179
timestamp 1698175906
transform 1 0 10696 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_185
timestamp 1698175906
transform 1 0 11032 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_193
timestamp 1698175906
transform 1 0 11480 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_197
timestamp 1698175906
transform 1 0 11704 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_199
timestamp 1698175906
transform 1 0 11816 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_229
timestamp 1698175906
transform 1 0 13496 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_233
timestamp 1698175906
transform 1 0 13720 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_241
timestamp 1698175906
transform 1 0 14168 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_247
timestamp 1698175906
transform 1 0 14504 0 1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_311
timestamp 1698175906
transform 1 0 18088 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_317
timestamp 1698175906
transform 1 0 18424 0 1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_2
timestamp 1698175906
transform 1 0 784 0 -1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_66
timestamp 1698175906
transform 1 0 4368 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_72
timestamp 1698175906
transform 1 0 4704 0 -1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_104
timestamp 1698175906
transform 1 0 6496 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_108
timestamp 1698175906
transform 1 0 6720 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_110
timestamp 1698175906
transform 1 0 6832 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_142
timestamp 1698175906
transform 1 0 8624 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_146
timestamp 1698175906
transform 1 0 8848 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_177
timestamp 1698175906
transform 1 0 10584 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_181
timestamp 1698175906
transform 1 0 10808 0 -1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_197
timestamp 1698175906
transform 1 0 11704 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_205
timestamp 1698175906
transform 1 0 12152 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_209
timestamp 1698175906
transform 1 0 12376 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_225
timestamp 1698175906
transform 1 0 13272 0 -1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_257
timestamp 1698175906
transform 1 0 15064 0 -1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_273
timestamp 1698175906
transform 1 0 15960 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_277
timestamp 1698175906
transform 1 0 16184 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_279
timestamp 1698175906
transform 1 0 16296 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_282
timestamp 1698175906
transform 1 0 16464 0 -1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_346
timestamp 1698175906
transform 1 0 20048 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_348
timestamp 1698175906
transform 1 0 20160 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_2
timestamp 1698175906
transform 1 0 784 0 1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698175906
transform 1 0 2576 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_37
timestamp 1698175906
transform 1 0 2744 0 1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_69
timestamp 1698175906
transform 1 0 4536 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_73
timestamp 1698175906
transform 1 0 4760 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_75
timestamp 1698175906
transform 1 0 4872 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_107
timestamp 1698175906
transform 1 0 6664 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_111
timestamp 1698175906
transform 1 0 6888 0 1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_127
timestamp 1698175906
transform 1 0 7784 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_131
timestamp 1698175906
transform 1 0 8008 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_138
timestamp 1698175906
transform 1 0 8400 0 1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_154
timestamp 1698175906
transform 1 0 9296 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_162
timestamp 1698175906
transform 1 0 9744 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_164
timestamp 1698175906
transform 1 0 9856 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_177
timestamp 1698175906
transform 1 0 10584 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_184
timestamp 1698175906
transform 1 0 10976 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_192
timestamp 1698175906
transform 1 0 11424 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_194
timestamp 1698175906
transform 1 0 11536 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_224
timestamp 1698175906
transform 1 0 13216 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_228
timestamp 1698175906
transform 1 0 13440 0 1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_244
timestamp 1698175906
transform 1 0 14336 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_247
timestamp 1698175906
transform 1 0 14504 0 1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_311
timestamp 1698175906
transform 1 0 18088 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_317
timestamp 1698175906
transform 1 0 18424 0 1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_28
timestamp 1698175906
transform 1 0 2240 0 -1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_60
timestamp 1698175906
transform 1 0 4032 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_68
timestamp 1698175906
transform 1 0 4480 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_72
timestamp 1698175906
transform 1 0 4704 0 -1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_88
timestamp 1698175906
transform 1 0 5600 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_119
timestamp 1698175906
transform 1 0 7336 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_123
timestamp 1698175906
transform 1 0 7560 0 -1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_139
timestamp 1698175906
transform 1 0 8456 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_148
timestamp 1698175906
transform 1 0 8960 0 -1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_164
timestamp 1698175906
transform 1 0 9856 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_194
timestamp 1698175906
transform 1 0 11536 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_198
timestamp 1698175906
transform 1 0 11760 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_202
timestamp 1698175906
transform 1 0 11984 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_208
timestamp 1698175906
transform 1 0 12320 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_212
timestamp 1698175906
transform 1 0 12544 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_220
timestamp 1698175906
transform 1 0 12992 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_227
timestamp 1698175906
transform 1 0 13384 0 -1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_259
timestamp 1698175906
transform 1 0 15176 0 -1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_275
timestamp 1698175906
transform 1 0 16072 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_279
timestamp 1698175906
transform 1 0 16296 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_282
timestamp 1698175906
transform 1 0 16464 0 -1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_314
timestamp 1698175906
transform 1 0 18256 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_322
timestamp 1698175906
transform 1 0 18704 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_28
timestamp 1698175906
transform 1 0 2240 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_32
timestamp 1698175906
transform 1 0 2464 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698175906
transform 1 0 2576 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_37
timestamp 1698175906
transform 1 0 2744 0 1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_69
timestamp 1698175906
transform 1 0 4536 0 1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_85
timestamp 1698175906
transform 1 0 5432 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_89
timestamp 1698175906
transform 1 0 5656 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_107
timestamp 1698175906
transform 1 0 6664 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_111
timestamp 1698175906
transform 1 0 6888 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_125
timestamp 1698175906
transform 1 0 7672 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_129
timestamp 1698175906
transform 1 0 7896 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_140
timestamp 1698175906
transform 1 0 8512 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_142
timestamp 1698175906
transform 1 0 8624 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_157
timestamp 1698175906
transform 1 0 9464 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_167
timestamp 1698175906
transform 1 0 10024 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_174
timestamp 1698175906
transform 1 0 10416 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_177
timestamp 1698175906
transform 1 0 10584 0 1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_193
timestamp 1698175906
transform 1 0 11480 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_201
timestamp 1698175906
transform 1 0 11928 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_211
timestamp 1698175906
transform 1 0 12488 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_241
timestamp 1698175906
transform 1 0 14168 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_247
timestamp 1698175906
transform 1 0 14504 0 1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_311
timestamp 1698175906
transform 1 0 18088 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_317
timestamp 1698175906
transform 1 0 18424 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_321
timestamp 1698175906
transform 1 0 18648 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_28
timestamp 1698175906
transform 1 0 2240 0 -1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_60
timestamp 1698175906
transform 1 0 4032 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_68
timestamp 1698175906
transform 1 0 4480 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_72
timestamp 1698175906
transform 1 0 4704 0 -1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_88
timestamp 1698175906
transform 1 0 5600 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_96
timestamp 1698175906
transform 1 0 6048 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_106
timestamp 1698175906
transform 1 0 6608 0 -1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_122
timestamp 1698175906
transform 1 0 7504 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_142
timestamp 1698175906
transform 1 0 8624 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_146
timestamp 1698175906
transform 1 0 8848 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_163
timestamp 1698175906
transform 1 0 9800 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_184
timestamp 1698175906
transform 1 0 10976 0 -1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_200
timestamp 1698175906
transform 1 0 11872 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_208
timestamp 1698175906
transform 1 0 12320 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_212
timestamp 1698175906
transform 1 0 12544 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_222
timestamp 1698175906
transform 1 0 13104 0 -1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_254
timestamp 1698175906
transform 1 0 14896 0 -1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_270
timestamp 1698175906
transform 1 0 15792 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_278
timestamp 1698175906
transform 1 0 16240 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_282
timestamp 1698175906
transform 1 0 16464 0 -1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_346
timestamp 1698175906
transform 1 0 20048 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_348
timestamp 1698175906
transform 1 0 20160 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_2
timestamp 1698175906
transform 1 0 784 0 1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698175906
transform 1 0 2576 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_37
timestamp 1698175906
transform 1 0 2744 0 1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_101
timestamp 1698175906
transform 1 0 6328 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_107
timestamp 1698175906
transform 1 0 6664 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_115
timestamp 1698175906
transform 1 0 7112 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_119
timestamp 1698175906
transform 1 0 7336 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_148
timestamp 1698175906
transform 1 0 8960 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_177
timestamp 1698175906
transform 1 0 10584 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_179
timestamp 1698175906
transform 1 0 10696 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_209
timestamp 1698175906
transform 1 0 12376 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_211
timestamp 1698175906
transform 1 0 12488 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_222
timestamp 1698175906
transform 1 0 13104 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_226
timestamp 1698175906
transform 1 0 13328 0 1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_242
timestamp 1698175906
transform 1 0 14224 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_244
timestamp 1698175906
transform 1 0 14336 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_247
timestamp 1698175906
transform 1 0 14504 0 1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_311
timestamp 1698175906
transform 1 0 18088 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_317
timestamp 1698175906
transform 1 0 18424 0 1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_2
timestamp 1698175906
transform 1 0 784 0 -1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_66
timestamp 1698175906
transform 1 0 4368 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_72
timestamp 1698175906
transform 1 0 4704 0 -1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_88
timestamp 1698175906
transform 1 0 5600 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_92
timestamp 1698175906
transform 1 0 5824 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_99
timestamp 1698175906
transform 1 0 6216 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_108
timestamp 1698175906
transform 1 0 6720 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_110
timestamp 1698175906
transform 1 0 6832 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_142
timestamp 1698175906
transform 1 0 8624 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_184
timestamp 1698175906
transform 1 0 10976 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_186
timestamp 1698175906
transform 1 0 11088 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_201
timestamp 1698175906
transform 1 0 11928 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_209
timestamp 1698175906
transform 1 0 12376 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_241
timestamp 1698175906
transform 1 0 14168 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_245
timestamp 1698175906
transform 1 0 14392 0 -1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_277
timestamp 1698175906
transform 1 0 16184 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_279
timestamp 1698175906
transform 1 0 16296 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_282
timestamp 1698175906
transform 1 0 16464 0 -1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_346
timestamp 1698175906
transform 1 0 20048 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_348
timestamp 1698175906
transform 1 0 20160 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_2
timestamp 1698175906
transform 1 0 784 0 1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698175906
transform 1 0 2576 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_37
timestamp 1698175906
transform 1 0 2744 0 1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_69
timestamp 1698175906
transform 1 0 4536 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_102
timestamp 1698175906
transform 1 0 6384 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_104
timestamp 1698175906
transform 1 0 6496 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_121
timestamp 1698175906
transform 1 0 7448 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_172
timestamp 1698175906
transform 1 0 10304 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_174
timestamp 1698175906
transform 1 0 10416 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_177
timestamp 1698175906
transform 1 0 10584 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_179
timestamp 1698175906
transform 1 0 10696 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_230
timestamp 1698175906
transform 1 0 13552 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_238
timestamp 1698175906
transform 1 0 14000 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_242
timestamp 1698175906
transform 1 0 14224 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_244
timestamp 1698175906
transform 1 0 14336 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_247
timestamp 1698175906
transform 1 0 14504 0 1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_311
timestamp 1698175906
transform 1 0 18088 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_317
timestamp 1698175906
transform 1 0 18424 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_321
timestamp 1698175906
transform 1 0 18648 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_28
timestamp 1698175906
transform 1 0 2240 0 -1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_60
timestamp 1698175906
transform 1 0 4032 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_68
timestamp 1698175906
transform 1 0 4480 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_72
timestamp 1698175906
transform 1 0 4704 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_76
timestamp 1698175906
transform 1 0 4928 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_106
timestamp 1698175906
transform 1 0 6608 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_108
timestamp 1698175906
transform 1 0 6720 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_127
timestamp 1698175906
transform 1 0 7784 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_142
timestamp 1698175906
transform 1 0 8624 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_144
timestamp 1698175906
transform 1 0 8736 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_197
timestamp 1698175906
transform 1 0 11704 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_205
timestamp 1698175906
transform 1 0 12152 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_209
timestamp 1698175906
transform 1 0 12376 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_241
timestamp 1698175906
transform 1 0 14168 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_245
timestamp 1698175906
transform 1 0 14392 0 -1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_277
timestamp 1698175906
transform 1 0 16184 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_279
timestamp 1698175906
transform 1 0 16296 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_282
timestamp 1698175906
transform 1 0 16464 0 -1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_314
timestamp 1698175906
transform 1 0 18256 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_322
timestamp 1698175906
transform 1 0 18704 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_2
timestamp 1698175906
transform 1 0 784 0 1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698175906
transform 1 0 2576 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_37
timestamp 1698175906
transform 1 0 2744 0 1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_69
timestamp 1698175906
transform 1 0 4536 0 1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_85
timestamp 1698175906
transform 1 0 5432 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_93
timestamp 1698175906
transform 1 0 5880 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_97
timestamp 1698175906
transform 1 0 6104 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_99
timestamp 1698175906
transform 1 0 6216 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_107
timestamp 1698175906
transform 1 0 6664 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_170
timestamp 1698175906
transform 1 0 10192 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_174
timestamp 1698175906
transform 1 0 10416 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_177
timestamp 1698175906
transform 1 0 10584 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_185
timestamp 1698175906
transform 1 0 11032 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_194
timestamp 1698175906
transform 1 0 11536 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_202
timestamp 1698175906
transform 1 0 11984 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_220
timestamp 1698175906
transform 1 0 12992 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_222
timestamp 1698175906
transform 1 0 13104 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_235
timestamp 1698175906
transform 1 0 13832 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_243
timestamp 1698175906
transform 1 0 14280 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_247
timestamp 1698175906
transform 1 0 14504 0 1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_311
timestamp 1698175906
transform 1 0 18088 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_317
timestamp 1698175906
transform 1 0 18424 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_321
timestamp 1698175906
transform 1 0 18648 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_2
timestamp 1698175906
transform 1 0 784 0 -1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_66
timestamp 1698175906
transform 1 0 4368 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_72
timestamp 1698175906
transform 1 0 4704 0 -1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_104
timestamp 1698175906
transform 1 0 6496 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_108
timestamp 1698175906
transform 1 0 6720 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_116
timestamp 1698175906
transform 1 0 7168 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_120
timestamp 1698175906
transform 1 0 7392 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_142
timestamp 1698175906
transform 1 0 8624 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_165
timestamp 1698175906
transform 1 0 9912 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_173
timestamp 1698175906
transform 1 0 10360 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_183
timestamp 1698175906
transform 1 0 10920 0 -1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_199
timestamp 1698175906
transform 1 0 11816 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_207
timestamp 1698175906
transform 1 0 12264 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_209
timestamp 1698175906
transform 1 0 12376 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_212
timestamp 1698175906
transform 1 0 12544 0 -1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_276
timestamp 1698175906
transform 1 0 16128 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_282
timestamp 1698175906
transform 1 0 16464 0 -1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_346
timestamp 1698175906
transform 1 0 20048 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_348
timestamp 1698175906
transform 1 0 20160 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_2
timestamp 1698175906
transform 1 0 784 0 1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698175906
transform 1 0 2576 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_37
timestamp 1698175906
transform 1 0 2744 0 1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_69
timestamp 1698175906
transform 1 0 4536 0 1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_85
timestamp 1698175906
transform 1 0 5432 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_93
timestamp 1698175906
transform 1 0 5880 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_97
timestamp 1698175906
transform 1 0 6104 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_99
timestamp 1698175906
transform 1 0 6216 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_115
timestamp 1698175906
transform 1 0 7112 0 1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_131
timestamp 1698175906
transform 1 0 8008 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_136
timestamp 1698175906
transform 1 0 8288 0 1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_168
timestamp 1698175906
transform 1 0 10080 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_172
timestamp 1698175906
transform 1 0 10304 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_174
timestamp 1698175906
transform 1 0 10416 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_195
timestamp 1698175906
transform 1 0 11592 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_199
timestamp 1698175906
transform 1 0 11816 0 1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_231
timestamp 1698175906
transform 1 0 13608 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_239
timestamp 1698175906
transform 1 0 14056 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_243
timestamp 1698175906
transform 1 0 14280 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_247
timestamp 1698175906
transform 1 0 14504 0 1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_311
timestamp 1698175906
transform 1 0 18088 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_317
timestamp 1698175906
transform 1 0 18424 0 1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_2
timestamp 1698175906
transform 1 0 784 0 -1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_66
timestamp 1698175906
transform 1 0 4368 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_72
timestamp 1698175906
transform 1 0 4704 0 -1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_88
timestamp 1698175906
transform 1 0 5600 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_92
timestamp 1698175906
transform 1 0 5824 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_127
timestamp 1698175906
transform 1 0 7784 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_131
timestamp 1698175906
transform 1 0 8008 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_139
timestamp 1698175906
transform 1 0 8456 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_151
timestamp 1698175906
transform 1 0 9128 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_159
timestamp 1698175906
transform 1 0 9576 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_202
timestamp 1698175906
transform 1 0 11984 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_212
timestamp 1698175906
transform 1 0 12544 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_221
timestamp 1698175906
transform 1 0 13048 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_232
timestamp 1698175906
transform 1 0 13664 0 -1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_264
timestamp 1698175906
transform 1 0 15456 0 -1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_282
timestamp 1698175906
transform 1 0 16464 0 -1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_346
timestamp 1698175906
transform 1 0 20048 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_348
timestamp 1698175906
transform 1 0 20160 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_28
timestamp 1698175906
transform 1 0 2240 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_32
timestamp 1698175906
transform 1 0 2464 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698175906
transform 1 0 2576 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_37
timestamp 1698175906
transform 1 0 2744 0 1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_69
timestamp 1698175906
transform 1 0 4536 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_73
timestamp 1698175906
transform 1 0 4760 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_75
timestamp 1698175906
transform 1 0 4872 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_115
timestamp 1698175906
transform 1 0 7112 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_123
timestamp 1698175906
transform 1 0 7560 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_125
timestamp 1698175906
transform 1 0 7672 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_155
timestamp 1698175906
transform 1 0 9352 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_159
timestamp 1698175906
transform 1 0 9576 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_161
timestamp 1698175906
transform 1 0 9688 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_168
timestamp 1698175906
transform 1 0 10080 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_172
timestamp 1698175906
transform 1 0 10304 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_174
timestamp 1698175906
transform 1 0 10416 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_177
timestamp 1698175906
transform 1 0 10584 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_207
timestamp 1698175906
transform 1 0 12264 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_240
timestamp 1698175906
transform 1 0 14112 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_244
timestamp 1698175906
transform 1 0 14336 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_247
timestamp 1698175906
transform 1 0 14504 0 1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_311
timestamp 1698175906
transform 1 0 18088 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_317
timestamp 1698175906
transform 1 0 18424 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_321
timestamp 1698175906
transform 1 0 18648 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_2
timestamp 1698175906
transform 1 0 784 0 -1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_66
timestamp 1698175906
transform 1 0 4368 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_72
timestamp 1698175906
transform 1 0 4704 0 -1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_104
timestamp 1698175906
transform 1 0 6496 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_107
timestamp 1698175906
transform 1 0 6664 0 -1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_123
timestamp 1698175906
transform 1 0 7560 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_131
timestamp 1698175906
transform 1 0 8008 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_150
timestamp 1698175906
transform 1 0 9072 0 -1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_182
timestamp 1698175906
transform 1 0 10864 0 -1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_198
timestamp 1698175906
transform 1 0 11760 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_206
timestamp 1698175906
transform 1 0 12208 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_247
timestamp 1698175906
transform 1 0 14504 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_251
timestamp 1698175906
transform 1 0 14728 0 -1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_267
timestamp 1698175906
transform 1 0 15624 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_275
timestamp 1698175906
transform 1 0 16072 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_279
timestamp 1698175906
transform 1 0 16296 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_282
timestamp 1698175906
transform 1 0 16464 0 -1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_314
timestamp 1698175906
transform 1 0 18256 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_322
timestamp 1698175906
transform 1 0 18704 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_2
timestamp 1698175906
transform 1 0 784 0 1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698175906
transform 1 0 2576 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_37
timestamp 1698175906
transform 1 0 2744 0 1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_101
timestamp 1698175906
transform 1 0 6328 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_107
timestamp 1698175906
transform 1 0 6664 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_111
timestamp 1698175906
transform 1 0 6888 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_148
timestamp 1698175906
transform 1 0 8960 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_152
timestamp 1698175906
transform 1 0 9184 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_154
timestamp 1698175906
transform 1 0 9296 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_160
timestamp 1698175906
transform 1 0 9632 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_164
timestamp 1698175906
transform 1 0 9856 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_171
timestamp 1698175906
transform 1 0 10248 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_177
timestamp 1698175906
transform 1 0 10584 0 1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_185
timestamp 1698175906
transform 1 0 11032 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_194
timestamp 1698175906
transform 1 0 11536 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_201
timestamp 1698175906
transform 1 0 11928 0 1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_217
timestamp 1698175906
transform 1 0 12824 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_226
timestamp 1698175906
transform 1 0 13328 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_230
timestamp 1698175906
transform 1 0 13552 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_238
timestamp 1698175906
transform 1 0 14000 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_242
timestamp 1698175906
transform 1 0 14224 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_244
timestamp 1698175906
transform 1 0 14336 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_247
timestamp 1698175906
transform 1 0 14504 0 1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_311
timestamp 1698175906
transform 1 0 18088 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_317
timestamp 1698175906
transform 1 0 18424 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_321
timestamp 1698175906
transform 1 0 18648 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_2
timestamp 1698175906
transform 1 0 784 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_66
timestamp 1698175906
transform 1 0 4368 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_72
timestamp 1698175906
transform 1 0 4704 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_136
timestamp 1698175906
transform 1 0 8288 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_142
timestamp 1698175906
transform 1 0 8624 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_144
timestamp 1698175906
transform 1 0 8736 0 -1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_176
timestamp 1698175906
transform 1 0 10528 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_178
timestamp 1698175906
transform 1 0 10640 0 -1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_208
timestamp 1698175906
transform 1 0 12320 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_212
timestamp 1698175906
transform 1 0 12544 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_216
timestamp 1698175906
transform 1 0 12768 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_282
timestamp 1698175906
transform 1 0 16464 0 -1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_314
timestamp 1698175906
transform 1 0 18256 0 -1 14112
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_322
timestamp 1698175906
transform 1 0 18704 0 -1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_2
timestamp 1698175906
transform 1 0 784 0 1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698175906
transform 1 0 2576 0 1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_37
timestamp 1698175906
transform 1 0 2744 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_101
timestamp 1698175906
transform 1 0 6328 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_107
timestamp 1698175906
transform 1 0 6664 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_171
timestamp 1698175906
transform 1 0 10248 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_177
timestamp 1698175906
transform 1 0 10584 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_241
timestamp 1698175906
transform 1 0 14168 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_247
timestamp 1698175906
transform 1 0 14504 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_311
timestamp 1698175906
transform 1 0 18088 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_317
timestamp 1698175906
transform 1 0 18424 0 1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_2
timestamp 1698175906
transform 1 0 784 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_66
timestamp 1698175906
transform 1 0 4368 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_72
timestamp 1698175906
transform 1 0 4704 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_136
timestamp 1698175906
transform 1 0 8288 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_142
timestamp 1698175906
transform 1 0 8624 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_206
timestamp 1698175906
transform 1 0 12208 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_212
timestamp 1698175906
transform 1 0 12544 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_276
timestamp 1698175906
transform 1 0 16128 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_282
timestamp 1698175906
transform 1 0 16464 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_346
timestamp 1698175906
transform 1 0 20048 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_348
timestamp 1698175906
transform 1 0 20160 0 -1 14896
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698175906
transform 1 0 784 0 1 14896
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698175906
transform 1 0 2576 0 1 14896
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_37
timestamp 1698175906
transform 1 0 2744 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_101
timestamp 1698175906
transform 1 0 6328 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_107
timestamp 1698175906
transform 1 0 6664 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_171
timestamp 1698175906
transform 1 0 10248 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_177
timestamp 1698175906
transform 1 0 10584 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_241
timestamp 1698175906
transform 1 0 14168 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_247
timestamp 1698175906
transform 1 0 14504 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_311
timestamp 1698175906
transform 1 0 18088 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_317
timestamp 1698175906
transform 1 0 18424 0 1 14896
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2
timestamp 1698175906
transform 1 0 784 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_66
timestamp 1698175906
transform 1 0 4368 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_72
timestamp 1698175906
transform 1 0 4704 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_136
timestamp 1698175906
transform 1 0 8288 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_142
timestamp 1698175906
transform 1 0 8624 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_206
timestamp 1698175906
transform 1 0 12208 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_212
timestamp 1698175906
transform 1 0 12544 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_276
timestamp 1698175906
transform 1 0 16128 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_282
timestamp 1698175906
transform 1 0 16464 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_346
timestamp 1698175906
transform 1 0 20048 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_348
timestamp 1698175906
transform 1 0 20160 0 -1 15680
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_2
timestamp 1698175906
transform 1 0 784 0 1 15680
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698175906
transform 1 0 2576 0 1 15680
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_37
timestamp 1698175906
transform 1 0 2744 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_101
timestamp 1698175906
transform 1 0 6328 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_107
timestamp 1698175906
transform 1 0 6664 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_171
timestamp 1698175906
transform 1 0 10248 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_177
timestamp 1698175906
transform 1 0 10584 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_241
timestamp 1698175906
transform 1 0 14168 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_247
timestamp 1698175906
transform 1 0 14504 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_311
timestamp 1698175906
transform 1 0 18088 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_317
timestamp 1698175906
transform 1 0 18424 0 1 15680
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2
timestamp 1698175906
transform 1 0 784 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_66
timestamp 1698175906
transform 1 0 4368 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_72
timestamp 1698175906
transform 1 0 4704 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_136
timestamp 1698175906
transform 1 0 8288 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_142
timestamp 1698175906
transform 1 0 8624 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_206
timestamp 1698175906
transform 1 0 12208 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_212
timestamp 1698175906
transform 1 0 12544 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_276
timestamp 1698175906
transform 1 0 16128 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_282
timestamp 1698175906
transform 1 0 16464 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_346
timestamp 1698175906
transform 1 0 20048 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_348
timestamp 1698175906
transform 1 0 20160 0 -1 16464
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698175906
transform 1 0 784 0 1 16464
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698175906
transform 1 0 2576 0 1 16464
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_37
timestamp 1698175906
transform 1 0 2744 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_101
timestamp 1698175906
transform 1 0 6328 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_107
timestamp 1698175906
transform 1 0 6664 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_171
timestamp 1698175906
transform 1 0 10248 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_177
timestamp 1698175906
transform 1 0 10584 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_241
timestamp 1698175906
transform 1 0 14168 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_247
timestamp 1698175906
transform 1 0 14504 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_311
timestamp 1698175906
transform 1 0 18088 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_317
timestamp 1698175906
transform 1 0 18424 0 1 16464
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_2
timestamp 1698175906
transform 1 0 784 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_66
timestamp 1698175906
transform 1 0 4368 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_72
timestamp 1698175906
transform 1 0 4704 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_136
timestamp 1698175906
transform 1 0 8288 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_142
timestamp 1698175906
transform 1 0 8624 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_206
timestamp 1698175906
transform 1 0 12208 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_212
timestamp 1698175906
transform 1 0 12544 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_276
timestamp 1698175906
transform 1 0 16128 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_282
timestamp 1698175906
transform 1 0 16464 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_346
timestamp 1698175906
transform 1 0 20048 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_348
timestamp 1698175906
transform 1 0 20160 0 -1 17248
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698175906
transform 1 0 784 0 1 17248
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698175906
transform 1 0 2576 0 1 17248
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_37
timestamp 1698175906
transform 1 0 2744 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_101
timestamp 1698175906
transform 1 0 6328 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_107
timestamp 1698175906
transform 1 0 6664 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_171
timestamp 1698175906
transform 1 0 10248 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_177
timestamp 1698175906
transform 1 0 10584 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_241
timestamp 1698175906
transform 1 0 14168 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_247
timestamp 1698175906
transform 1 0 14504 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_311
timestamp 1698175906
transform 1 0 18088 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_317
timestamp 1698175906
transform 1 0 18424 0 1 17248
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2
timestamp 1698175906
transform 1 0 784 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1698175906
transform 1 0 4368 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_72
timestamp 1698175906
transform 1 0 4704 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_136
timestamp 1698175906
transform 1 0 8288 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_142
timestamp 1698175906
transform 1 0 8624 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_206
timestamp 1698175906
transform 1 0 12208 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_212
timestamp 1698175906
transform 1 0 12544 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_276
timestamp 1698175906
transform 1 0 16128 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_282
timestamp 1698175906
transform 1 0 16464 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_346
timestamp 1698175906
transform 1 0 20048 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_348
timestamp 1698175906
transform 1 0 20160 0 -1 18032
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_2
timestamp 1698175906
transform 1 0 784 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698175906
transform 1 0 2576 0 1 18032
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_37
timestamp 1698175906
transform 1 0 2744 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_101
timestamp 1698175906
transform 1 0 6328 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_107
timestamp 1698175906
transform 1 0 6664 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_171
timestamp 1698175906
transform 1 0 10248 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_177
timestamp 1698175906
transform 1 0 10584 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_241
timestamp 1698175906
transform 1 0 14168 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_247
timestamp 1698175906
transform 1 0 14504 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_311
timestamp 1698175906
transform 1 0 18088 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_317
timestamp 1698175906
transform 1 0 18424 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_2
timestamp 1698175906
transform 1 0 784 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_66
timestamp 1698175906
transform 1 0 4368 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_72
timestamp 1698175906
transform 1 0 4704 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_136
timestamp 1698175906
transform 1 0 8288 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_168
timestamp 1698175906
transform 1 0 10080 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_172
timestamp 1698175906
transform 1 0 10304 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_174
timestamp 1698175906
transform 1 0 10416 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_201
timestamp 1698175906
transform 1 0 11928 0 -1 18816
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_209
timestamp 1698175906
transform 1 0 12376 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_238
timestamp 1698175906
transform 1 0 14000 0 -1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_270
timestamp 1698175906
transform 1 0 15792 0 -1 18816
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_278
timestamp 1698175906
transform 1 0 16240 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_282
timestamp 1698175906
transform 1 0 16464 0 -1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_314
timestamp 1698175906
transform 1 0 18256 0 -1 18816
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_330
timestamp 1698175906
transform 1 0 19152 0 -1 18816
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_338
timestamp 1698175906
transform 1 0 19600 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_342
timestamp 1698175906
transform 1 0 19824 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_344
timestamp 1698175906
transform 1 0 19936 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_2
timestamp 1698175906
transform 1 0 784 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_36
timestamp 1698175906
transform 1 0 2688 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_70
timestamp 1698175906
transform 1 0 4592 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_104
timestamp 1698175906
transform 1 0 6496 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_138
timestamp 1698175906
transform 1 0 8400 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_142
timestamp 1698175906
transform 1 0 8624 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_176
timestamp 1698175906
transform 1 0 10528 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_232
timestamp 1698175906
transform 1 0 13664 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_236
timestamp 1698175906
transform 1 0 13888 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_240
timestamp 1698175906
transform 1 0 14112 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_274
timestamp 1698175906
transform 1 0 16016 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_308
timestamp 1698175906
transform 1 0 17920 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_342
timestamp 1698175906
transform 1 0 19824 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_346
timestamp 1698175906
transform 1 0 20048 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_348
timestamp 1698175906
transform 1 0 20160 0 1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita2_24 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 3976 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita2_25
timestamp 1698175906
transform -1 0 10528 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita2_26
timestamp 1698175906
transform 1 0 19992 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10640 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output2
timestamp 1698175906
transform 1 0 18760 0 1 10976
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output3
timestamp 1698175906
transform 1 0 8624 0 -1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output4
timestamp 1698175906
transform 1 0 10808 0 -1 2352
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output5
timestamp 1698175906
transform 1 0 18760 0 -1 14112
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output6
timestamp 1698175906
transform -1 0 2240 0 -1 9408
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output7
timestamp 1698175906
transform 1 0 18760 0 -1 13328
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output8
timestamp 1698175906
transform 1 0 18760 0 -1 10976
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output9
timestamp 1698175906
transform 1 0 18760 0 1 10192
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output10
timestamp 1698175906
transform 1 0 12544 0 -1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output11
timestamp 1698175906
transform 1 0 18760 0 1 12544
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output12
timestamp 1698175906
transform -1 0 2240 0 -1 10976
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output13
timestamp 1698175906
transform 1 0 10640 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output14
timestamp 1698175906
transform -1 0 14000 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output15
timestamp 1698175906
transform 1 0 10472 0 -1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output16
timestamp 1698175906
transform 1 0 18760 0 1 8624
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output17
timestamp 1698175906
transform 1 0 12208 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output18
timestamp 1698175906
transform -1 0 2240 0 1 8624
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output19
timestamp 1698175906
transform 1 0 18760 0 1 13328
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output20
timestamp 1698175906
transform 1 0 8736 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output21
timestamp 1698175906
transform -1 0 2240 0 1 12544
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output22
timestamp 1698175906
transform -1 0 2240 0 -1 8624
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output23
timestamp 1698175906
transform 1 0 18760 0 -1 8624
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_45 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 672 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698175906
transform -1 0 20328 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_46
timestamp 1698175906
transform 1 0 672 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698175906
transform -1 0 20328 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_47
timestamp 1698175906
transform 1 0 672 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698175906
transform -1 0 20328 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_48
timestamp 1698175906
transform 1 0 672 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698175906
transform -1 0 20328 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_49
timestamp 1698175906
transform 1 0 672 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698175906
transform -1 0 20328 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_50
timestamp 1698175906
transform 1 0 672 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698175906
transform -1 0 20328 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_51
timestamp 1698175906
transform 1 0 672 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698175906
transform -1 0 20328 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_52
timestamp 1698175906
transform 1 0 672 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698175906
transform -1 0 20328 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_53
timestamp 1698175906
transform 1 0 672 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698175906
transform -1 0 20328 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_54
timestamp 1698175906
transform 1 0 672 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698175906
transform -1 0 20328 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_55
timestamp 1698175906
transform 1 0 672 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698175906
transform -1 0 20328 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_56
timestamp 1698175906
transform 1 0 672 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698175906
transform -1 0 20328 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_57
timestamp 1698175906
transform 1 0 672 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698175906
transform -1 0 20328 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_58
timestamp 1698175906
transform 1 0 672 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698175906
transform -1 0 20328 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_59
timestamp 1698175906
transform 1 0 672 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698175906
transform -1 0 20328 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_60
timestamp 1698175906
transform 1 0 672 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698175906
transform -1 0 20328 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_61
timestamp 1698175906
transform 1 0 672 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698175906
transform -1 0 20328 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_62
timestamp 1698175906
transform 1 0 672 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698175906
transform -1 0 20328 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_63
timestamp 1698175906
transform 1 0 672 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698175906
transform -1 0 20328 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_64
timestamp 1698175906
transform 1 0 672 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698175906
transform -1 0 20328 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_65
timestamp 1698175906
transform 1 0 672 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698175906
transform -1 0 20328 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_66
timestamp 1698175906
transform 1 0 672 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698175906
transform -1 0 20328 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_67
timestamp 1698175906
transform 1 0 672 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698175906
transform -1 0 20328 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_68
timestamp 1698175906
transform 1 0 672 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698175906
transform -1 0 20328 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_69
timestamp 1698175906
transform 1 0 672 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698175906
transform -1 0 20328 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_70
timestamp 1698175906
transform 1 0 672 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698175906
transform -1 0 20328 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_71
timestamp 1698175906
transform 1 0 672 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698175906
transform -1 0 20328 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_72
timestamp 1698175906
transform 1 0 672 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698175906
transform -1 0 20328 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_73
timestamp 1698175906
transform 1 0 672 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698175906
transform -1 0 20328 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_74
timestamp 1698175906
transform 1 0 672 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698175906
transform -1 0 20328 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_75
timestamp 1698175906
transform 1 0 672 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698175906
transform -1 0 20328 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_76
timestamp 1698175906
transform 1 0 672 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698175906
transform -1 0 20328 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_77
timestamp 1698175906
transform 1 0 672 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698175906
transform -1 0 20328 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_78
timestamp 1698175906
transform 1 0 672 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698175906
transform -1 0 20328 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_79
timestamp 1698175906
transform 1 0 672 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698175906
transform -1 0 20328 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_80
timestamp 1698175906
transform 1 0 672 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698175906
transform -1 0 20328 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_81
timestamp 1698175906
transform 1 0 672 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698175906
transform -1 0 20328 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_82
timestamp 1698175906
transform 1 0 672 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698175906
transform -1 0 20328 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_83
timestamp 1698175906
transform 1 0 672 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698175906
transform -1 0 20328 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_84
timestamp 1698175906
transform 1 0 672 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698175906
transform -1 0 20328 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_85
timestamp 1698175906
transform 1 0 672 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698175906
transform -1 0 20328 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_86
timestamp 1698175906
transform 1 0 672 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698175906
transform -1 0 20328 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_87
timestamp 1698175906
transform 1 0 672 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698175906
transform -1 0 20328 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_88
timestamp 1698175906
transform 1 0 672 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698175906
transform -1 0 20328 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_89
timestamp 1698175906
transform 1 0 672 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698175906
transform -1 0 20328 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_90 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 2576 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_91
timestamp 1698175906
transform 1 0 4480 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_92
timestamp 1698175906
transform 1 0 6384 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_93
timestamp 1698175906
transform 1 0 8288 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_94
timestamp 1698175906
transform 1 0 10192 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_95
timestamp 1698175906
transform 1 0 12096 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_96
timestamp 1698175906
transform 1 0 14000 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_97
timestamp 1698175906
transform 1 0 15904 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_98
timestamp 1698175906
transform 1 0 17808 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_99
timestamp 1698175906
transform 1 0 19712 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_100
timestamp 1698175906
transform 1 0 4592 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_101
timestamp 1698175906
transform 1 0 8512 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_102
timestamp 1698175906
transform 1 0 12432 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_103
timestamp 1698175906
transform 1 0 16352 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_104
timestamp 1698175906
transform 1 0 2632 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_105
timestamp 1698175906
transform 1 0 6552 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_106
timestamp 1698175906
transform 1 0 10472 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_107
timestamp 1698175906
transform 1 0 14392 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_108
timestamp 1698175906
transform 1 0 18312 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_109
timestamp 1698175906
transform 1 0 4592 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_110
timestamp 1698175906
transform 1 0 8512 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_111
timestamp 1698175906
transform 1 0 12432 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_112
timestamp 1698175906
transform 1 0 16352 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_113
timestamp 1698175906
transform 1 0 2632 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_114
timestamp 1698175906
transform 1 0 6552 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_115
timestamp 1698175906
transform 1 0 10472 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_116
timestamp 1698175906
transform 1 0 14392 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_117
timestamp 1698175906
transform 1 0 18312 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_118
timestamp 1698175906
transform 1 0 4592 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_119
timestamp 1698175906
transform 1 0 8512 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_120
timestamp 1698175906
transform 1 0 12432 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_121
timestamp 1698175906
transform 1 0 16352 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_122
timestamp 1698175906
transform 1 0 2632 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_123
timestamp 1698175906
transform 1 0 6552 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_124
timestamp 1698175906
transform 1 0 10472 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_125
timestamp 1698175906
transform 1 0 14392 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_126
timestamp 1698175906
transform 1 0 18312 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_127
timestamp 1698175906
transform 1 0 4592 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_128
timestamp 1698175906
transform 1 0 8512 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_129
timestamp 1698175906
transform 1 0 12432 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_130
timestamp 1698175906
transform 1 0 16352 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_131
timestamp 1698175906
transform 1 0 2632 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_132
timestamp 1698175906
transform 1 0 6552 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_133
timestamp 1698175906
transform 1 0 10472 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_134
timestamp 1698175906
transform 1 0 14392 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_135
timestamp 1698175906
transform 1 0 18312 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_136
timestamp 1698175906
transform 1 0 4592 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_137
timestamp 1698175906
transform 1 0 8512 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_138
timestamp 1698175906
transform 1 0 12432 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_139
timestamp 1698175906
transform 1 0 16352 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_140
timestamp 1698175906
transform 1 0 2632 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_141
timestamp 1698175906
transform 1 0 6552 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_142
timestamp 1698175906
transform 1 0 10472 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_143
timestamp 1698175906
transform 1 0 14392 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_144
timestamp 1698175906
transform 1 0 18312 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_145
timestamp 1698175906
transform 1 0 4592 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_146
timestamp 1698175906
transform 1 0 8512 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_147
timestamp 1698175906
transform 1 0 12432 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_148
timestamp 1698175906
transform 1 0 16352 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_149
timestamp 1698175906
transform 1 0 2632 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_150
timestamp 1698175906
transform 1 0 6552 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_151
timestamp 1698175906
transform 1 0 10472 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_152
timestamp 1698175906
transform 1 0 14392 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_153
timestamp 1698175906
transform 1 0 18312 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_154
timestamp 1698175906
transform 1 0 4592 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_155
timestamp 1698175906
transform 1 0 8512 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_156
timestamp 1698175906
transform 1 0 12432 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_157
timestamp 1698175906
transform 1 0 16352 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_158
timestamp 1698175906
transform 1 0 2632 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_159
timestamp 1698175906
transform 1 0 6552 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_160
timestamp 1698175906
transform 1 0 10472 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_161
timestamp 1698175906
transform 1 0 14392 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_162
timestamp 1698175906
transform 1 0 18312 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_163
timestamp 1698175906
transform 1 0 4592 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_164
timestamp 1698175906
transform 1 0 8512 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_165
timestamp 1698175906
transform 1 0 12432 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_166
timestamp 1698175906
transform 1 0 16352 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_167
timestamp 1698175906
transform 1 0 2632 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_168
timestamp 1698175906
transform 1 0 6552 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_169
timestamp 1698175906
transform 1 0 10472 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_170
timestamp 1698175906
transform 1 0 14392 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_171
timestamp 1698175906
transform 1 0 18312 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_172
timestamp 1698175906
transform 1 0 4592 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_173
timestamp 1698175906
transform 1 0 8512 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_174
timestamp 1698175906
transform 1 0 12432 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_175
timestamp 1698175906
transform 1 0 16352 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_176
timestamp 1698175906
transform 1 0 2632 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_177
timestamp 1698175906
transform 1 0 6552 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_178
timestamp 1698175906
transform 1 0 10472 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_179
timestamp 1698175906
transform 1 0 14392 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_180
timestamp 1698175906
transform 1 0 18312 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_181
timestamp 1698175906
transform 1 0 4592 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_182
timestamp 1698175906
transform 1 0 8512 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_183
timestamp 1698175906
transform 1 0 12432 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_184
timestamp 1698175906
transform 1 0 16352 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_185
timestamp 1698175906
transform 1 0 2632 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_186
timestamp 1698175906
transform 1 0 6552 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_187
timestamp 1698175906
transform 1 0 10472 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_188
timestamp 1698175906
transform 1 0 14392 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_189
timestamp 1698175906
transform 1 0 18312 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_190
timestamp 1698175906
transform 1 0 4592 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_191
timestamp 1698175906
transform 1 0 8512 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_192
timestamp 1698175906
transform 1 0 12432 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_193
timestamp 1698175906
transform 1 0 16352 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_194
timestamp 1698175906
transform 1 0 2632 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_195
timestamp 1698175906
transform 1 0 6552 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_196
timestamp 1698175906
transform 1 0 10472 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_197
timestamp 1698175906
transform 1 0 14392 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_198
timestamp 1698175906
transform 1 0 18312 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_199
timestamp 1698175906
transform 1 0 4592 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_200
timestamp 1698175906
transform 1 0 8512 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_201
timestamp 1698175906
transform 1 0 12432 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_202
timestamp 1698175906
transform 1 0 16352 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_203
timestamp 1698175906
transform 1 0 2632 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_204
timestamp 1698175906
transform 1 0 6552 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_205
timestamp 1698175906
transform 1 0 10472 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_206
timestamp 1698175906
transform 1 0 14392 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_207
timestamp 1698175906
transform 1 0 18312 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_208
timestamp 1698175906
transform 1 0 4592 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_209
timestamp 1698175906
transform 1 0 8512 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_210
timestamp 1698175906
transform 1 0 12432 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_211
timestamp 1698175906
transform 1 0 16352 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_212
timestamp 1698175906
transform 1 0 2632 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_213
timestamp 1698175906
transform 1 0 6552 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_214
timestamp 1698175906
transform 1 0 10472 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_215
timestamp 1698175906
transform 1 0 14392 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_216
timestamp 1698175906
transform 1 0 18312 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_217
timestamp 1698175906
transform 1 0 4592 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_218
timestamp 1698175906
transform 1 0 8512 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_219
timestamp 1698175906
transform 1 0 12432 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_220
timestamp 1698175906
transform 1 0 16352 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_221
timestamp 1698175906
transform 1 0 2632 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_222
timestamp 1698175906
transform 1 0 6552 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_223
timestamp 1698175906
transform 1 0 10472 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_224
timestamp 1698175906
transform 1 0 14392 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_225
timestamp 1698175906
transform 1 0 18312 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_226
timestamp 1698175906
transform 1 0 4592 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_227
timestamp 1698175906
transform 1 0 8512 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_228
timestamp 1698175906
transform 1 0 12432 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_229
timestamp 1698175906
transform 1 0 16352 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_230
timestamp 1698175906
transform 1 0 2632 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_231
timestamp 1698175906
transform 1 0 6552 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_232
timestamp 1698175906
transform 1 0 10472 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_233
timestamp 1698175906
transform 1 0 14392 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_234
timestamp 1698175906
transform 1 0 18312 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_235
timestamp 1698175906
transform 1 0 4592 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_236
timestamp 1698175906
transform 1 0 8512 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_237
timestamp 1698175906
transform 1 0 12432 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_238
timestamp 1698175906
transform 1 0 16352 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_239
timestamp 1698175906
transform 1 0 2632 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_240
timestamp 1698175906
transform 1 0 6552 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_241
timestamp 1698175906
transform 1 0 10472 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_242
timestamp 1698175906
transform 1 0 14392 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_243
timestamp 1698175906
transform 1 0 18312 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_244
timestamp 1698175906
transform 1 0 4592 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_245
timestamp 1698175906
transform 1 0 8512 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_246
timestamp 1698175906
transform 1 0 12432 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_247
timestamp 1698175906
transform 1 0 16352 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_248
timestamp 1698175906
transform 1 0 2632 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_249
timestamp 1698175906
transform 1 0 6552 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_250
timestamp 1698175906
transform 1 0 10472 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_251
timestamp 1698175906
transform 1 0 14392 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_252
timestamp 1698175906
transform 1 0 18312 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_253
timestamp 1698175906
transform 1 0 4592 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_254
timestamp 1698175906
transform 1 0 8512 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_255
timestamp 1698175906
transform 1 0 12432 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_256
timestamp 1698175906
transform 1 0 16352 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_257
timestamp 1698175906
transform 1 0 2632 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_258
timestamp 1698175906
transform 1 0 6552 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_259
timestamp 1698175906
transform 1 0 10472 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_260
timestamp 1698175906
transform 1 0 14392 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_261
timestamp 1698175906
transform 1 0 18312 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_262
timestamp 1698175906
transform 1 0 4592 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_263
timestamp 1698175906
transform 1 0 8512 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_264
timestamp 1698175906
transform 1 0 12432 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_265
timestamp 1698175906
transform 1 0 16352 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_266
timestamp 1698175906
transform 1 0 2632 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_267
timestamp 1698175906
transform 1 0 6552 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_268
timestamp 1698175906
transform 1 0 10472 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_269
timestamp 1698175906
transform 1 0 14392 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_270
timestamp 1698175906
transform 1 0 18312 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_271
timestamp 1698175906
transform 1 0 4592 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_272
timestamp 1698175906
transform 1 0 8512 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_273
timestamp 1698175906
transform 1 0 12432 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_274
timestamp 1698175906
transform 1 0 16352 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_275
timestamp 1698175906
transform 1 0 2632 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_276
timestamp 1698175906
transform 1 0 6552 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_277
timestamp 1698175906
transform 1 0 10472 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_278
timestamp 1698175906
transform 1 0 14392 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_279
timestamp 1698175906
transform 1 0 18312 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_280
timestamp 1698175906
transform 1 0 4592 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_281
timestamp 1698175906
transform 1 0 8512 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_282
timestamp 1698175906
transform 1 0 12432 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_283
timestamp 1698175906
transform 1 0 16352 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_284
timestamp 1698175906
transform 1 0 2632 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_285
timestamp 1698175906
transform 1 0 6552 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_286
timestamp 1698175906
transform 1 0 10472 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_287
timestamp 1698175906
transform 1 0 14392 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_288
timestamp 1698175906
transform 1 0 18312 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_289
timestamp 1698175906
transform 1 0 4592 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_290
timestamp 1698175906
transform 1 0 8512 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_291
timestamp 1698175906
transform 1 0 12432 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_292
timestamp 1698175906
transform 1 0 16352 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_293
timestamp 1698175906
transform 1 0 2576 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_294
timestamp 1698175906
transform 1 0 4480 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_295
timestamp 1698175906
transform 1 0 6384 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_296
timestamp 1698175906
transform 1 0 8288 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_297
timestamp 1698175906
transform 1 0 10192 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_298
timestamp 1698175906
transform 1 0 12096 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_299
timestamp 1698175906
transform 1 0 14000 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_300
timestamp 1698175906
transform 1 0 15904 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_301
timestamp 1698175906
transform 1 0 17808 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_302
timestamp 1698175906
transform 1 0 19712 0 1 18816
box -43 -43 155 435
<< labels >>
flabel metal3 s 0 13776 400 13832 0 FreeSans 224 0 0 0 clk
port 0 nsew signal input
flabel metal2 s 3696 0 3752 400 0 FreeSans 224 90 0 0 segm[0]
port 1 nsew signal tristate
flabel metal2 s 11088 20600 11144 21000 0 FreeSans 224 90 0 0 segm[10]
port 2 nsew signal tristate
flabel metal3 s 20600 10752 21000 10808 0 FreeSans 224 0 0 0 segm[11]
port 3 nsew signal tristate
flabel metal2 s 8400 20600 8456 21000 0 FreeSans 224 90 0 0 segm[12]
port 4 nsew signal tristate
flabel metal2 s 10752 0 10808 400 0 FreeSans 224 90 0 0 segm[13]
port 5 nsew signal tristate
flabel metal3 s 20600 13440 21000 13496 0 FreeSans 224 0 0 0 segm[1]
port 6 nsew signal tristate
flabel metal3 s 0 9072 400 9128 0 FreeSans 224 0 0 0 segm[2]
port 7 nsew signal tristate
flabel metal2 s 9408 20600 9464 21000 0 FreeSans 224 90 0 0 segm[3]
port 8 nsew signal tristate
flabel metal3 s 20600 12768 21000 12824 0 FreeSans 224 0 0 0 segm[4]
port 9 nsew signal tristate
flabel metal3 s 20600 18480 21000 18536 0 FreeSans 224 0 0 0 segm[5]
port 10 nsew signal tristate
flabel metal3 s 20600 10416 21000 10472 0 FreeSans 224 0 0 0 segm[6]
port 11 nsew signal tristate
flabel metal3 s 20600 10080 21000 10136 0 FreeSans 224 0 0 0 segm[7]
port 12 nsew signal tristate
flabel metal2 s 12096 20600 12152 21000 0 FreeSans 224 90 0 0 segm[8]
port 13 nsew signal tristate
flabel metal3 s 20600 12432 21000 12488 0 FreeSans 224 0 0 0 segm[9]
port 14 nsew signal tristate
flabel metal3 s 0 10416 400 10472 0 FreeSans 224 0 0 0 sel[0]
port 15 nsew signal tristate
flabel metal2 s 11088 0 11144 400 0 FreeSans 224 90 0 0 sel[10]
port 16 nsew signal tristate
flabel metal2 s 12768 0 12824 400 0 FreeSans 224 90 0 0 sel[11]
port 17 nsew signal tristate
flabel metal2 s 10416 20600 10472 21000 0 FreeSans 224 90 0 0 sel[1]
port 18 nsew signal tristate
flabel metal3 s 20600 8736 21000 8792 0 FreeSans 224 0 0 0 sel[2]
port 19 nsew signal tristate
flabel metal2 s 11760 20600 11816 21000 0 FreeSans 224 90 0 0 sel[3]
port 20 nsew signal tristate
flabel metal3 s 0 8736 400 8792 0 FreeSans 224 0 0 0 sel[4]
port 21 nsew signal tristate
flabel metal3 s 20600 13104 21000 13160 0 FreeSans 224 0 0 0 sel[5]
port 22 nsew signal tristate
flabel metal2 s 9072 20600 9128 21000 0 FreeSans 224 90 0 0 sel[6]
port 23 nsew signal tristate
flabel metal3 s 0 12432 400 12488 0 FreeSans 224 0 0 0 sel[7]
port 24 nsew signal tristate
flabel metal3 s 0 8400 400 8456 0 FreeSans 224 0 0 0 sel[8]
port 25 nsew signal tristate
flabel metal3 s 20600 8400 21000 8456 0 FreeSans 224 0 0 0 sel[9]
port 26 nsew signal tristate
flabel metal4 s 2224 1538 2384 19238 0 FreeSans 640 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 17584 1538 17744 19238 0 FreeSans 640 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 9904 1538 10064 19238 0 FreeSans 640 90 0 0 vss
port 28 nsew ground bidirectional
rlabel metal1 10500 19208 10500 19208 0 vdd
rlabel metal1 10500 18816 10500 18816 0 vss
rlabel metal3 6524 12684 6524 12684 0 _000_
rlabel metal2 9380 13692 9380 13692 0 _001_
rlabel metal2 5908 10206 5908 10206 0 _002_
rlabel metal2 13188 12236 13188 12236 0 _003_
rlabel metal2 7476 13356 7476 13356 0 _004_
rlabel metal2 11284 13692 11284 13692 0 _005_
rlabel metal2 10220 7140 10220 7140 0 _006_
rlabel metal3 12740 7588 12740 7588 0 _007_
rlabel metal2 13020 9716 13020 9716 0 _008_
rlabel metal2 11200 9660 11200 9660 0 _009_
rlabel metal3 11312 11900 11312 11900 0 _010_
rlabel metal2 10780 11984 10780 11984 0 _011_
rlabel metal2 13020 10948 13020 10948 0 _012_
rlabel metal2 11060 8792 11060 8792 0 _013_
rlabel metal2 12796 12768 12796 12768 0 _014_
rlabel metal2 6860 8512 6860 8512 0 _015_
rlabel metal2 12068 8204 12068 8204 0 _016_
rlabel metal3 8512 13524 8512 13524 0 _017_
rlabel metal2 6020 8092 6020 8092 0 _018_
rlabel metal2 10080 7924 10080 7924 0 _019_
rlabel metal2 8148 8428 8148 8428 0 _020_
rlabel metal2 6132 10948 6132 10948 0 _021_
rlabel metal2 6804 12152 6804 12152 0 _022_
rlabel metal2 13020 8932 13020 8932 0 _023_
rlabel metal3 13440 12460 13440 12460 0 _024_
rlabel metal2 7420 9352 7420 9352 0 _025_
rlabel metal2 12740 9492 12740 9492 0 _026_
rlabel metal2 12068 11480 12068 11480 0 _027_
rlabel metal2 12404 11816 12404 11816 0 _028_
rlabel metal3 8540 13132 8540 13132 0 _029_
rlabel metal2 11564 13468 11564 13468 0 _030_
rlabel metal2 10696 7812 10696 7812 0 _031_
rlabel metal3 9800 9604 9800 9604 0 _032_
rlabel metal2 10164 7896 10164 7896 0 _033_
rlabel metal2 10164 8148 10164 8148 0 _034_
rlabel metal3 12992 7644 12992 7644 0 _035_
rlabel metal3 10696 9548 10696 9548 0 _036_
rlabel metal3 10220 11956 10220 11956 0 _037_
rlabel metal2 13636 10808 13636 10808 0 _038_
rlabel metal3 11844 9996 11844 9996 0 _039_
rlabel metal2 11284 10612 11284 10612 0 _040_
rlabel metal2 10836 9408 10836 9408 0 _041_
rlabel metal2 11732 12208 11732 12208 0 _042_
rlabel metal2 10836 11676 10836 11676 0 _043_
rlabel metal2 8316 9884 8316 9884 0 _044_
rlabel metal2 12824 11284 12824 11284 0 _045_
rlabel metal2 10724 9296 10724 9296 0 _046_
rlabel metal2 13076 13160 13076 13160 0 _047_
rlabel metal2 7364 8764 7364 8764 0 _048_
rlabel metal2 12236 8596 12236 8596 0 _049_
rlabel metal2 8484 10584 8484 10584 0 _050_
rlabel metal2 9828 11256 9828 11256 0 _051_
rlabel metal2 8036 8652 8036 8652 0 _052_
rlabel metal3 7896 10444 7896 10444 0 _053_
rlabel metal2 8820 12488 8820 12488 0 _054_
rlabel metal2 8092 9184 8092 9184 0 _055_
rlabel metal3 8540 10052 8540 10052 0 _056_
rlabel metal2 8820 13328 8820 13328 0 _057_
rlabel metal2 7252 10780 7252 10780 0 _058_
rlabel metal2 6804 10976 6804 10976 0 _059_
rlabel metal2 6972 10724 6972 10724 0 _060_
rlabel metal2 8148 11368 8148 11368 0 _061_
rlabel metal2 9212 10584 9212 10584 0 _062_
rlabel via2 9100 9100 9100 9100 0 _063_
rlabel metal2 7112 10500 7112 10500 0 _064_
rlabel metal3 8904 10836 8904 10836 0 _065_
rlabel metal2 7980 9940 7980 9940 0 _066_
rlabel metal2 10444 9072 10444 9072 0 _067_
rlabel metal2 9632 9156 9632 9156 0 _068_
rlabel metal2 8680 13468 8680 13468 0 _069_
rlabel metal2 9352 10500 9352 10500 0 _070_
rlabel metal2 5880 8820 5880 8820 0 _071_
rlabel metal2 7476 11340 7476 11340 0 _072_
rlabel metal2 7476 9856 7476 9856 0 _073_
rlabel metal2 6132 8820 6132 8820 0 _074_
rlabel metal2 8148 7308 8148 7308 0 _075_
rlabel metal2 7868 10696 7868 10696 0 _076_
rlabel metal2 6748 11816 6748 11816 0 _077_
rlabel metal2 6496 11116 6496 11116 0 _078_
rlabel metal2 6916 10668 6916 10668 0 _079_
rlabel metal2 6888 11956 6888 11956 0 _080_
rlabel metal2 7084 12096 7084 12096 0 _081_
rlabel metal2 12068 9044 12068 9044 0 _082_
rlabel metal2 7812 9072 7812 9072 0 _083_
rlabel metal2 10948 7406 10948 7406 0 _084_
rlabel metal2 13188 8316 13188 8316 0 _085_
rlabel metal2 6440 12068 6440 12068 0 _086_
rlabel metal2 9520 13188 9520 13188 0 _087_
rlabel metal2 13356 13468 13356 13468 0 _088_
rlabel metal2 9772 13468 9772 13468 0 _089_
rlabel metal3 6496 10276 6496 10276 0 _090_
rlabel metal3 1239 13804 1239 13804 0 clk
rlabel metal2 10836 10556 10836 10556 0 clknet_0_clk
rlabel metal2 6636 11256 6636 11256 0 clknet_1_0__leaf_clk
rlabel metal2 14644 12852 14644 12852 0 clknet_1_1__leaf_clk
rlabel metal2 9044 7756 9044 7756 0 dut2.count\[0\]
rlabel metal2 8456 7308 8456 7308 0 dut2.count\[1\]
rlabel metal3 6020 10108 6020 10108 0 dut2.count\[2\]
rlabel metal2 7420 11368 7420 11368 0 dut2.count\[3\]
rlabel metal2 10696 15960 10696 15960 0 net1
rlabel metal2 12180 13020 12180 13020 0 net10
rlabel metal2 14028 12768 14028 12768 0 net11
rlabel metal2 4844 10416 4844 10416 0 net12
rlabel metal2 10724 2982 10724 2982 0 net13
rlabel metal2 13692 2982 13692 2982 0 net14
rlabel metal2 10108 13664 10108 13664 0 net15
rlabel metal2 14084 8904 14084 8904 0 net16
rlabel metal2 11788 13664 11788 13664 0 net17
rlabel metal2 6356 9044 6356 9044 0 net18
rlabel metal3 15190 13188 15190 13188 0 net19
rlabel metal2 14084 10948 14084 10948 0 net2
rlabel metal2 9044 17486 9044 17486 0 net20
rlabel metal3 3178 12740 3178 12740 0 net21
rlabel metal2 5796 8540 5796 8540 0 net22
rlabel metal3 15960 8484 15960 8484 0 net23
rlabel metal2 3724 1015 3724 1015 0 net24
rlabel metal2 9436 19789 9436 19789 0 net25
rlabel metal2 20132 18592 20132 18592 0 net26
rlabel metal2 8540 14770 8540 14770 0 net3
rlabel metal3 10696 2156 10696 2156 0 net4
rlabel metal2 18956 13692 18956 13692 0 net5
rlabel metal2 5012 8652 5012 8652 0 net6
rlabel metal2 14084 13104 14084 13104 0 net7
rlabel metal2 13748 10976 13748 10976 0 net8
rlabel metal2 18844 10024 18844 10024 0 net9
rlabel metal2 11116 19873 11116 19873 0 segm[10]
rlabel metal2 20020 11004 20020 11004 0 segm[11]
rlabel metal2 8428 19677 8428 19677 0 segm[12]
rlabel metal2 10780 1211 10780 1211 0 segm[13]
rlabel metal2 19964 13664 19964 13664 0 segm[1]
rlabel metal3 679 9100 679 9100 0 segm[2]
rlabel metal2 19964 12936 19964 12936 0 segm[4]
rlabel metal2 19964 10584 19964 10584 0 segm[6]
rlabel metal2 20020 10276 20020 10276 0 segm[7]
rlabel metal2 12124 19677 12124 19677 0 segm[8]
rlabel metal2 20020 12628 20020 12628 0 segm[9]
rlabel metal3 679 10444 679 10444 0 sel[0]
rlabel metal2 11116 1015 11116 1015 0 sel[10]
rlabel metal2 12796 1099 12796 1099 0 sel[11]
rlabel metal2 10444 19677 10444 19677 0 sel[1]
rlabel metal2 20020 8820 20020 8820 0 sel[2]
rlabel metal2 11788 19873 11788 19873 0 sel[3]
rlabel metal3 679 8764 679 8764 0 sel[4]
rlabel metal2 20020 13356 20020 13356 0 sel[5]
rlabel metal2 9100 19873 9100 19873 0 sel[6]
rlabel metal3 679 12460 679 12460 0 sel[7]
rlabel metal3 679 8428 679 8428 0 sel[8]
rlabel metal2 20020 8400 20020 8400 0 sel[9]
<< properties >>
string FIXED_BBOX 0 0 21000 21000
<< end >>
