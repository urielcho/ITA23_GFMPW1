// This is the unpowered netlist.
module ita (clk,
    io_oeb,
    itasegm,
    itasel,
    nsel,
    segm,
    sel);
 input clk;
 output [37:0] io_oeb;
 input [895:0] itasegm;
 input [767:0] itasel;
 input [5:0] nsel;
 output [13:0] segm;
 output [11:0] sel;

 wire net1855;
 wire net1865;
 wire net1866;
 wire net1829;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1856;
 wire net1837;
 wire net1838;
 wire net1839;
 wire net1840;
 wire net1841;
 wire net1842;
 wire net1843;
 wire net1844;
 wire net1845;
 wire net1846;
 wire net1857;
 wire net1847;
 wire net1848;
 wire net1849;
 wire net1850;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1858;
 wire net1859;
 wire net1860;
 wire net1861;
 wire net1862;
 wire net1863;
 wire net1864;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire net1;
 wire net10;
 wire net100;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net101;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net102;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net103;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net104;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net105;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net106;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net107;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net108;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net109;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net11;
 wire net110;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net111;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net112;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net113;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net114;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net115;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net116;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net117;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net118;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net119;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net12;
 wire net120;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net121;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net122;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net123;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net124;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net125;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net126;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net127;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net128;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net129;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net13;
 wire net130;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net131;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net132;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net133;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net134;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net135;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net136;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net137;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net138;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net139;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net14;
 wire net140;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net141;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net142;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net143;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net144;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net145;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net146;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net147;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net148;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net149;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net15;
 wire net150;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net151;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net152;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net153;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net154;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net155;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net156;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net157;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net158;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net159;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net16;
 wire net160;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net161;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net162;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net163;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net164;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net165;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net166;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net167;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net168;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net169;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net17;
 wire net170;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net171;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net172;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net173;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net174;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net175;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net176;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net177;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net178;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net179;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net18;
 wire net180;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net181;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net182;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net73;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net74;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net75;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net76;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net77;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net78;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net79;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net8;
 wire net80;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net81;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net82;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net83;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net84;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net85;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net86;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net87;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net88;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net89;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net9;
 wire net90;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net91;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net92;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net93;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net94;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net95;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net96;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net97;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net98;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net99;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;

 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_1 (.I(_0050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_10 (.I(net749));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_11 (.I(net749));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_12 (.I(net749));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_13 (.I(net749));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_14 (.I(net749));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_15 (.I(net758));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_16 (.I(net758));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_17 (.I(net989));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_18 (.I(net989));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_19 (.I(net1517));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_2 (.I(_0050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_20 (.I(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_21 (.I(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_22 (.I(_1806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_23 (.I(net126));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_24 (.I(net126));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_25 (.I(net748));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_26 (.I(net748));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_27 (.I(net750));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_28 (.I(net750));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_29 (.I(net751));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_3 (.I(_0050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_30 (.I(net751));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_31 (.I(net751));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_32 (.I(net751));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_33 (.I(net752));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_34 (.I(net752));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_35 (.I(net752));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_36 (.I(net752));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_37 (.I(net752));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_38 (.I(net994));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_39 (.I(net994));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_4 (.I(_0226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_40 (.I(net1685));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_41 (.I(net1685));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_42 (.I(net1685));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_43 (.I(net1685));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_5 (.I(_0226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_6 (.I(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_7 (.I(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_8 (.I(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_9 (.I(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2335__I (.I(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2336__I (.I(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2337__I (.I(_0207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2338__I (.I(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2339__I (.I(_0151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2340__I (.I(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2343__A1 (.I(net862));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2343__B2 (.I(net785));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2343__C (.I(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2344__I (.I(_0227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2346__I (.I(_0231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2349__I (.I(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2350__I (.I(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2354__A1 (.I(_0969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2354__A3 (.I(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2354__B2 (.I(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2355__A1 (.I(net801));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2355__B2 (.I(net816));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2355__C (.I(_0975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2357__I (.I(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2359__I (.I(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2361__I (.I(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2362__I (.I(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2363__I (.I(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2364__I (.I(_0984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2366__B2 (.I(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2367__A1 (.I(net179));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2367__A2 (.I(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2367__B1 (.I(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2367__B2 (.I(net888));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2367__C (.I(_0987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2368__I (.I(_0261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2369__I (.I(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2370__I (.I(_0264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2371__I (.I(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2373__I (.I(_0268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2374__I (.I(_0994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2375__I (.I(_0271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2376__I (.I(_0996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2378__A1 (.I(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2379__B2 (.I(net753));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2379__C (.I(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2380__A1 (.I(net1813));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2380__A2 (.I(net1811));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2380__A4 (.I(_1000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2382__I (.I(_1002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2384__I (.I(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2387__I (.I(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2389__I (.I(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2390__A1 (.I(net645));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2390__B2 (.I(net536));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2392__I (.I(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2394__I (.I(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2397__I (.I(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2399__I (.I(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2400__A1 (.I(net412));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2400__B2 (.I(net583));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2401__A1 (.I(_1006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2401__A2 (.I(_1011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2401__A3 (.I(_1016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2406__A1 (.I(net303));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2406__A2 (.I(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2406__B1 (.I(_1026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2408__I (.I(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2411__A1 (.I(net318));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2411__A2 (.I(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2411__B1 (.I(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2413__I (.I(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2416__A2 (.I(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2416__B1 (.I(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2419__I (.I(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2420__I (.I(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2421__A2 (.I(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2421__B2 (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2422__A1 (.I(_1027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2422__A2 (.I(_1032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2422__A3 (.I(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2422__A4 (.I(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2423__A2 (.I(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2424__A1 (.I(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2424__B1 (.I(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2424__B2 (.I(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2425__I (.I(net896));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2427__A1 (.I(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2428__A1 (.I(net521));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2433__A2 (.I(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2433__A3 (.I(_1050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2433__A4 (.I(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2434__I (.I(net460));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2440__A1 (.I(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2440__A2 (.I(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2440__A3 (.I(_0890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2441__A2 (.I(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2441__B1 (.I(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2441__C (.I(_1060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2444__A2 (.I(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2444__B1 (.I(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2445__A2 (.I(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2445__B1 (.I(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2445__C (.I(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2446__A1 (.I(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2446__A2 (.I(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2446__A3 (.I(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2446__A4 (.I(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2447__A1 (.I(net467));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2447__A2 (.I(_0911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2447__B1 (.I(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2447__B2 (.I(net102));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2448__A1 (.I(net661));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2448__B2 (.I(net133));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2450__A2 (.I(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2450__B1 (.I(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2451__A1 (.I(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2451__A3 (.I(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2451__A4 (.I(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2452__A2 (.I(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2452__B2 (.I(net739));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2453__A1 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2453__B2 (.I(net311));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2454__A1 (.I(net366));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2454__B1 (.I(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2454__B2 (.I(net273));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2455__A1 (.I(net336));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2456__A1 (.I(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2456__A2 (.I(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2456__A4 (.I(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2457__A2 (.I(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2461__A1 (.I(net863));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2461__B2 (.I(net786));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2461__C (.I(_1080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2464__A1 (.I(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2464__A3 (.I(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2464__B2 (.I(_1083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2465__A1 (.I(net802));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2465__B2 (.I(net817));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2465__C (.I(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2468__B2 (.I(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2469__A1 (.I(net180));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2469__A2 (.I(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2469__B1 (.I(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2469__B2 (.I(net889));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2469__C (.I(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2472__A1 (.I(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2473__B2 (.I(net754));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2473__C (.I(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2474__A1 (.I(net1809));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2474__A2 (.I(net1807));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2474__A4 (.I(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2476__A1 (.I(net646));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2476__B2 (.I(net537));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2478__A1 (.I(net413));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2478__B2 (.I(net584));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2479__A1 (.I(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2479__A2 (.I(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2479__A3 (.I(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2480__A1 (.I(net304));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2480__A2 (.I(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2480__B1 (.I(_1026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2481__A1 (.I(net319));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2481__A2 (.I(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2481__B1 (.I(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2482__A2 (.I(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2482__B1 (.I(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2483__A2 (.I(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2483__B2 (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2484__A1 (.I(_1100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2484__A2 (.I(_1101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2484__A3 (.I(_1102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2484__A4 (.I(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2485__A2 (.I(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2486__B1 (.I(_1077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2486__B2 (.I(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2489__A1 (.I(_1107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2490__A1 (.I(net523));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2493__A3 (.I(_1111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2496__A2 (.I(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2496__A3 (.I(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2496__A4 (.I(_1114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2497__I (.I(net461));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2499__A1 (.I(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2502__I (.I(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2504__A1 (.I(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2504__A3 (.I(_0890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2504__B2 (.I(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2505__A2 (.I(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2505__B1 (.I(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2505__C (.I(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2508__A2 (.I(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2508__B1 (.I(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2509__A2 (.I(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2509__B1 (.I(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2509__C (.I(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2510__A1 (.I(_1115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2510__A2 (.I(_1119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2510__A3 (.I(_1124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2510__A4 (.I(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2511__A1 (.I(net478));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2511__A2 (.I(_0911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2511__B1 (.I(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2511__B2 (.I(net103));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2512__A1 (.I(net662));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2512__B2 (.I(net135));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2514__A2 (.I(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2514__B1 (.I(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2515__A1 (.I(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2515__A3 (.I(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2515__A4 (.I(_1133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2516__A2 (.I(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2516__B2 (.I(net740));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2517__B2 (.I(net322));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2518__A1 (.I(net368));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2518__B1 (.I(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2518__B2 (.I(net274));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2519__I (.I(_0012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2520__A1 (.I(net337));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2521__A1 (.I(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2521__A2 (.I(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2521__A4 (.I(_1139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2522__A2 (.I(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2526__A1 (.I(net864));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2526__B2 (.I(net787));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2526__C (.I(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2528__I (.I(_0066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2531__A1 (.I(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2531__A3 (.I(_1148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2531__B2 (.I(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2532__A1 (.I(net803));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2532__B2 (.I(net818));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2532__C (.I(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2535__B2 (.I(_1153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2536__A1 (.I(net181));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2536__A2 (.I(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2536__B1 (.I(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2536__B2 (.I(net890));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2536__C (.I(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2539__A1 (.I(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2540__B2 (.I(net756));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2540__C (.I(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2541__A1 (.I(net1805));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2541__A2 (.I(net1803));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2541__A4 (.I(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2543__A1 (.I(net647));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2543__B2 (.I(net538));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2545__A1 (.I(net414));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2545__B2 (.I(net585));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2546__A1 (.I(_1161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2546__A2 (.I(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2546__A3 (.I(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2547__A1 (.I(net305));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2547__A2 (.I(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2547__B1 (.I(_1026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2548__A1 (.I(net320));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2548__A2 (.I(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2548__B1 (.I(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2549__A2 (.I(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2549__B1 (.I(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2550__A2 (.I(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2551__A4 (.I(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2552__A2 (.I(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2552__A3 (.I(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2553__A1 (.I(_1106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2553__B1 (.I(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2553__B2 (.I(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2556__A1 (.I(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2557__A1 (.I(net524));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2559__A3 (.I(_1111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2562__A2 (.I(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2562__A3 (.I(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2562__A4 (.I(_1179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2563__I (.I(net462));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2565__A1 (.I(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2569__A1 (.I(_1185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2569__A3 (.I(_0890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2569__B2 (.I(_1186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2570__A2 (.I(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2570__B1 (.I(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2570__C (.I(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2573__A2 (.I(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2573__B1 (.I(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2574__A2 (.I(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2574__B1 (.I(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2574__C (.I(_1191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2575__A1 (.I(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2575__A2 (.I(_1184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2575__A3 (.I(_1188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2575__A4 (.I(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2576__A1 (.I(net489));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2576__A2 (.I(_0911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2576__B1 (.I(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2576__B2 (.I(net104));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2577__A1 (.I(net663));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2577__B2 (.I(net136));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2579__A2 (.I(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2579__B1 (.I(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2580__A1 (.I(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2580__A3 (.I(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2580__A4 (.I(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2581__A2 (.I(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2581__B2 (.I(net741));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2582__A1 (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2582__B2 (.I(net333));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2583__A1 (.I(net369));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2583__B1 (.I(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2583__B2 (.I(net275));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2585__A1 (.I(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2585__A2 (.I(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2586__A2 (.I(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2590__A1 (.I(net865));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2590__B2 (.I(net788));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2590__C (.I(_1207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2593__A1 (.I(_1209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2593__A3 (.I(_1148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2593__B2 (.I(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2594__A1 (.I(net804));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2594__B2 (.I(net819));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2594__C (.I(_1211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2597__B2 (.I(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2598__A1 (.I(net182));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2598__A2 (.I(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2598__B1 (.I(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2598__B2 (.I(net891));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2598__C (.I(_1215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2601__A1 (.I(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2602__A1 (.I(net800));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2602__B2 (.I(net757));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2602__C (.I(_1219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2603__A1 (.I(net1801));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2603__A2 (.I(net1799));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2603__A4 (.I(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2605__A1 (.I(net648));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2605__B2 (.I(net539));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2607__A1 (.I(net415));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2607__B2 (.I(net586));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2608__A1 (.I(_1222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2608__A2 (.I(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2608__A3 (.I(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2609__A1 (.I(net306));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2609__A2 (.I(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2609__B1 (.I(_1026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2610__A1 (.I(net321));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2610__A2 (.I(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2610__B1 (.I(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2611__A2 (.I(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2611__B1 (.I(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2612__A2 (.I(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2612__B2 (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2613__A2 (.I(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2613__A4 (.I(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2614__A2 (.I(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2614__A3 (.I(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2615__A1 (.I(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2615__B1 (.I(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2615__B2 (.I(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2617__I (.I(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2619__I (.I(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2620__I (.I(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2621__A2 (.I(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2621__A3 (.I(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2622__I (.I(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2623__I (.I(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2624__A1 (.I(net525));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2626__I (.I(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2627__A2 (.I(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2627__A3 (.I(_1111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2629__I (.I(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2630__I (.I(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2632__A2 (.I(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2632__A3 (.I(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2633__I (.I(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2634__I (.I(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2635__I (.I(net463));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2636__I (.I(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2637__I (.I(_0079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2638__I (.I(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2640__A1 (.I(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2640__B2 (.I(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2641__A2 (.I(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2641__B1 (.I(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2641__B2 (.I(net431));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2645__I (.I(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2646__I (.I(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2648__A1 (.I(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2648__B2 (.I(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2649__A2 (.I(_1259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2649__B1 (.I(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2649__C (.I(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2650__I (.I(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2651__I (.I(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2653__I (.I(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2654__I (.I(_0127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2655__I (.I(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2657__A2 (.I(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2657__A3 (.I(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2657__B1 (.I(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2658__A2 (.I(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2658__B1 (.I(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2658__C (.I(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2659__A1 (.I(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2659__A2 (.I(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2659__A3 (.I(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2659__A4 (.I(_1275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2660__I (.I(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2661__I (.I(_0912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2662__A1 (.I(net500));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2662__B2 (.I(net105));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2663__I (.I(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2664__I (.I(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2665__A1 (.I(net664));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2665__B2 (.I(net137));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2668__A1 (.I(net727));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2668__A2 (.I(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2668__B1 (.I(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2671__A2 (.I(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2671__B1 (.I(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2672__A1 (.I(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2672__A3 (.I(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2672__A4 (.I(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2673__I (.I(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2674__I (.I(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2675__A2 (.I(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2675__B1 (.I(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2675__B2 (.I(net742));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2676__I (.I(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2677__I (.I(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2678__A2 (.I(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2678__B1 (.I(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2678__B2 (.I(net345));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2679__I (.I(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2680__I (.I(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2681__A1 (.I(net370));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2681__A2 (.I(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2681__B1 (.I(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2681__B2 (.I(net276));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2682__I (.I(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2683__A2 (.I(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2684__A2 (.I(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2685__A2 (.I(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2685__A3 (.I(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2686__I (.I(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2687__I (.I(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2689__I (.I(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2690__I (.I(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2691__I (.I(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2692__A1 (.I(net882));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2692__A2 (.I(_1307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2692__A3 (.I(_1308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2693__A2 (.I(_1306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2694__A1 (.I(net867));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2694__A2 (.I(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2694__B1 (.I(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2694__B2 (.I(net790));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2694__C (.I(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2698__I (.I(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2700__I (.I(net836));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2701__A1 (.I(_1314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2701__A3 (.I(_1148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2702__A1 (.I(net805));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2702__B2 (.I(net820));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2702__C (.I(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2703__I (.I(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2704__I (.I(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2706__I (.I(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2707__I (.I(_0984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2709__A1 (.I(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2709__B2 (.I(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2710__A1 (.I(net183));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2710__B2 (.I(net892));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2710__C (.I(_1326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2711__I (.I(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2712__I (.I(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2714__I (.I(_0994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2715__I (.I(_0996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2717__A1 (.I(_1330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2717__A2 (.I(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2717__B1 (.I(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2718__B2 (.I(net758));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2719__A1 (.I(net1797));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2719__A2 (.I(net1795));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2719__A4 (.I(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2720__I (.I(_1002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2721__I (.I(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2722__A2 (.I(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2722__B1 (.I(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2723__I (.I(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2724__I (.I(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2725__A1 (.I(net649));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2725__B1 (.I(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2726__I (.I(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2727__I (.I(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2728__A2 (.I(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2728__B1 (.I(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2729__I (.I(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2730__I (.I(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2731__A1 (.I(net416));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2731__A2 (.I(_1346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2731__B1 (.I(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2731__B2 (.I(net587));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2732__A1 (.I(_1339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2732__A2 (.I(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2732__A3 (.I(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2735__A1 (.I(net307));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2735__A2 (.I(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2735__B1 (.I(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2735__B2 (.I(net59));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2736__I (.I(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2738__A1 (.I(net323));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2738__B2 (.I(net74));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2739__I (.I(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2741__A2 (.I(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2741__B1 (.I(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2743__I (.I(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2744__A2 (.I(_1359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2744__B1 (.I(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2744__B2 (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2745__A3 (.I(_1358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2745__A4 (.I(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2746__A2 (.I(_1349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2747__A1 (.I(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2747__B1 (.I(net1704));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2747__B2 (.I(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2748__I (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2750__A2 (.I(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2750__A3 (.I(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2751__A1 (.I(net526));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2753__A2 (.I(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2753__A3 (.I(_1111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2756__A2 (.I(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2756__A3 (.I(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2757__I (.I(net464));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2759__A1 (.I(_1373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2759__B2 (.I(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2760__A2 (.I(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2760__B1 (.I(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2760__B2 (.I(net432));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2763__A1 (.I(_1377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2763__B2 (.I(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2764__A2 (.I(_1259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2764__B1 (.I(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2764__C (.I(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2767__A2 (.I(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2767__A3 (.I(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2767__B1 (.I(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2768__A2 (.I(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2768__B1 (.I(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2768__C (.I(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2769__A1 (.I(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2769__A2 (.I(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2769__A3 (.I(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2769__A4 (.I(_1384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2770__A1 (.I(net511));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2770__B2 (.I(net106));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2771__A1 (.I(net665));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2771__B2 (.I(net138));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2772__A1 (.I(net728));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2772__A2 (.I(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2772__B1 (.I(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2773__A2 (.I(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2773__B1 (.I(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2774__A1 (.I(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2774__A3 (.I(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2774__A4 (.I(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2775__A2 (.I(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2775__B1 (.I(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2775__B2 (.I(net743));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2776__A2 (.I(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2776__B1 (.I(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2776__B2 (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2777__A1 (.I(net371));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2777__A2 (.I(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2777__B1 (.I(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2777__B2 (.I(net277));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2778__A2 (.I(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2779__A2 (.I(_1392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2780__A2 (.I(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2782__A1 (.I(net883));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2782__A2 (.I(_1307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2782__A3 (.I(_1308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2783__A2 (.I(_1306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2784__A1 (.I(net868));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2784__A2 (.I(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2784__B1 (.I(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2784__B2 (.I(net791));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2784__C (.I(_1399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2787__A1 (.I(_1401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2787__A3 (.I(_1148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2787__B2 (.I(_1402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2788__A1 (.I(net806));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2788__B2 (.I(net821));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2788__C (.I(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2791__A1 (.I(_1405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2791__B2 (.I(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2792__A1 (.I(net184));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2792__B2 (.I(net893));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2792__C (.I(_1407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2795__A1 (.I(_1409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2795__A2 (.I(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2795__B1 (.I(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2796__B2 (.I(net759));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2797__A1 (.I(net1793));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2797__A2 (.I(net1791));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2797__A4 (.I(_1412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2798__A2 (.I(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2798__B1 (.I(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2799__A1 (.I(net650));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2799__B1 (.I(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2800__A2 (.I(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2800__B1 (.I(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2801__A1 (.I(net417));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2801__A2 (.I(_1346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2801__B1 (.I(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2801__B2 (.I(net588));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2802__A1 (.I(_1414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2802__A2 (.I(_1415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2802__A3 (.I(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2803__A1 (.I(net308));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2803__A2 (.I(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2803__B1 (.I(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2803__B2 (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2804__A1 (.I(net324));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2804__B2 (.I(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2805__A2 (.I(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2805__B1 (.I(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2805__B2 (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2806__A2 (.I(_1359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2806__B1 (.I(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2806__B2 (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2807__A3 (.I(_1421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2807__A4 (.I(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2808__A2 (.I(_1418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2809__B1 (.I(_1396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2809__B2 (.I(_1424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2810__I (.I(net897));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2812__A1 (.I(_1426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2812__A2 (.I(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2812__A3 (.I(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2813__A1 (.I(net1319));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2815__I (.I(_0028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2816__A2 (.I(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2818__A1 (.I(_1432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2819__A2 (.I(_1428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2819__A3 (.I(_1431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2820__I (.I(net1266));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2822__A1 (.I(_1435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2823__A1 (.I(net1212));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2823__A2 (.I(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2823__B1 (.I(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2825__I (.I(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2827__A1 (.I(_1439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2828__A2 (.I(_1259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2828__B1 (.I(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2828__C (.I(_1442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2831__A2 (.I(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2831__A3 (.I(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2831__B1 (.I(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2832__A2 (.I(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2832__B1 (.I(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2832__C (.I(_1446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2833__A1 (.I(net1790));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2833__A2 (.I(net1789));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2833__A3 (.I(_1443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2834__A1 (.I(net1196));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2835__A1 (.I(net1438));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2835__B2 (.I(net986));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2836__A2 (.I(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2836__B1 (.I(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2837__A2 (.I(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2837__B1 (.I(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2838__A1 (.I(_1449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2838__A3 (.I(_1451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2838__A4 (.I(_1452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2839__A2 (.I(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2839__B1 (.I(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2839__B2 (.I(net1505));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2840__A2 (.I(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2840__B1 (.I(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2840__B2 (.I(net1063));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2841__A1 (.I(net1186));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2841__A2 (.I(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2841__B1 (.I(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2841__B2 (.I(net1105));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2843__A1 (.I(net1159));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2843__A2 (.I(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2844__A1 (.I(_1454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2844__A2 (.I(_1455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2844__A3 (.I(_1456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2845__A2 (.I(_1453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2845__A3 (.I(_1459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2847__A2 (.I(_1307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2847__A3 (.I(_1308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2848__A2 (.I(_1306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2849__A1 (.I(net1612));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2849__A2 (.I(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2849__B1 (.I(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2849__B2 (.I(net1545));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2849__C (.I(_1463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2853__A1 (.I(_1465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2854__A1 (.I(net1558));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2854__B2 (.I(net1572));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2854__C (.I(_1468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2855__I (.I(net1039));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2857__B2 (.I(_1471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2858__A1 (.I(net1026));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2858__B2 (.I(net1596));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2858__C (.I(_1472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2861__A1 (.I(_1474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2861__A2 (.I(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2861__B1 (.I(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2862__A1 (.I(net1463));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2862__B2 (.I(net1519));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2862__C (.I(_1476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2863__A1 (.I(net1787));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2863__A2 (.I(net1785));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2863__A4 (.I(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2864__A2 (.I(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2864__B1 (.I(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2865__A1 (.I(net1425));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2865__B1 (.I(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2865__B2 (.I(net1332));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2866__A2 (.I(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2866__B1 (.I(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2867__A1 (.I(net1225));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2867__A2 (.I(_1346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2867__B1 (.I(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2867__B2 (.I(net1372));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2868__A1 (.I(_1479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2868__A2 (.I(_1480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2868__A3 (.I(_1481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2869__A1 (.I(net1133));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2869__A2 (.I(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2869__B1 (.I(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2869__B2 (.I(net920));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2870__A1 (.I(net1146));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2870__B2 (.I(net933));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2871__A2 (.I(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2871__B1 (.I(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2872__A2 (.I(_1359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2872__B1 (.I(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2873__A3 (.I(_1486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2873__A4 (.I(_1487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2874__A1 (.I(_1478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2874__A2 (.I(_1483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2875__A1 (.I(_1425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2875__B1 (.I(_1460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2875__B2 (.I(_1489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2878__A2 (.I(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2878__A3 (.I(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2879__A1 (.I(net1320));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2881__A2 (.I(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2883__A1 (.I(_1496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2884__A2 (.I(_1493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2885__I (.I(net1267));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2887__A1 (.I(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2888__A2 (.I(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2888__B1 (.I(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2891__A1 (.I(_1503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2892__A2 (.I(_1259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2892__B1 (.I(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2892__C (.I(_1505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2895__A2 (.I(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2895__A3 (.I(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2895__B1 (.I(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2896__A2 (.I(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2896__B1 (.I(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2896__C (.I(_1509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2897__A1 (.I(net1784));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2897__A2 (.I(net1783));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2897__A3 (.I(_1506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2898__A1 (.I(net1207));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2898__B2 (.I(net960));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2899__A1 (.I(net1439));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2899__B2 (.I(net987));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2900__A2 (.I(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2900__B1 (.I(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2901__A2 (.I(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2901__B1 (.I(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2902__A1 (.I(_1512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2902__A3 (.I(_1514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2902__A4 (.I(_1515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2903__A2 (.I(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2903__B1 (.I(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2903__B2 (.I(net1506));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2904__A2 (.I(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2904__B1 (.I(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2904__B2 (.I(net1074));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2905__A1 (.I(net1187));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2905__A2 (.I(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2905__B1 (.I(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2905__B2 (.I(net1106));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2906__A1 (.I(net1160));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2906__A2 (.I(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2907__A1 (.I(_1517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2907__A2 (.I(_1518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2907__A3 (.I(_1519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2908__A2 (.I(_1516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2910__A2 (.I(_1307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2910__A3 (.I(_1308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2911__A2 (.I(_1306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2912__A1 (.I(net1613));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2912__A2 (.I(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2912__B1 (.I(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2912__B2 (.I(net1546));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2912__C (.I(_1525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2915__A1 (.I(_1527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2916__A1 (.I(net1559));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2916__B2 (.I(net1573));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2916__C (.I(_1529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2917__I (.I(net1040));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2919__B2 (.I(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2920__A1 (.I(net1027));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2920__B2 (.I(net1607));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2920__C (.I(_1533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2921__I (.I(net941));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2923__A1 (.I(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2923__A2 (.I(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2923__B1 (.I(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2924__A1 (.I(net1474));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2924__B2 (.I(net1520));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2924__C (.I(_1537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2925__A1 (.I(net1781));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2925__A2 (.I(net1779));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2925__A4 (.I(_1538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2926__A2 (.I(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2926__B1 (.I(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2927__A1 (.I(net1426));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2927__B1 (.I(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2927__B2 (.I(net1333));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2928__A2 (.I(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2928__B1 (.I(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2929__A1 (.I(net1226));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2929__A2 (.I(_1346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2929__B1 (.I(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2929__B2 (.I(net1373));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2930__A1 (.I(_1540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2930__A2 (.I(_1541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2930__A3 (.I(_1542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2931__A1 (.I(net1134));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2931__A2 (.I(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2931__B1 (.I(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2931__B2 (.I(net921));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2932__A1 (.I(net1147));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2932__B2 (.I(net934));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2933__A2 (.I(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2933__B1 (.I(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2934__A2 (.I(_1359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2934__B1 (.I(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2935__A3 (.I(_1547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2935__A4 (.I(_1548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2936__A2 (.I(_1544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2937__A1 (.I(_1490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2937__B1 (.I(_1522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2937__B2 (.I(_1550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2939__I (.I(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2941__I (.I(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2942__I (.I(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2944__I (.I(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2945__I (.I(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2946__A1 (.I(net1321));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2948__I (.I(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2951__I (.I(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2952__I (.I(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2954__A2 (.I(_1559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2954__A3 (.I(_1562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2955__I (.I(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2956__I (.I(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2957__I (.I(net1268));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2958__I (.I(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2959__I (.I(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2960__I (.I(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2962__B2 (.I(_1574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2963__B2 (.I(net1242));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2967__I (.I(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2968__I (.I(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2970__A1 (.I(_1579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2971__C (.I(_1583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2972__I (.I(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2973__I (.I(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2974__I (.I(net1015));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2975__I (.I(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2976__I (.I(_0102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2977__I (.I(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2978__I (.I(net1001));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2980__C (.I(_1592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2981__A1 (.I(_1567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2981__A2 (.I(_1576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2981__A3 (.I(_1584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2981__A4 (.I(_1593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2982__I (.I(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2983__I (.I(_0912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2984__A1 (.I(net1218));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2984__B2 (.I(net961));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2985__I (.I(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2986__I (.I(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2987__A1 (.I(net1441));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2987__B2 (.I(net988));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2994__A1 (.I(_1597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2994__A3 (.I(_1603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2994__A4 (.I(_1606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2995__I (.I(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2996__I (.I(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2997__B2 (.I(net1508));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2998__I (.I(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2999__I (.I(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3000__A1 (.I(net1649));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3000__B2 (.I(net1085));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3001__I (.I(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3002__I (.I(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3003__A1 (.I(net1188));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3003__B2 (.I(net1108));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3004__I (.I(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3005__A1 (.I(net1161));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3006__A1 (.I(_1610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3006__A2 (.I(_1613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3007__A2 (.I(_1607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3008__I (.I(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3009__I (.I(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3011__I (.I(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3012__I (.I(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3013__I (.I(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3016__A1 (.I(net1614));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3016__B2 (.I(net1547));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3016__C (.I(_1628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3020__I (.I(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3023__A1 (.I(_1632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3024__A1 (.I(net1560));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3024__B2 (.I(net1575));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3024__C (.I(_1636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3025__I (.I(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3026__I (.I(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3028__I (.I(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3029__I (.I(_0984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3031__B2 (.I(_1643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3032__A1 (.I(net1028));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3032__B2 (.I(net1618));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3033__I (.I(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3034__I (.I(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3036__I (.I(_0994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3037__I (.I(_0996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3039__A1 (.I(_1648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3040__B2 (.I(net1521));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3041__A1 (.I(net1778));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3041__A2 (.I(net1777));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3041__A3 (.I(_1645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3041__A4 (.I(net1776));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3042__I (.I(_1002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3043__I (.I(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3044__A2 (.I(_1655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3044__B1 (.I(_1656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3045__I (.I(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3046__I (.I(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3047__A1 (.I(net1427));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3048__I (.I(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3049__I (.I(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3051__I (.I(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3052__I (.I(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3053__A1 (.I(net1227));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3053__A2 (.I(_1664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3053__B2 (.I(net1375));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3054__A1 (.I(_1657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3054__A3 (.I(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3057__A1 (.I(net1135));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3057__B2 (.I(net922));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3058__I (.I(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3060__A1 (.I(net1148));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3060__B2 (.I(net935));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3061__I (.I(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3065__I (.I(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3067__A4 (.I(_1679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3068__A2 (.I(_1667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3068__A3 (.I(_1680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3069__A1 (.I(_1551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3070__I (.I(net1230));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3073__A1 (.I(net1322));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3078__A2 (.I(_1685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3078__A3 (.I(_1687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3079__I (.I(net1269));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3081__B2 (.I(_1692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3082__B2 (.I(net1243));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3085__A1 (.I(_1695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3086__C (.I(_1697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3087__I (.I(net1016));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3088__I (.I(net1002));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3090__C (.I(_1701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3091__A1 (.I(net1775));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3091__A2 (.I(net1774));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3091__A3 (.I(_1698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3092__A1 (.I(net1229));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3092__B2 (.I(net962));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3093__A1 (.I(net1442));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3093__B2 (.I(net989));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3096__A1 (.I(_1704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3096__A3 (.I(_1706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3096__A4 (.I(_1707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3097__B2 (.I(net1509));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3098__A1 (.I(net1650));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3098__B2 (.I(net1096));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3099__A1 (.I(net1189));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3099__B2 (.I(net1109));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3100__A1 (.I(net1162));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3101__A1 (.I(_1709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3101__A2 (.I(_1710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3102__A1 (.I(_1703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3102__A2 (.I(_1708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3106__A1 (.I(net1615));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3106__B2 (.I(net1548));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3106__C (.I(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3109__A1 (.I(_1719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3110__A1 (.I(net1561));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3110__B2 (.I(net1576));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3110__C (.I(_1721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3113__B2 (.I(_1724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3114__A1 (.I(net1029));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3114__B2 (.I(net1629));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3117__A1 (.I(_1727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3118__B2 (.I(net1522));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3119__A1 (.I(net1773));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3119__A2 (.I(net1772));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3119__A3 (.I(_1726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3119__A4 (.I(net1771));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3120__A2 (.I(_1655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3120__B1 (.I(_1656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3121__A1 (.I(net1428));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3123__A1 (.I(net1228));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3123__A2 (.I(_1664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3123__B2 (.I(net1376));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3124__A1 (.I(_1732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3125__A1 (.I(net1136));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3125__B2 (.I(net923));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3126__A1 (.I(net1149));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3126__B2 (.I(net936));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3129__A4 (.I(_1740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3130__A2 (.I(_1736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3130__A3 (.I(_1741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3131__A1 (.I(_1682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3131__B1 (.I(_1714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3132__I (.I(net1341));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3135__A1 (.I(net1323));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3137__I (.I(_0028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3141__A2 (.I(_1746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3141__A3 (.I(_1749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3142__I (.I(net1270));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3143__I (.I(net1257));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3145__B2 (.I(net1244));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3147__I (.I(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3149__A1 (.I(_1757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3150__B2 (.I(net1070));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3150__C (.I(_1760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3151__I (.I(net1017));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3152__I (.I(net1003));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3154__C (.I(_1764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3155__A1 (.I(_1752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3155__A2 (.I(_1756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3155__A3 (.I(_1761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3155__A4 (.I(_1765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3156__A1 (.I(net1241));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3156__B2 (.I(net964));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3157__A1 (.I(net1443));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3157__B2 (.I(net990));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3160__A1 (.I(_1767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3160__A3 (.I(_1769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3160__A4 (.I(_1770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3161__B2 (.I(net1510));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3162__A1 (.I(net1651));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3162__B2 (.I(net1107));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3163__A1 (.I(net1190));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3163__B2 (.I(net1110));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3165__A1 (.I(net1164));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3166__A1 (.I(_1772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3166__A2 (.I(_1773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3167__A2 (.I(_1771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3171__A1 (.I(net1616));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3171__B2 (.I(net1549));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3171__C (.I(_1781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3175__A1 (.I(_1783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3176__A1 (.I(net1564));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3176__B2 (.I(net1577));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3176__C (.I(_1786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3179__B2 (.I(_1789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3180__A1 (.I(net1031));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3180__B2 (.I(net1638));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3183__A1 (.I(_1792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3184__B2 (.I(net1523));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3185__A1 (.I(net1770));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3185__A2 (.I(net1769));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3185__A3 (.I(_1791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3185__A4 (.I(net1768));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3186__A2 (.I(_1655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3186__B1 (.I(_1656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3187__A1 (.I(net1430));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3189__A1 (.I(net1231));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3189__A2 (.I(_1664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3189__B2 (.I(net1377));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3190__A1 (.I(_1797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3191__A1 (.I(net1137));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3191__B2 (.I(net924));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3192__A1 (.I(net1150));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3192__B2 (.I(net937));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3195__A4 (.I(_1805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3196__A2 (.I(_1801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3196__A3 (.I(_1806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3197__B1 (.I(_1778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3198__I (.I(net1452));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3200__A1 (.I(_1809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3201__A1 (.I(net1324));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3206__A2 (.I(_1811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3206__A3 (.I(_1813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3206__A4 (.I(_1815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3207__I (.I(net1271));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3208__I (.I(net1258));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3210__B2 (.I(net1245));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3210__C (.I(_1819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3213__A1 (.I(_1821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3214__C (.I(_1823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3215__I (.I(net1018));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3216__I (.I(net1004));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3218__A1 (.I(net1098));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3218__C (.I(_1827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3219__A1 (.I(_1816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3219__A2 (.I(_1820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3219__A3 (.I(_1824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3219__A4 (.I(_1828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3220__A1 (.I(net1252));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3220__B2 (.I(net965));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3221__A1 (.I(net1444));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3221__B2 (.I(net991));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3224__A1 (.I(_1830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3224__A3 (.I(_1832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3224__A4 (.I(_1833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3225__B2 (.I(net1511));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3226__A1 (.I(net1652));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3226__B2 (.I(net1118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3227__A1 (.I(net1191));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3227__B2 (.I(net1111));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3228__A1 (.I(net1165));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3229__A1 (.I(_1835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3229__A2 (.I(_1836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3230__A2 (.I(_1834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3234__A1 (.I(net1617));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3234__B2 (.I(net1550));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3234__C (.I(_1843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3237__A1 (.I(_1845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3238__A1 (.I(net1565));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3238__B2 (.I(net1578));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3238__C (.I(_1847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3241__B2 (.I(_1850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3242__A1 (.I(net1032));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3242__B2 (.I(net1639));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3242__C (.I(_1851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3245__A1 (.I(_1853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3246__B2 (.I(net1524));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3247__A1 (.I(net1767));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3247__A2 (.I(net1766));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3247__A3 (.I(_1852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3247__A4 (.I(net1765));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3248__A2 (.I(_1655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3248__B1 (.I(_1656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3249__A1 (.I(net1431));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3251__A1 (.I(net1232));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3251__A2 (.I(_1664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3251__B2 (.I(net1378));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3252__A1 (.I(_1858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3253__A1 (.I(net1138));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3253__B2 (.I(net925));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3254__A1 (.I(net1151));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3254__B2 (.I(net938));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3257__A4 (.I(_1866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3258__A2 (.I(_1862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3258__A3 (.I(_1867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3260__I (.I(net1563));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3261__I (.I(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3263__I (.I(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3264__I (.I(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3265__A3 (.I(_1873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3266__I (.I(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3267__I (.I(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3268__A1 (.I(net1325));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3270__I (.I(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3273__I (.I(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3274__I (.I(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3276__A2 (.I(_1877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3276__A3 (.I(_1880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3277__I (.I(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3278__I (.I(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3279__I (.I(net1272));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3280__I (.I(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3281__I (.I(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3282__I (.I(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3289__I (.I(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3290__I (.I(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3292__A1 (.I(_1897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3293__A2 (.I(_1895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3293__B1 (.I(_1896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3293__C (.I(_1901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3294__I (.I(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3295__I (.I(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3296__I (.I(net1020));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3297__I (.I(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3298__I (.I(_0102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3299__I (.I(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3300__I (.I(net1005));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3302__C (.I(_1910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3303__A1 (.I(_1885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3303__A2 (.I(_1894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3303__A3 (.I(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3303__A4 (.I(_1911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3304__I (.I(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3305__I (.I(_0912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3306__A1 (.I(net1263));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3307__I (.I(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3308__I (.I(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3309__A1 (.I(net1445));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3309__B2 (.I(net992));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3316__A1 (.I(_1915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3316__A3 (.I(_1921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3316__A4 (.I(_1924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3317__I (.I(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3318__I (.I(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3319__B2 (.I(net1512));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3320__I (.I(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3321__I (.I(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3322__B2 (.I(net1130));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3323__I (.I(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3324__I (.I(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3325__A1 (.I(net1192));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3325__B2 (.I(net1112));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3326__I (.I(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3328__A2 (.I(_1931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3329__A3 (.I(_1937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3330__I (.I(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3331__I (.I(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3333__I (.I(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3334__I (.I(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3335__I (.I(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3338__A1 (.I(net1619));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3338__B2 (.I(net1552));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3338__C (.I(_1946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3342__I (.I(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3345__A1 (.I(_1950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3346__A1 (.I(net1566));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3346__B2 (.I(net1579));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3346__C (.I(_1954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3347__I (.I(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3348__I (.I(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3350__I (.I(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3351__I (.I(_0984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3353__B2 (.I(_1961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3354__A2 (.I(_1956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3354__B1 (.I(_1957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3354__B2 (.I(net1640));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3355__I (.I(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3356__I (.I(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3357__I (.I(net996));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3358__I (.I(_0994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3359__I (.I(_0996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3361__A1 (.I(_1966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3362__B2 (.I(net1525));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3363__A1 (.I(net1764));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3363__A2 (.I(net1763));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3363__A3 (.I(_1963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3363__A4 (.I(net1762));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3364__I (.I(_1002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3365__I (.I(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3367__I (.I(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3368__I (.I(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3369__A1 (.I(net1432));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3370__I (.I(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3371__I (.I(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3373__I (.I(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3374__I (.I(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3375__A1 (.I(net1233));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3375__B2 (.I(net1379));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3376__A1 (.I(_1975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3379__A1 (.I(net1139));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3379__A2 (.I(_1986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3379__B1 (.I(_1987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3380__I (.I(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3382__A1 (.I(net1153));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3382__B1 (.I(_1990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3383__I (.I(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3385__B1 (.I(_1993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3387__I (.I(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3389__A4 (.I(_1997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3390__A2 (.I(_1985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3390__A3 (.I(_1998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3391__A2 (.I(_1870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3391__B1 (.I(_1938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3392__I (.I(net1642));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3394__A3 (.I(_1873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3395__A1 (.I(net1326));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3400__A2 (.I(_2003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3400__A3 (.I(_2005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3401__I (.I(net1273));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3402__I (.I(net1260));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3406__I (.I(net1206));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3407__A1 (.I(_2013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3408__A2 (.I(_1895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3408__B1 (.I(_1896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3408__C (.I(_2015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3409__I (.I(net1021));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3410__I (.I(net1006));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3412__C (.I(_2019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3413__A1 (.I(_2008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3413__A2 (.I(_2012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3413__A3 (.I(_2016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3413__A4 (.I(_2020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3414__A1 (.I(net1274));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3415__A1 (.I(net1446));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3415__B2 (.I(net993));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3418__A1 (.I(_2022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3418__A3 (.I(_2024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3418__A4 (.I(_2025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3419__B2 (.I(net1513));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3420__B2 (.I(net1141));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3421__A1 (.I(net1193));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3421__B2 (.I(net1113));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3423__A2 (.I(_2028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3424__A2 (.I(_2026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3424__A3 (.I(_2031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3428__A1 (.I(net1620));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3428__B2 (.I(net1553));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3428__C (.I(_2035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3431__A1 (.I(_2037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3432__A1 (.I(net1567));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3432__B2 (.I(net1580));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3432__C (.I(_2039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3435__B2 (.I(_2042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3436__A2 (.I(_1956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3436__B1 (.I(_1957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3436__B2 (.I(net1641));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3437__I (.I(net1007));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3440__B2 (.I(net1526));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3441__A1 (.I(net1761));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3441__A2 (.I(net1760));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3441__A3 (.I(_2044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3441__A4 (.I(net1759));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3443__A1 (.I(net1433));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3445__A1 (.I(net1234));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3445__B2 (.I(net1380));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3446__A1 (.I(_2050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3446__A3 (.I(_2052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3447__A1 (.I(net1140));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3447__A2 (.I(_1986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3447__B1 (.I(_1987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3448__A1 (.I(net1154));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3448__B1 (.I(_1990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3449__B1 (.I(_1993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3451__A4 (.I(_2058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3452__A2 (.I(_2054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3452__A3 (.I(_2059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3453__A2 (.I(_1870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3453__B1 (.I(_2032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3454__I (.I(net1653));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3456__A3 (.I(_1873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3457__A1 (.I(net1327));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3459__I (.I(_0028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3463__A2 (.I(_2064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3463__A3 (.I(_2067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3464__I (.I(net1275));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3465__I (.I(net1261));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3469__I (.I(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3470__I (.I(net1208));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3471__A1 (.I(_2075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3471__A2 (.I(_2076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3472__A2 (.I(_1895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3472__B1 (.I(_1896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3472__C (.I(_2078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3473__I (.I(net1022));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3474__I (.I(net1009));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3476__C (.I(_2082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3477__A1 (.I(_2070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3477__A2 (.I(_2074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3477__A3 (.I(_2079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3477__A4 (.I(_2083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3478__A1 (.I(net1285));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3479__A1 (.I(net1447));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3479__B2 (.I(net994));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3482__A1 (.I(_2085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3482__A3 (.I(_2087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3482__A4 (.I(_2088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3483__B2 (.I(net1514));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3484__B2 (.I(net1152));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3485__A1 (.I(net1194));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3485__B2 (.I(net1114));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3487__B (.I(_2093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3488__A2 (.I(_2091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3489__A3 (.I(_2095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3493__A1 (.I(net1621));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3493__B2 (.I(net1554));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3493__C (.I(_2099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3497__A1 (.I(_2101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3498__A1 (.I(net1568));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3498__B2 (.I(net1581));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3498__C (.I(_2104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3501__B2 (.I(_2107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3502__A2 (.I(_1956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3502__B1 (.I(_1957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3502__B2 (.I(net1643));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3503__I (.I(net1019));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3504__I (.I(net1418));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3506__B2 (.I(net1527));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3507__A1 (.I(net1758));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3507__A2 (.I(net1757));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3507__A3 (.I(_2109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3507__A4 (.I(net1756));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3509__A1 (.I(net1434));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3511__A1 (.I(net1235));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3511__B2 (.I(net1381));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3512__A1 (.I(_2115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3512__A3 (.I(_2117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3513__A1 (.I(net1142));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3513__A2 (.I(_1986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3513__B1 (.I(_1987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3514__A1 (.I(net1155));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3514__B1 (.I(_1990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3515__B1 (.I(_1993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3517__A4 (.I(_2123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3518__A2 (.I(_2119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3518__A3 (.I(_2124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3519__A2 (.I(_1870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3519__B1 (.I(_2096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3520__I (.I(net1664));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3522__A3 (.I(_1873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3523__A1 (.I(net1328));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3528__A2 (.I(_2129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3528__A3 (.I(_2131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3529__I (.I(net1276));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3531__B2 (.I(_2136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3534__I (.I(net1209));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3535__A1 (.I(_2139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3535__A2 (.I(_2076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3536__A2 (.I(_1895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3536__B1 (.I(_1896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3536__C (.I(_2141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3537__I (.I(net1023));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3538__I (.I(net1010));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3540__C (.I(_2145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3541__A1 (.I(_2134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3541__A2 (.I(_2138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3541__A3 (.I(_2142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3541__A4 (.I(_2146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3542__A1 (.I(net1296));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3543__A1 (.I(net1448));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3543__B2 (.I(net995));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3546__A1 (.I(_2148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3546__A3 (.I(_2150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3546__A4 (.I(_2151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3547__B2 (.I(net1515));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3548__B2 (.I(net1163));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3549__A1 (.I(net1195));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3549__B2 (.I(net1115));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3550__B (.I(_2093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3551__A2 (.I(_2154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3552__A3 (.I(_2157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3556__A1 (.I(net1622));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3556__B2 (.I(net1555));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3556__C (.I(_2161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3559__A1 (.I(_2163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3560__A1 (.I(net1569));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3560__B2 (.I(net1582));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3560__C (.I(_2165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3563__B2 (.I(_2168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3564__A1 (.I(net1036));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3564__A2 (.I(_1956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3564__B1 (.I(_1957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3564__B2 (.I(net1644));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3565__I (.I(net1030));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3568__B2 (.I(net1528));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3569__A1 (.I(net1755));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3569__A2 (.I(net1754));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3569__A3 (.I(_2170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3569__A4 (.I(net1753));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3571__A1 (.I(net1435));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3573__A1 (.I(net1236));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3573__B2 (.I(net1382));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3574__A1 (.I(_2176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3574__A3 (.I(_2178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3575__A1 (.I(net1143));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3575__A2 (.I(_1986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3575__B1 (.I(_1987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3576__A1 (.I(net1156));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3576__B1 (.I(_1990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3577__B1 (.I(_1993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3579__A3 (.I(_2183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3579__A4 (.I(_2184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3580__A2 (.I(_2180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3580__A3 (.I(_2185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3581__A2 (.I(_1870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3581__B1 (.I(_2158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3582__I (.I(net908));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3583__I (.I(net1316));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3584__A2 (.I(_0023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3584__A3 (.I(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3585__A1 (.I(net1330));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3585__A2 (.I(_0033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3585__A3 (.I(_0040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3586__I (.I(net1397));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3587__A2 (.I(_0051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3588__I (.I(net1303));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3589__A1 (.I(_2193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3589__A2 (.I(_0060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3589__A3 (.I(_0054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3591__I (.I(net1277));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3592__I (.I(net1264));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3593__A2 (.I(_0077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3593__A3 (.I(_0062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3593__B1 (.I(_0084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3594__A1 (.I(net1223));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3594__B2 (.I(net1250));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3596__I (.I(net1210));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3597__A1 (.I(_2200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3597__A2 (.I(_2076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3597__A3 (.I(_0105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3597__B1 (.I(_0111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3598__A2 (.I(_0092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3598__B1 (.I(_0099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3598__C (.I(net1828));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3599__I (.I(net1024));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3600__I (.I(net1011));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3601__A3 (.I(_0103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3602__A1 (.I(net1103));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3602__B2 (.I(net1090));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3603__A1 (.I(_2195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3603__A2 (.I(_2199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3603__A3 (.I(_2203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3603__A4 (.I(_2207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3604__A1 (.I(net1307));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3604__A2 (.I(_0138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3604__B1 (.I(_0142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3605__A1 (.I(net1449));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3605__A2 (.I(_0148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3605__B1 (.I(_0153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3605__B2 (.I(net997));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3606__A2 (.I(_0157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3606__B1 (.I(_0162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3607__A2 (.I(_0166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3607__B1 (.I(_0169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3608__A1 (.I(net1822));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3608__A4 (.I(_2212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3609__A2 (.I(_0175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3609__B1 (.I(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3609__B2 (.I(net1516));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3610__A1 (.I(net1658));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3610__A2 (.I(_0182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3610__B1 (.I(_0185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3610__B2 (.I(net1174));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3611__A1 (.I(net1197));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3611__A2 (.I(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3611__B1 (.I(_0196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3611__B2 (.I(net1116));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3612__A1 (.I(net1170));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3612__A2 (.I(_0201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3612__B (.I(_2093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3613__A1 (.I(_2214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3613__A2 (.I(_2215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3614__A2 (.I(_2213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3615__I (.I(net1610));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3616__A1 (.I(net1636));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3616__A2 (.I(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3616__A3 (.I(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3617__A2 (.I(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3618__A1 (.I(net1623));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3618__A2 (.I(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3618__B1 (.I(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3618__B2 (.I(net1556));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3620__I (.I(net1597));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3621__A1 (.I(_2224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3621__A2 (.I(_0235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3621__B1 (.I(_0240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3622__A2 (.I(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3622__B1 (.I(_0232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3622__B2 (.I(net1583));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3622__C (.I(_2226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3625__A2 (.I(_0253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3625__B1 (.I(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3625__B2 (.I(_2229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3626__A1 (.I(net1037));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3626__A2 (.I(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3626__B1 (.I(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3626__B2 (.I(net1645));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3626__C (.I(_2230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3628__I (.I(net1440));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3629__A1 (.I(_2232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3629__A2 (.I(_0269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3629__B1 (.I(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3630__A1 (.I(net1574));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3630__B2 (.I(net1530));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3630__C (.I(_2234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3631__A1 (.I(net1821));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3631__A2 (.I(net1820));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3631__A3 (.I(_2231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3631__A4 (.I(net1819));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3632__A2 (.I(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3632__B1 (.I(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3633__A1 (.I(net1436));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3633__A2 (.I(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3633__B1 (.I(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3633__B2 (.I(net1344));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3634__A1 (.I(net1357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3634__A2 (.I(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3634__B1 (.I(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3635__A1 (.I(net1237));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3635__A2 (.I(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3635__B1 (.I(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3635__B2 (.I(net1383));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3636__A1 (.I(_2237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3636__A2 (.I(_2238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3637__A1 (.I(net1144));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3637__A2 (.I(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3637__B1 (.I(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3637__B2 (.I(net931));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3638__A1 (.I(net1157));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3638__A2 (.I(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3638__B1 (.I(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3639__A1 (.I(net904));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3639__A2 (.I(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3639__B1 (.I(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3639__B2 (.I(net917));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3641__A4 (.I(_2245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3642__A2 (.I(_2241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3642__A3 (.I(_2246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3643__A2 (.I(_0014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3643__B1 (.I(_2219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3644__I (.I(net919));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3645__I (.I(net1317));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3646__A2 (.I(_0023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3646__A3 (.I(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3647__A1 (.I(net1331));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3647__A2 (.I(_0033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3647__A3 (.I(_0040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3648__I (.I(net1398));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3649__A2 (.I(_0051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3650__I (.I(net1304));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3651__A1 (.I(_2254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3651__A2 (.I(_0060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3651__A3 (.I(_0054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3653__I (.I(net1278));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3654__I (.I(net1265));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3655__A2 (.I(_0077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3655__A3 (.I(_0062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3655__B1 (.I(_0084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3656__A1 (.I(net1224));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3656__B2 (.I(net1251));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3658__I (.I(net1211));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3659__A1 (.I(_2261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3659__A2 (.I(_2076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3659__A3 (.I(_0105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3659__B1 (.I(_0111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3660__A2 (.I(_0092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3660__B1 (.I(_0099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3660__C (.I(net1827));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3661__I (.I(net1025));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3662__I (.I(net1012));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3663__A3 (.I(_0103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3664__A1 (.I(net1104));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3664__B2 (.I(net1091));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3664__C (.I(_2267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3665__A1 (.I(_2256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3665__A2 (.I(_2260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3665__A3 (.I(_2264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3665__A4 (.I(_2268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3666__A1 (.I(net1318));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3666__A2 (.I(_0138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3666__B1 (.I(_0142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3667__A1 (.I(net1450));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3667__A2 (.I(_0148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3667__B1 (.I(_0153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3667__B2 (.I(net998));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3668__A2 (.I(_0157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3668__B1 (.I(_0162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3669__A2 (.I(_0166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3669__B1 (.I(_0169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3670__A1 (.I(net1818));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3670__A4 (.I(_2273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3671__A2 (.I(_0175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3671__B1 (.I(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3671__B2 (.I(net1517));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3672__A1 (.I(net1659));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3672__A2 (.I(_0182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3672__B1 (.I(_0185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3672__B2 (.I(net1185));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3673__A1 (.I(net1198));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3673__A2 (.I(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3673__B1 (.I(_0196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3673__B2 (.I(net1117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3674__A1 (.I(net1171));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3674__A2 (.I(_0201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3674__B (.I(_2093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3675__A1 (.I(_2275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3675__A2 (.I(_2276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3676__A2 (.I(_2274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3677__I (.I(net1611));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3678__A1 (.I(net1637));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3678__A2 (.I(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3678__A3 (.I(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3679__A2 (.I(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3680__A1 (.I(net1624));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3680__A2 (.I(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3680__B1 (.I(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3680__B2 (.I(net1557));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3681__I (.I(net1291));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3682__I (.I(net1598));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3683__A1 (.I(_2285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3683__A2 (.I(_0235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3683__B1 (.I(_0240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3684__A2 (.I(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3684__B1 (.I(_0232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3684__B2 (.I(net1584));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3684__C (.I(_2287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3687__A2 (.I(_0253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3687__B1 (.I(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3687__B2 (.I(_2290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3688__A1 (.I(net1038));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3688__A2 (.I(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3688__B1 (.I(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3688__B2 (.I(net1646));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3688__C (.I(_2291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3690__I (.I(net1451));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3691__A1 (.I(_2293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3691__A2 (.I(_0269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3691__B1 (.I(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3692__A1 (.I(net1585));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3692__B2 (.I(net1531));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3692__C (.I(_2295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3693__A1 (.I(net1817));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3693__A2 (.I(net1816));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3693__A3 (.I(_2292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3693__A4 (.I(net1815));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3694__A2 (.I(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3694__B1 (.I(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3695__A1 (.I(net1437));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3695__A2 (.I(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3695__B1 (.I(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3695__B2 (.I(net1345));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3696__A1 (.I(net1358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3696__A2 (.I(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3696__B1 (.I(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3697__A1 (.I(net1238));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3697__A2 (.I(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3697__B1 (.I(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3697__B2 (.I(net1384));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3698__A1 (.I(_2298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3698__A2 (.I(_2299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3699__A1 (.I(net1145));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3699__A2 (.I(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3699__B1 (.I(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3700__A1 (.I(net1158));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3700__A2 (.I(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3700__B1 (.I(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3701__A1 (.I(net905));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3701__A2 (.I(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3701__B1 (.I(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3701__B2 (.I(net918));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3703__A4 (.I(_2306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3704__A2 (.I(_2302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3704__A3 (.I(_2307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3705__A2 (.I(_0014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3707__I (.I(net1666));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3708__A1 (.I(net1665));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3710__A1 (.I(net1668));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3710__A2 (.I(net1667));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3712__A1 (.I(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3712__A2 (.I(_0005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3713__I (.I(net1670));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3714__I (.I(net1669));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3716__I (.I(_0009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3717__A1 (.I(_0006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3717__A2 (.I(_0010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3719__I (.I(_0012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3720__I (.I(_0013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3721__I (.I(_0014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3722__I (.I(net496));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3723__I (.I(net1668));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3725__I (.I(net1667));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3726__A1 (.I(net1665));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3727__A1 (.I(_0018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3727__A2 (.I(_0019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3727__A3 (.I(_0020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3728__I (.I(_0021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3729__I (.I(_0022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3730__I (.I(_0023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3731__A1 (.I(net1670));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3733__I (.I(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3734__I (.I(_0027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3735__I (.I(_0028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3736__A1 (.I(_0016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3737__I (.I(net1669));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3739__I (.I(_0032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3740__I (.I(_0033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3741__I (.I(net1668));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3742__I (.I(net1667));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3745__A3 (.I(_0038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3746__I (.I(_0039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3747__I (.I(_0040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3748__A1 (.I(net512));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3749__I (.I(net590));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3750__I (.I(net1665));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3752__I (.I(net1666));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3756__A1 (.I(_0045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3756__A2 (.I(_0047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3756__A3 (.I(_0049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3757__I (.I(_0050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3758__I (.I(_0051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3759__I (.I(_0027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3761__A3 (.I(_0054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3762__I (.I(net481));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3765__A1 (.I(_0018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3765__A2 (.I(_0019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3766__I (.I(_0059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3767__I (.I(_0060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3768__I (.I(_0027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3769__I (.I(_0062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3771__A3 (.I(_0055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3771__A4 (.I(_0064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3773__A1 (.I(_0006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3773__A2 (.I(_0066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3777__A3 (.I(_0070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3778__A1 (.I(_0071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3778__A2 (.I(_0066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3781__I (.I(net450));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3782__A1 (.I(_0018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3782__A2 (.I(_0019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3783__I (.I(_0076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3784__I (.I(_0077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3785__I (.I(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3786__I (.I(_0079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3787__I (.I(net1670));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3788__I (.I(_0020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3789__A3 (.I(_0070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3790__I (.I(_0083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3791__I (.I(_0084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3792__I (.I(net434));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3793__B2 (.I(_0086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3794__A1 (.I(net387));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3794__B2 (.I(net418));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3795__A2 (.I(net1669));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3796__I (.I(_0089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3797__A1 (.I(_0090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3797__A2 (.I(_0076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3799__I (.I(_0092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3802__I (.I(_0089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3804__A1 (.I(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3804__A2 (.I(_0097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3806__I (.I(_0099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3809__I (.I(_0102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3811__I (.I(_0104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3812__I (.I(_0105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3815__A1 (.I(net1668));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3815__A3 (.I(net1665));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3816__A3 (.I(_0109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3817__I (.I(_0110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3818__I (.I(_0111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3819__I (.I(net372));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3820__A1 (.I(_0101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3820__A2 (.I(_0103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3820__B2 (.I(_0113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3821__B2 (.I(net216));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3821__C (.I(_0114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3822__A1 (.I(_0021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3822__A2 (.I(_0090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3825__I (.I(_0059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3826__A1 (.I(_0090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3826__A2 (.I(_0119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3829__I (.I(net154));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3830__A1 (.I(_0045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3830__A2 (.I(_0047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3830__A3 (.I(_0070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3831__I (.I(_0124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3833__I (.I(_0090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3834__I (.I(_0127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3835__A3 (.I(_0038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3835__A4 (.I(_0070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3836__I (.I(_0129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3838__I (.I(net139));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3840__A1 (.I(net248));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3840__A2 (.I(_0118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3840__B1 (.I(_0122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3840__B2 (.I(net232));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3840__C (.I(_0133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3841__A1 (.I(_0065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3841__A2 (.I(_0088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3841__A3 (.I(_0115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3841__A4 (.I(_0134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3842__A1 (.I(_0005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3843__A1 (.I(_0010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3843__A2 (.I(_0136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3845__I (.I(_0138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3846__I (.I(_0009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3847__A1 (.I(_0140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3847__A2 (.I(_0050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3849__I (.I(_0142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3850__A1 (.I(net367));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3850__B2 (.I(net92));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3851__A2 (.I(net1669));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3853__A1 (.I(_0146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3853__A2 (.I(_0124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3854__I (.I(_0147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3855__I (.I(_0148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3857__I (.I(_0109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3858__A1 (.I(_0150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3858__A2 (.I(_0151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3859__I (.I(_0152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3860__I (.I(_0153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3861__A1 (.I(net651));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3861__B2 (.I(net124));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3862__A1 (.I(_0146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3862__A2 (.I(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3864__I (.I(_0157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3866__I (.I(_0159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3867__A1 (.I(_0160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3867__A2 (.I(_0076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3869__I (.I(_0162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3871__A1 (.I(_0146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3871__A2 (.I(_0071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3873__I (.I(_0166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3874__A1 (.I(_0136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3874__A2 (.I(_0160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3876__I (.I(_0169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3878__A1 (.I(net1752));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3878__A4 (.I(_0171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3880__A1 (.I(_0050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3880__A2 (.I(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3882__I (.I(_0175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3883__A1 (.I(_0160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3883__A2 (.I(_0119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3884__I (.I(_0177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3885__I (.I(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3886__B2 (.I(net729));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3887__A1 (.I(_0140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3887__A2 (.I(_0022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3889__I (.I(_0182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3890__A1 (.I(_0140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3890__A2 (.I(_0071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3892__I (.I(_0185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3893__A1 (.I(net894));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3893__B2 (.I(net211));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3895__A3 (.I(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3896__I (.I(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3897__I (.I(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3900__A3 (.I(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3901__A1 (.I(_0097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3901__A2 (.I(_0194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3902__I (.I(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3903__I (.I(_0196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3904__A1 (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3904__B2 (.I(net263));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3905__A1 (.I(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3905__A2 (.I(_0049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3906__A1 (.I(_0097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3906__A2 (.I(_0199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3908__I (.I(_0201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3909__A1 (.I(net325));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3909__B (.I(_0013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3910__A1 (.I(_0180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3910__A2 (.I(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3911__A2 (.I(_0172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3913__I (.I(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3914__A1 (.I(_0207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3914__A2 (.I(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3916__I (.I(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3917__I (.I(_0104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3918__A1 (.I(_0146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3918__A2 (.I(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3919__I (.I(_0212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3920__I (.I(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3922__A1 (.I(_0045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3922__A2 (.I(_0047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3922__A3 (.I(_0049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3922__A4 (.I(_0207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3923__I (.I(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3924__I (.I(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3925__I (.I(_0207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3926__I (.I(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3927__I (.I(_0151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3928__I (.I(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3931__A1 (.I(net853));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3931__B2 (.I(net775));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3931__C (.I(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3933__A1 (.I(_0159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3933__A2 (.I(_0226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3934__I (.I(_0227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3935__I (.I(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3937__A1 (.I(_0159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3937__A2 (.I(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3938__I (.I(_0231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3939__I (.I(_0232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3940__I (.I(net465));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3942__I (.I(_0235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3943__I (.I(_0066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3944__I (.I(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3945__A1 (.I(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3945__A2 (.I(_0049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3945__A3 (.I(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3947__I (.I(_0240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3948__I (.I(net823));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3949__A1 (.I(_0234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3949__A3 (.I(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3950__A1 (.I(net792));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3950__B2 (.I(net807));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3951__A1 (.I(_0071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3951__A2 (.I(_0097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3953__I (.I(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3954__A1 (.I(_0010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3954__A2 (.I(_0119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3956__I (.I(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3958__A3 (.I(_0005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3959__I (.I(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3960__I (.I(_0253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3961__A3 (.I(_0038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3961__A4 (.I(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3962__I (.I(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3963__I (.I(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3965__B2 (.I(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3966__A1 (.I(net170));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3966__B2 (.I(net833));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3966__C (.I(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3967__A1 (.I(_0010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3967__A2 (.I(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3968__I (.I(_0261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3970__A1 (.I(_0159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3970__A2 (.I(_0022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3971__I (.I(_0264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3974__A1 (.I(_0045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3974__A2 (.I(_0047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3974__A3 (.I(_0005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3974__A4 (.I(_0150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3975__I (.I(_0268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3976__I (.I(_0269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3977__A1 (.I(_0018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3977__A2 (.I(_0019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3977__A3 (.I(_0038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3977__A4 (.I(_0150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3978__I (.I(_0271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3979__I (.I(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3981__A1 (.I(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3982__B2 (.I(net745));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3983__A1 (.I(net1750));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3983__A2 (.I(net1748));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3983__A4 (.I(net1747));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3984__A1 (.I(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3984__A2 (.I(_0032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3986__I (.I(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3987__A1 (.I(_0151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3987__A2 (.I(_0032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3989__I (.I(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3991__A1 (.I(_0006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3991__A2 (.I(_0160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3993__I (.I(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3994__I (.I(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3995__A1 (.I(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3995__A2 (.I(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3997__I (.I(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3998__A1 (.I(net636));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3999__I (.I(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4000__A1 (.I(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4000__A2 (.I(_0226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4002__I (.I(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4003__A1 (.I(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4003__A2 (.I(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4005__I (.I(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4007__A1 (.I(_0124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4007__A2 (.I(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4009__I (.I(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4010__A1 (.I(_0199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4010__A2 (.I(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4012__I (.I(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4013__A1 (.I(net403));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4013__B2 (.I(net574));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4014__A1 (.I(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4015__A1 (.I(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4015__A2 (.I(_0226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4017__I (.I(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4018__I (.I(_0009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4019__A1 (.I(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4019__A2 (.I(_0226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4021__I (.I(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4022__A1 (.I(net294));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4023__A1 (.I(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4023__A2 (.I(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4025__I (.I(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4026__A1 (.I(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4026__A2 (.I(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4028__I (.I(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4029__A1 (.I(net309));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4030__A1 (.I(_0140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4030__A2 (.I(_0194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4032__I (.I(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4033__A1 (.I(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4033__A2 (.I(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4035__I (.I(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4037__A1 (.I(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4037__A2 (.I(_0199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4040__A1 (.I(_0150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4040__A2 (.I(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4041__I (.I(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4044__A4 (.I(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4045__A1 (.I(_0277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4045__A2 (.I(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4046__B1 (.I(_0205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4046__B2 (.I(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4048__I (.I(net497));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4049__A1 (.I(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4050__A1 (.I(net513));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4051__I (.I(net591));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4052__A3 (.I(_0054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4053__I (.I(net482));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4055__A3 (.I(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4056__I (.I(net451));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4057__I (.I(net435));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4059__A1 (.I(net388));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4059__B2 (.I(net419));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4061__I (.I(net373));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4062__A1 (.I(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4062__A2 (.I(_0103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4062__B2 (.I(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4063__C (.I(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4064__I (.I(net155));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4065__I (.I(net140));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4067__A1 (.I(net249));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4067__A2 (.I(_0118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4067__B1 (.I(_0122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4067__B2 (.I(net233));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4068__A1 (.I(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4068__A2 (.I(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4068__A3 (.I(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4068__A4 (.I(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4069__A1 (.I(net378));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4069__B2 (.I(net93));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4070__A1 (.I(net652));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4070__B2 (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4073__A1 (.I(net1746));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4073__A3 (.I(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4073__A4 (.I(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4074__B2 (.I(net730));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4075__A1 (.I(net895));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4075__B2 (.I(net222));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4076__A1 (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4076__B2 (.I(net264));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4077__A1 (.I(net326));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4077__B (.I(_0013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4078__A1 (.I(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4078__A2 (.I(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4079__A2 (.I(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4083__A1 (.I(net854));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4083__B2 (.I(net776));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4083__C (.I(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4084__I (.I(net466));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4085__I (.I(net824));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4086__A1 (.I(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4086__A3 (.I(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4087__A1 (.I(net793));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4087__B2 (.I(net808));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4087__C (.I(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4090__B2 (.I(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4091__A1 (.I(net171));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4091__B2 (.I(net844));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4091__C (.I(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4094__A1 (.I(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4095__B2 (.I(net746));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4096__A1 (.I(net1744));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4096__A2 (.I(net1742));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4096__A4 (.I(net1741));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4098__A1 (.I(net637));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4100__A1 (.I(net404));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4100__B2 (.I(net575));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4101__A1 (.I(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4102__A1 (.I(net295));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4103__A1 (.I(net310));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4106__A2 (.I(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4106__A4 (.I(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4107__A1 (.I(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4107__A2 (.I(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4108__B1 (.I(net1703));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4108__B2 (.I(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4110__I (.I(net498));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4111__A1 (.I(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4112__A1 (.I(net514));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4113__I (.I(net592));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4116__I (.I(net483));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4118__A3 (.I(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4118__A4 (.I(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4119__I (.I(net452));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4120__I (.I(net436));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4122__A1 (.I(net390));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4122__B2 (.I(net420));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4124__I (.I(_0102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4125__I (.I(net374));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4127__C (.I(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4128__I (.I(net157));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4129__I (.I(net141));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4131__A1 (.I(net250));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4131__A2 (.I(_0118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4131__B1 (.I(_0122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4131__B2 (.I(net235));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4132__A1 (.I(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4132__A2 (.I(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4132__A3 (.I(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4132__A4 (.I(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4133__A1 (.I(net389));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4133__B2 (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4134__A1 (.I(net653));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4134__B2 (.I(net126));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4137__A1 (.I(net1740));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4137__A3 (.I(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4137__A4 (.I(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4138__B2 (.I(net731));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4139__A1 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4139__B2 (.I(net234));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4140__A1 (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4140__B2 (.I(net265));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4141__I (.I(_0012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4142__A1 (.I(net327));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4143__A1 (.I(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4143__A2 (.I(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4144__A2 (.I(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4148__A1 (.I(net856));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4148__B2 (.I(net779));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4148__C (.I(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4149__I (.I(net468));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4150__I (.I(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4151__I (.I(net825));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4152__A1 (.I(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4152__A3 (.I(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4153__A1 (.I(net794));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4153__B2 (.I(net809));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4153__C (.I(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4156__B2 (.I(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4157__A1 (.I(net172));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4157__B2 (.I(net855));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4160__A1 (.I(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4161__B2 (.I(net747));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4162__A1 (.I(net1738));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4162__A2 (.I(net1736));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4162__A4 (.I(net1735));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4164__A1 (.I(net638));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4166__A1 (.I(net405));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4166__B2 (.I(net576));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4167__A1 (.I(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4168__A1 (.I(net296));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4169__A1 (.I(net312));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4172__A4 (.I(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4173__A1 (.I(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4173__A2 (.I(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4174__B1 (.I(net1702));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4174__B2 (.I(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4176__I (.I(net499));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4177__A1 (.I(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4178__A1 (.I(net515));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4179__I (.I(net593));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4181__I (.I(net484));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4183__A3 (.I(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4183__A4 (.I(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4184__I (.I(net453));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4186__B2 (.I(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4187__A1 (.I(net391));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4187__B2 (.I(net421));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4189__I (.I(net375));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4190__A1 (.I(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4191__C (.I(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4192__I (.I(net158));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4193__I (.I(net142));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4195__A1 (.I(net251));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4195__A2 (.I(_0118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4195__B1 (.I(_0122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4195__B2 (.I(net236));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4195__C (.I(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4196__A1 (.I(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4196__A2 (.I(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4196__A3 (.I(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4196__A4 (.I(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4197__A1 (.I(net400));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4197__B2 (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4198__A1 (.I(net654));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4198__B2 (.I(net127));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4201__A1 (.I(net1734));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4201__A3 (.I(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4201__A4 (.I(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4202__B2 (.I(net732));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4203__A1 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4203__B2 (.I(net245));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4204__A1 (.I(net360));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4204__B2 (.I(net266));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4205__A1 (.I(net328));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4206__A1 (.I(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4206__A2 (.I(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4206__A3 (.I(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4207__A2 (.I(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4211__A1 (.I(net857));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4211__B2 (.I(net780));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4211__C (.I(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4212__I (.I(net469));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4213__I (.I(net826));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4214__A1 (.I(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4214__A3 (.I(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4215__A1 (.I(net795));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4215__B2 (.I(net810));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4215__C (.I(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4218__B2 (.I(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4219__A1 (.I(net173));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4219__B2 (.I(net866));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4222__A1 (.I(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4223__B2 (.I(net748));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4224__A1 (.I(net1732));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4224__A2 (.I(net1730));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4224__A4 (.I(net1729));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4226__A1 (.I(net639));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4227__B2 (.I(net562));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4228__A1 (.I(net406));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4228__B2 (.I(net577));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4229__A1 (.I(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4230__A1 (.I(net297));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4231__A1 (.I(net313));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4234__A2 (.I(_0522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4234__A4 (.I(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4235__A1 (.I(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4235__A2 (.I(_0520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4236__B1 (.I(net1701));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4236__B2 (.I(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4237__I (.I(net445));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4238__I (.I(_0014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4239__I (.I(net501));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4240__I (.I(_0023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4241__I (.I(_0027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4242__I (.I(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4244__I (.I(_0033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4245__I (.I(_0040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4246__A1 (.I(net516));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4248__I (.I(_0051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4249__A1 (.I(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4250__I (.I(net485));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4251__I (.I(_0060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4252__I (.I(_0062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4257__I (.I(net454));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4258__I (.I(_0077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4259__I (.I(_0079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4260__I (.I(_0084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4263__B2 (.I(net423));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4264__I (.I(_0092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4265__I (.I(_0099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4267__I (.I(_0105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4268__I (.I(_0111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4269__I (.I(net376));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4271__C (.I(net1826));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4274__I (.I(net159));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4276__I (.I(_0127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4278__I (.I(net143));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4280__A1 (.I(net252));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4280__B2 (.I(net237));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4280__C (.I(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4281__A1 (.I(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4281__A2 (.I(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4281__A3 (.I(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4281__A4 (.I(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4282__I (.I(_0138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4283__I (.I(_0142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4284__A1 (.I(net411));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4285__I (.I(_0148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4286__I (.I(_0153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4287__A1 (.I(net656));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4287__B2 (.I(net128));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4288__I (.I(_0157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4289__I (.I(_0162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4291__I (.I(_0166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4292__I (.I(_0169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4294__A1 (.I(net1728));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4294__A3 (.I(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4294__A4 (.I(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4295__I (.I(_0175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4296__I (.I(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4297__B2 (.I(net734));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4298__I (.I(_0182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4299__I (.I(_0185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4300__A1 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4300__B2 (.I(net256));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4301__I (.I(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4302__I (.I(_0196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4303__A1 (.I(net361));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4303__B2 (.I(net268));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4304__I (.I(_0201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4305__A1 (.I(net329));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4305__A2 (.I(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4306__A1 (.I(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4306__A2 (.I(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4307__A2 (.I(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4307__A3 (.I(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4308__I (.I(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4309__I (.I(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4311__I (.I(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4312__I (.I(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4313__I (.I(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4316__A1 (.I(net858));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4316__B2 (.I(net781));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4317__I (.I(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4318__I (.I(_0232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4320__I (.I(_0235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4321__I (.I(_0240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4323__A1 (.I(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4323__A3 (.I(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4324__B2 (.I(net812));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4324__C (.I(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4325__I (.I(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4326__I (.I(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4328__I (.I(_0253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4329__I (.I(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4331__B2 (.I(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4332__A1 (.I(net174));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4332__B2 (.I(net877));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4332__C (.I(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4336__I (.I(_0269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4337__I (.I(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4338__I (.I(net567));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4339__A1 (.I(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4340__A1 (.I(net722));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4340__B2 (.I(net749));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4341__A1 (.I(net1726));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4341__A2 (.I(net1724));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4341__A4 (.I(net1723));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4342__I (.I(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4343__I (.I(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4344__A1 (.I(net609));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4345__I (.I(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4346__I (.I(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4347__A1 (.I(net640));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4347__B2 (.I(net531));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4348__I (.I(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4349__I (.I(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4350__A1 (.I(net547));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4351__I (.I(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4352__I (.I(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4353__A1 (.I(net407));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4353__B2 (.I(net579));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4354__A1 (.I(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4354__A2 (.I(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4355__I (.I(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4356__I (.I(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4357__A1 (.I(net298));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4358__I (.I(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4359__I (.I(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4360__A1 (.I(net314));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4360__B2 (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4361__I (.I(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4362__I (.I(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4363__A1 (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4363__B2 (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4366__A2 (.I(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4367__A4 (.I(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4368__A1 (.I(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4368__A2 (.I(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4369__B1 (.I(net1700));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4369__B2 (.I(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4370__I (.I(net556));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4371__I (.I(net502));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4373__A1 (.I(net517));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4374__I (.I(net595));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4376__I (.I(net486));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4378__A3 (.I(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4379__I (.I(net455));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4382__B2 (.I(net424));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4384__I (.I(net377));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4385__A1 (.I(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4386__C (.I(net1825));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4387__I (.I(net160));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4388__I (.I(net144));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4390__A1 (.I(net253));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4390__B2 (.I(net238));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4390__C (.I(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4391__A1 (.I(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4391__A2 (.I(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4391__A3 (.I(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4391__A4 (.I(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4392__A1 (.I(net422));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4393__A1 (.I(net657));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4393__B2 (.I(net129));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4396__A1 (.I(net1722));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4396__A3 (.I(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4396__A4 (.I(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4397__B2 (.I(net735));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4398__A1 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4398__B2 (.I(net267));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4399__A1 (.I(net362));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4399__B2 (.I(net269));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4400__A1 (.I(net330));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4400__A2 (.I(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4401__A1 (.I(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4401__A2 (.I(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4402__A2 (.I(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4402__A3 (.I(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4403__I (.I(net843));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4404__A1 (.I(net874));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4406__A1 (.I(net859));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4406__B2 (.I(net782));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4409__A1 (.I(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4409__A3 (.I(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4410__A1 (.I(net797));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4410__B2 (.I(net813));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4410__C (.I(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4413__B2 (.I(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4414__A1 (.I(net175));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4414__B2 (.I(net884));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4414__C (.I(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4416__I (.I(net578));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4417__A1 (.I(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4418__A1 (.I(net733));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4418__B2 (.I(net750));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4419__A1 (.I(net1720));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4419__A2 (.I(net1718));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4419__A4 (.I(net1717));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4420__A1 (.I(net610));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4421__A1 (.I(net641));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4421__B2 (.I(net532));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4422__A1 (.I(net548));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4423__A1 (.I(net408));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4423__B2 (.I(net580));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4424__A1 (.I(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4424__A2 (.I(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4425__A1 (.I(net299));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4426__A1 (.I(net315));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4426__B2 (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4427__A1 (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4427__B2 (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4428__A2 (.I(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4429__A4 (.I(_0717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4430__A1 (.I(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4430__A2 (.I(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4431__B1 (.I(net1699));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4431__B2 (.I(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4432__I (.I(net667));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4433__I (.I(net503));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4435__A1 (.I(net518));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4436__I (.I(net596));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4439__I (.I(net487));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4442__I (.I(net457));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4445__B2 (.I(net425));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4448__I (.I(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4449__I (.I(net379));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4450__A1 (.I(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4450__A2 (.I(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4451__C (.I(net1824));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4452__I (.I(net161));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4453__I (.I(net146));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4455__A1 (.I(net254));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4455__B2 (.I(net239));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4455__C (.I(_0742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4456__A1 (.I(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4456__A2 (.I(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4456__A3 (.I(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4456__A4 (.I(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4457__A1 (.I(net433));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4458__A1 (.I(net658));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4458__B2 (.I(net130));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4461__A1 (.I(net1716));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4461__A4 (.I(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4462__B2 (.I(net736));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4463__A1 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4463__B2 (.I(net278));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4464__A1 (.I(net363));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4464__B2 (.I(net270));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4465__I (.I(_0012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4466__A1 (.I(net331));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4466__A2 (.I(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4467__A1 (.I(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4467__A2 (.I(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4468__A2 (.I(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4469__I (.I(net845));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4470__A1 (.I(net875));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4472__A1 (.I(net860));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4472__B2 (.I(net783));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4474__I (.I(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4476__A1 (.I(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4476__A3 (.I(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4477__A1 (.I(net798));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4477__B2 (.I(net814));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4477__C (.I(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4480__B2 (.I(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4481__A1 (.I(net176));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4481__B2 (.I(net886));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4481__C (.I(_0768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4483__I (.I(net589));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4484__A1 (.I(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4485__A1 (.I(net744));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4485__B2 (.I(net751));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4486__A1 (.I(net1714));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4486__A2 (.I(net1712));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4486__A4 (.I(net1711));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4487__A1 (.I(net612));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4488__A1 (.I(net642));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4488__B2 (.I(net534));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4489__A1 (.I(net549));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4490__A1 (.I(net409));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4490__B2 (.I(net581));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4491__A1 (.I(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4491__A2 (.I(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4492__A1 (.I(net301));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4493__A1 (.I(net316));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4493__B2 (.I(net68));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4494__A1 (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4494__B2 (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4495__A2 (.I(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4496__A4 (.I(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4497__A1 (.I(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4497__A2 (.I(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4498__B1 (.I(net1698));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4498__B2 (.I(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4500__I (.I(net504));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4502__A1 (.I(net519));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4503__I (.I(net597));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4505__I (.I(net488));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4508__I (.I(net458));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4511__A1 (.I(net395));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4511__B2 (.I(net426));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4513__I (.I(net380));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4514__A1 (.I(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4514__A2 (.I(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4515__C (.I(net1823));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4516__I (.I(net162));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4517__I (.I(net147));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4519__A1 (.I(net255));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4519__B2 (.I(net240));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4519__C (.I(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4520__A1 (.I(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4520__A2 (.I(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4520__A3 (.I(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4520__A4 (.I(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4521__A1 (.I(net444));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4522__A1 (.I(net659));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4522__B2 (.I(net131));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4525__A1 (.I(net1710));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4525__A4 (.I(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4526__B2 (.I(net737));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4527__A1 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4527__B2 (.I(net289));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4528__A1 (.I(net364));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4528__B2 (.I(net271));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4529__A1 (.I(net332));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4529__A2 (.I(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4530__A1 (.I(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4530__A2 (.I(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4531__A2 (.I(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4531__A3 (.I(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4532__I (.I(net846));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4533__A1 (.I(net876));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4535__A1 (.I(net861));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4535__B2 (.I(net784));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4538__A1 (.I(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4538__A3 (.I(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4539__A1 (.I(net799));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4539__B2 (.I(net815));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4539__C (.I(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4542__B2 (.I(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4543__A1 (.I(net177));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4543__B2 (.I(net887));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4543__C (.I(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4545__I (.I(net600));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4546__A1 (.I(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4547__A1 (.I(net755));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4547__B2 (.I(net752));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4548__A1 (.I(net1708));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4548__A2 (.I(net1706));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4548__A4 (.I(net1705));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4550__A1 (.I(net643));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4550__B2 (.I(net535));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4551__A1 (.I(net550));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4552__A1 (.I(net410));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4552__B2 (.I(net582));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4553__A1 (.I(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4553__A2 (.I(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4554__A1 (.I(net302));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4555__A1 (.I(net317));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4555__B2 (.I(net69));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4556__A1 (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4556__B2 (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4557__A2 (.I(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4558__A4 (.I(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4559__A1 (.I(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4559__A2 (.I(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4560__B1 (.I(net1697));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4560__B2 (.I(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4562__I (.I(_0013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4563__I (.I(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4565__I (.I(_0022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4566__I (.I(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4567__I (.I(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4568__A1 (.I(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4569__I (.I(_0032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4570__I (.I(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4571__I (.I(_0039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4572__I (.I(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4573__A1 (.I(net520));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4575__I (.I(_0050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4576__I (.I(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4579__I (.I(_0119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4580__I (.I(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4581__I (.I(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4582__I (.I(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4584__A2 (.I(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4584__A3 (.I(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4584__A4 (.I(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4586__I (.I(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4588__I (.I(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4589__I (.I(net459));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4590__I (.I(_0076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4591__I (.I(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4592__I (.I(_0079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4593__I (.I(_0083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4594__I (.I(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4603__I (.I(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4604__I (.I(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4605__I (.I(_0110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4606__I (.I(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4608__A1 (.I(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4608__A2 (.I(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4608__A3 (.I(_0890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4609__A2 (.I(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4609__B1 (.I(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4609__C (.I(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4611__I (.I(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4613__I (.I(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4615__I (.I(_0124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4616__I (.I(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4617__I (.I(_0127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4618__I (.I(_0129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4619__I (.I(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4621__A2 (.I(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4621__B1 (.I(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4622__A1 (.I(net257));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4622__A2 (.I(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4622__B1 (.I(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4622__C (.I(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4623__A1 (.I(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4623__A2 (.I(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4623__A3 (.I(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4623__A4 (.I(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4625__I (.I(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4627__I (.I(_0912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4628__A1 (.I(net456));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4628__A2 (.I(_0911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4628__B1 (.I(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4628__B2 (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4629__I (.I(_0147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4630__I (.I(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4631__I (.I(_0152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4632__I (.I(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4633__A1 (.I(net660));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4633__B2 (.I(net132));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4643__A2 (.I(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4643__B1 (.I(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4644__A1 (.I(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4644__A3 (.I(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4644__A4 (.I(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4646__I (.I(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4647__I (.I(_0177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4648__I (.I(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4649__A2 (.I(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4649__B2 (.I(net738));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4651__I (.I(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4653__I (.I(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4654__A1 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4654__B2 (.I(net300));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4655__I (.I(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4656__I (.I(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4657__I (.I(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4658__I (.I(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4659__A1 (.I(net365));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4659__B1 (.I(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4659__B2 (.I(net272));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4661__I (.I(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4662__A1 (.I(net335));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4663__A1 (.I(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4663__A2 (.I(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4663__A4 (.I(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4666__I (.I(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4667__I (.I(_0212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4668__I (.I(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4670__CLK (.I(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4671__CLK (.I(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4672__CLK (.I(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4672__D (.I(_2327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4673__CLK (.I(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4673__D (.I(_2328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4674__CLK (.I(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4674__D (.I(_2329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4675__CLK (.I(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4675__D (.I(_2330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4676__CLK (.I(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4677__CLK (.I(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4678__CLK (.I(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4679__CLK (.I(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4680__CLK (.I(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4681__CLK (.I(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4682__CLK (.I(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4682__D (.I(_2309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4683__CLK (.I(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4683__D (.I(_2314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4684__CLK (.I(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4684__D (.I(_2315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4685__CLK (.I(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4685__D (.I(_2316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4686__CLK (.I(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4686__D (.I(_2317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4687__CLK (.I(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4687__D (.I(_2318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4688__CLK (.I(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4688__D (.I(_2319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4689__CLK (.I(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4689__D (.I(_2320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4690__CLK (.I(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4690__D (.I(_2321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4691__CLK (.I(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4691__D (.I(_2322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4692__CLK (.I(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4692__D (.I(_2310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4693__CLK (.I(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4693__D (.I(_2311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4694__CLK (.I(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4694__D (.I(_2312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4695__CLK (.I(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4695__D (.I(_2313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_0_clk_I (.I(clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_1_0__f_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_1_1__f_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1000_I (.I(itasel[193]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1001_I (.I(itasel[194]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1002_I (.I(itasel[195]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1003_I (.I(itasel[196]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1004_I (.I(itasel[197]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1005_I (.I(itasel[198]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1006_I (.I(itasel[199]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1007_I (.I(itasel[19]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1008_I (.I(itasel[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1009_I (.I(itasel[200]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input100_I (.I(itasegm[18]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1010_I (.I(itasel[201]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1011_I (.I(itasel[202]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1012_I (.I(itasel[203]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1013_I (.I(itasel[204]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1014_I (.I(itasel[205]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1015_I (.I(itasel[206]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1016_I (.I(itasel[207]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1017_I (.I(itasel[208]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1018_I (.I(itasel[209]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1019_I (.I(itasel[20]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input101_I (.I(itasegm[190]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1020_I (.I(itasel[210]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1021_I (.I(itasel[211]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1022_I (.I(itasel[212]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1023_I (.I(itasel[213]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1024_I (.I(itasel[214]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1025_I (.I(itasel[215]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1026_I (.I(itasel[216]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1027_I (.I(itasel[217]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1028_I (.I(itasel[218]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1029_I (.I(itasel[219]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input102_I (.I(itasegm[191]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1030_I (.I(itasel[21]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1031_I (.I(itasel[220]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1032_I (.I(itasel[221]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1033_I (.I(itasel[222]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1034_I (.I(itasel[223]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1035_I (.I(itasel[224]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1036_I (.I(itasel[225]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1037_I (.I(itasel[226]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1038_I (.I(itasel[227]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1039_I (.I(itasel[228]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input103_I (.I(itasegm[192]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1040_I (.I(itasel[229]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1041_I (.I(itasel[22]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1042_I (.I(itasel[230]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1043_I (.I(itasel[231]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1044_I (.I(itasel[232]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1045_I (.I(itasel[233]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1046_I (.I(itasel[234]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1047_I (.I(itasel[235]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1048_I (.I(itasel[236]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1049_I (.I(itasel[237]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input104_I (.I(itasegm[193]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1050_I (.I(itasel[238]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1051_I (.I(itasel[239]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1052_I (.I(itasel[23]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1053_I (.I(itasel[240]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1054_I (.I(itasel[241]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1055_I (.I(itasel[242]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1056_I (.I(itasel[243]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1057_I (.I(itasel[244]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1058_I (.I(itasel[245]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1059_I (.I(itasel[246]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input105_I (.I(itasegm[194]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1060_I (.I(itasel[247]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1061_I (.I(itasel[248]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1062_I (.I(itasel[249]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1063_I (.I(itasel[24]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1064_I (.I(itasel[250]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1065_I (.I(itasel[251]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1066_I (.I(itasel[252]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1067_I (.I(itasel[253]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1068_I (.I(itasel[254]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1069_I (.I(itasel[255]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input106_I (.I(itasegm[195]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1070_I (.I(itasel[256]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1071_I (.I(itasel[257]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1072_I (.I(itasel[258]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1073_I (.I(itasel[259]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1074_I (.I(itasel[25]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1075_I (.I(itasel[260]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1076_I (.I(itasel[261]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1077_I (.I(itasel[262]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1078_I (.I(itasel[263]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1079_I (.I(itasel[264]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input107_I (.I(itasegm[196]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1080_I (.I(itasel[265]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1081_I (.I(itasel[266]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1082_I (.I(itasel[267]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1083_I (.I(itasel[268]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1084_I (.I(itasel[269]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1085_I (.I(itasel[26]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1086_I (.I(itasel[270]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1087_I (.I(itasel[271]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1088_I (.I(itasel[272]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1089_I (.I(itasel[273]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input108_I (.I(itasegm[197]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1090_I (.I(itasel[274]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1091_I (.I(itasel[275]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1092_I (.I(itasel[276]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1093_I (.I(itasel[277]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1094_I (.I(itasel[278]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1095_I (.I(itasel[279]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1096_I (.I(itasel[27]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1097_I (.I(itasel[280]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1098_I (.I(itasel[281]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1099_I (.I(itasel[282]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input109_I (.I(itasegm[198]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input10_I (.I(itasegm[108]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1100_I (.I(itasel[283]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1101_I (.I(itasel[284]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1102_I (.I(itasel[285]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1103_I (.I(itasel[286]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1104_I (.I(itasel[287]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1105_I (.I(itasel[288]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1106_I (.I(itasel[289]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1107_I (.I(itasel[28]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1108_I (.I(itasel[290]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1109_I (.I(itasel[291]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input110_I (.I(itasegm[199]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1110_I (.I(itasel[292]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1111_I (.I(itasel[293]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1112_I (.I(itasel[294]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1113_I (.I(itasel[295]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1114_I (.I(itasel[296]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1115_I (.I(itasel[297]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1116_I (.I(itasel[298]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1117_I (.I(itasel[299]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1118_I (.I(itasel[29]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1119_I (.I(itasel[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input111_I (.I(itasegm[19]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1120_I (.I(itasel[300]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1121_I (.I(itasel[301]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1122_I (.I(itasel[302]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1123_I (.I(itasel[303]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1124_I (.I(itasel[304]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1125_I (.I(itasel[305]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1126_I (.I(itasel[306]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1127_I (.I(itasel[307]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1128_I (.I(itasel[308]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1129_I (.I(itasel[309]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input112_I (.I(itasegm[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1130_I (.I(itasel[30]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1131_I (.I(itasel[310]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1132_I (.I(itasel[311]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1133_I (.I(itasel[312]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1134_I (.I(itasel[313]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1135_I (.I(itasel[314]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1136_I (.I(itasel[315]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1137_I (.I(itasel[316]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1138_I (.I(itasel[317]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1139_I (.I(itasel[318]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input113_I (.I(itasegm[200]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1140_I (.I(itasel[319]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1141_I (.I(itasel[31]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1142_I (.I(itasel[320]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1143_I (.I(itasel[321]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1144_I (.I(itasel[322]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1145_I (.I(itasel[323]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1146_I (.I(itasel[324]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1147_I (.I(itasel[325]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1148_I (.I(itasel[326]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1149_I (.I(itasel[327]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input114_I (.I(itasegm[201]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1150_I (.I(itasel[328]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1151_I (.I(itasel[329]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1152_I (.I(itasel[32]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1153_I (.I(itasel[330]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1154_I (.I(itasel[331]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1155_I (.I(itasel[332]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1156_I (.I(itasel[333]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1157_I (.I(itasel[334]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1158_I (.I(itasel[335]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1159_I (.I(itasel[336]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input115_I (.I(itasegm[202]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1160_I (.I(itasel[337]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1161_I (.I(itasel[338]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1162_I (.I(itasel[339]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1163_I (.I(itasel[33]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1164_I (.I(itasel[340]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1165_I (.I(itasel[341]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1166_I (.I(itasel[342]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1167_I (.I(itasel[343]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1168_I (.I(itasel[344]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1169_I (.I(itasel[345]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input116_I (.I(itasegm[203]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1170_I (.I(itasel[346]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1171_I (.I(itasel[347]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1172_I (.I(itasel[348]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1173_I (.I(itasel[349]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1174_I (.I(itasel[34]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1175_I (.I(itasel[350]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1176_I (.I(itasel[351]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1177_I (.I(itasel[352]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1178_I (.I(itasel[353]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1179_I (.I(itasel[354]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input117_I (.I(itasegm[204]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1180_I (.I(itasel[355]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1181_I (.I(itasel[356]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1182_I (.I(itasel[357]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1183_I (.I(itasel[358]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1184_I (.I(itasel[359]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1185_I (.I(itasel[35]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1186_I (.I(itasel[360]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1187_I (.I(itasel[361]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1188_I (.I(itasel[362]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1189_I (.I(itasel[363]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input118_I (.I(itasegm[205]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1190_I (.I(itasel[364]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1191_I (.I(itasel[365]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1192_I (.I(itasel[366]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1193_I (.I(itasel[367]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1194_I (.I(itasel[368]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1195_I (.I(itasel[369]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1196_I (.I(itasel[36]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1197_I (.I(itasel[370]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1198_I (.I(itasel[371]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1199_I (.I(itasel[372]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input119_I (.I(itasegm[206]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input11_I (.I(itasegm[109]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1200_I (.I(itasel[373]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1201_I (.I(itasel[374]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1202_I (.I(itasel[375]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1203_I (.I(itasel[376]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1204_I (.I(itasel[377]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1205_I (.I(itasel[378]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1206_I (.I(itasel[379]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1207_I (.I(itasel[37]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1208_I (.I(itasel[380]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1209_I (.I(itasel[381]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input120_I (.I(itasegm[207]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1210_I (.I(itasel[382]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1211_I (.I(itasel[383]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1212_I (.I(itasel[384]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1213_I (.I(itasel[385]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1214_I (.I(itasel[386]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1215_I (.I(itasel[387]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1216_I (.I(itasel[388]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1217_I (.I(itasel[389]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1218_I (.I(itasel[38]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1219_I (.I(itasel[390]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input121_I (.I(itasegm[208]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1220_I (.I(itasel[391]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1221_I (.I(itasel[392]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1222_I (.I(itasel[393]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1223_I (.I(itasel[394]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1224_I (.I(itasel[395]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1225_I (.I(itasel[396]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1226_I (.I(itasel[397]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1227_I (.I(itasel[398]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1228_I (.I(itasel[399]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1229_I (.I(itasel[39]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input122_I (.I(itasegm[209]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1230_I (.I(itasel[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1231_I (.I(itasel[400]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1232_I (.I(itasel[401]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1233_I (.I(itasel[402]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1234_I (.I(itasel[403]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1235_I (.I(itasel[404]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1236_I (.I(itasel[405]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1237_I (.I(itasel[406]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1238_I (.I(itasel[407]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1239_I (.I(itasel[408]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input123_I (.I(itasegm[20]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1240_I (.I(itasel[409]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1241_I (.I(itasel[40]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1242_I (.I(itasel[410]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1243_I (.I(itasel[411]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1244_I (.I(itasel[412]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1245_I (.I(itasel[413]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1246_I (.I(itasel[414]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1247_I (.I(itasel[415]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1248_I (.I(itasel[416]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1249_I (.I(itasel[417]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input124_I (.I(itasegm[210]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1250_I (.I(itasel[418]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1251_I (.I(itasel[419]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1252_I (.I(itasel[41]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1253_I (.I(itasel[420]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1254_I (.I(itasel[421]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1255_I (.I(itasel[422]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1256_I (.I(itasel[423]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1257_I (.I(itasel[424]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1258_I (.I(itasel[425]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1259_I (.I(itasel[426]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input125_I (.I(itasegm[211]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1260_I (.I(itasel[427]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1261_I (.I(itasel[428]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1262_I (.I(itasel[429]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1263_I (.I(itasel[42]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1264_I (.I(itasel[430]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1265_I (.I(itasel[431]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1266_I (.I(itasel[432]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1267_I (.I(itasel[433]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1268_I (.I(itasel[434]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1269_I (.I(itasel[435]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input126_I (.I(itasegm[212]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1270_I (.I(itasel[436]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1271_I (.I(itasel[437]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1272_I (.I(itasel[438]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1273_I (.I(itasel[439]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1274_I (.I(itasel[43]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1275_I (.I(itasel[440]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1276_I (.I(itasel[441]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1277_I (.I(itasel[442]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1278_I (.I(itasel[443]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1279_I (.I(itasel[444]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input127_I (.I(itasegm[213]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1280_I (.I(itasel[445]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1281_I (.I(itasel[446]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1282_I (.I(itasel[447]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1283_I (.I(itasel[448]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1284_I (.I(itasel[449]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1285_I (.I(itasel[44]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1286_I (.I(itasel[450]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1287_I (.I(itasel[451]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1288_I (.I(itasel[452]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1289_I (.I(itasel[453]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input128_I (.I(itasegm[214]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1290_I (.I(itasel[454]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1291_I (.I(itasel[455]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1292_I (.I(itasel[456]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1293_I (.I(itasel[457]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1294_I (.I(itasel[458]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1295_I (.I(itasel[459]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1296_I (.I(itasel[45]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1297_I (.I(itasel[460]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1298_I (.I(itasel[461]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1299_I (.I(itasel[462]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input129_I (.I(itasegm[215]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input12_I (.I(itasegm[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1300_I (.I(itasel[463]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1301_I (.I(itasel[464]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1302_I (.I(itasel[465]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1303_I (.I(itasel[466]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1304_I (.I(itasel[467]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1305_I (.I(itasel[468]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1306_I (.I(itasel[469]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1307_I (.I(itasel[46]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1308_I (.I(itasel[470]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1309_I (.I(itasel[471]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input130_I (.I(itasegm[216]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1310_I (.I(itasel[472]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1311_I (.I(itasel[473]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1312_I (.I(itasel[474]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1313_I (.I(itasel[475]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1314_I (.I(itasel[476]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1315_I (.I(itasel[477]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1316_I (.I(itasel[478]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1317_I (.I(itasel[479]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1318_I (.I(itasel[47]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1319_I (.I(itasel[480]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input131_I (.I(itasegm[217]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1320_I (.I(itasel[481]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1321_I (.I(itasel[482]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1322_I (.I(itasel[483]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1323_I (.I(itasel[484]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1324_I (.I(itasel[485]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1325_I (.I(itasel[486]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1326_I (.I(itasel[487]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1327_I (.I(itasel[488]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1328_I (.I(itasel[489]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1329_I (.I(itasel[48]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input132_I (.I(itasegm[218]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1330_I (.I(itasel[490]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1331_I (.I(itasel[491]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1332_I (.I(itasel[492]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1333_I (.I(itasel[493]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1334_I (.I(itasel[494]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1335_I (.I(itasel[495]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1336_I (.I(itasel[496]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1337_I (.I(itasel[497]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1338_I (.I(itasel[498]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1339_I (.I(itasel[499]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input133_I (.I(itasegm[219]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1340_I (.I(itasel[49]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1341_I (.I(itasel[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1342_I (.I(itasel[500]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1343_I (.I(itasel[501]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1344_I (.I(itasel[502]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1345_I (.I(itasel[503]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1346_I (.I(itasel[504]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1347_I (.I(itasel[505]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1348_I (.I(itasel[506]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1349_I (.I(itasel[507]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input134_I (.I(itasegm[21]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1350_I (.I(itasel[508]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1351_I (.I(itasel[509]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1352_I (.I(itasel[50]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1353_I (.I(itasel[510]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1354_I (.I(itasel[511]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1355_I (.I(itasel[512]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1356_I (.I(itasel[513]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1357_I (.I(itasel[514]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1358_I (.I(itasel[515]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1359_I (.I(itasel[516]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input135_I (.I(itasegm[220]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1360_I (.I(itasel[517]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1361_I (.I(itasel[518]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1362_I (.I(itasel[519]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1363_I (.I(itasel[51]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1364_I (.I(itasel[520]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1365_I (.I(itasel[521]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1366_I (.I(itasel[522]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1367_I (.I(itasel[523]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1368_I (.I(itasel[524]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1369_I (.I(itasel[525]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input136_I (.I(itasegm[221]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1370_I (.I(itasel[526]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1371_I (.I(itasel[527]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1372_I (.I(itasel[528]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1373_I (.I(itasel[529]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1374_I (.I(itasel[52]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1375_I (.I(itasel[530]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1376_I (.I(itasel[531]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1377_I (.I(itasel[532]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1378_I (.I(itasel[533]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1379_I (.I(itasel[534]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input137_I (.I(itasegm[222]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1380_I (.I(itasel[535]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1381_I (.I(itasel[536]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1382_I (.I(itasel[537]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1383_I (.I(itasel[538]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1384_I (.I(itasel[539]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1385_I (.I(itasel[53]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1386_I (.I(itasel[540]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1387_I (.I(itasel[541]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1388_I (.I(itasel[542]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1389_I (.I(itasel[543]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input138_I (.I(itasegm[223]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1390_I (.I(itasel[544]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1391_I (.I(itasel[545]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1392_I (.I(itasel[546]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1393_I (.I(itasel[547]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1394_I (.I(itasel[548]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1395_I (.I(itasel[549]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1396_I (.I(itasel[54]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1397_I (.I(itasel[550]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1398_I (.I(itasel[551]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1399_I (.I(itasel[552]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input139_I (.I(itasegm[224]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input13_I (.I(itasegm[110]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1400_I (.I(itasel[553]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1401_I (.I(itasel[554]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1402_I (.I(itasel[555]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1403_I (.I(itasel[556]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1404_I (.I(itasel[557]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1405_I (.I(itasel[558]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1406_I (.I(itasel[559]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1407_I (.I(itasel[55]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1408_I (.I(itasel[560]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1409_I (.I(itasel[561]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input140_I (.I(itasegm[225]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1410_I (.I(itasel[562]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1411_I (.I(itasel[563]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1412_I (.I(itasel[564]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1413_I (.I(itasel[565]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1414_I (.I(itasel[566]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1415_I (.I(itasel[567]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1416_I (.I(itasel[568]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1417_I (.I(itasel[569]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1418_I (.I(itasel[56]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1419_I (.I(itasel[570]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input141_I (.I(itasegm[226]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1420_I (.I(itasel[571]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1421_I (.I(itasel[572]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1422_I (.I(itasel[573]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1423_I (.I(itasel[574]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1424_I (.I(itasel[575]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1425_I (.I(itasel[576]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1426_I (.I(itasel[577]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1427_I (.I(itasel[578]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1428_I (.I(itasel[579]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1429_I (.I(itasel[57]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input142_I (.I(itasegm[227]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1430_I (.I(itasel[580]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1431_I (.I(itasel[581]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1432_I (.I(itasel[582]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1433_I (.I(itasel[583]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1434_I (.I(itasel[584]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1435_I (.I(itasel[585]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1436_I (.I(itasel[586]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1437_I (.I(itasel[587]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1438_I (.I(itasel[588]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1439_I (.I(itasel[589]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input143_I (.I(itasegm[228]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1440_I (.I(itasel[58]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1441_I (.I(itasel[590]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1442_I (.I(itasel[591]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1443_I (.I(itasel[592]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1444_I (.I(itasel[593]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1445_I (.I(itasel[594]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1446_I (.I(itasel[595]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1447_I (.I(itasel[596]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1448_I (.I(itasel[597]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1449_I (.I(itasel[598]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input144_I (.I(itasegm[229]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1450_I (.I(itasel[599]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1451_I (.I(itasel[59]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1452_I (.I(itasel[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1453_I (.I(itasel[600]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1454_I (.I(itasel[601]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1455_I (.I(itasel[602]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1456_I (.I(itasel[603]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1457_I (.I(itasel[604]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1458_I (.I(itasel[605]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1459_I (.I(itasel[606]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input145_I (.I(itasegm[22]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1460_I (.I(itasel[607]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1461_I (.I(itasel[608]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1462_I (.I(itasel[609]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1463_I (.I(itasel[60]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1464_I (.I(itasel[610]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1465_I (.I(itasel[611]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1466_I (.I(itasel[612]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1467_I (.I(itasel[613]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1468_I (.I(itasel[614]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1469_I (.I(itasel[615]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input146_I (.I(itasegm[230]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1470_I (.I(itasel[616]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1471_I (.I(itasel[617]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1472_I (.I(itasel[618]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1473_I (.I(itasel[619]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1474_I (.I(itasel[61]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1475_I (.I(itasel[620]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1476_I (.I(itasel[621]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1477_I (.I(itasel[622]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1478_I (.I(itasel[623]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1479_I (.I(itasel[624]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input147_I (.I(itasegm[231]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1480_I (.I(itasel[625]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1481_I (.I(itasel[626]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1482_I (.I(itasel[627]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1483_I (.I(itasel[628]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1484_I (.I(itasel[629]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1485_I (.I(itasel[62]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1486_I (.I(itasel[630]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1487_I (.I(itasel[631]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1488_I (.I(itasel[632]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1489_I (.I(itasel[633]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input148_I (.I(itasegm[232]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1490_I (.I(itasel[634]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1491_I (.I(itasel[635]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1492_I (.I(itasel[636]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1493_I (.I(itasel[637]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1494_I (.I(itasel[638]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1495_I (.I(itasel[639]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1496_I (.I(itasel[63]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1497_I (.I(itasel[640]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1498_I (.I(itasel[641]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1499_I (.I(itasel[642]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input149_I (.I(itasegm[233]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input14_I (.I(itasegm[111]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1500_I (.I(itasel[643]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1501_I (.I(itasel[644]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1502_I (.I(itasel[645]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1503_I (.I(itasel[646]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1504_I (.I(itasel[647]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1505_I (.I(itasel[648]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1506_I (.I(itasel[649]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1507_I (.I(itasel[64]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1508_I (.I(itasel[650]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1509_I (.I(itasel[651]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input150_I (.I(itasegm[234]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1510_I (.I(itasel[652]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1511_I (.I(itasel[653]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1512_I (.I(itasel[654]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1513_I (.I(itasel[655]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1514_I (.I(itasel[656]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1515_I (.I(itasel[657]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1516_I (.I(itasel[658]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1517_I (.I(itasel[659]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1518_I (.I(itasel[65]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1519_I (.I(itasel[660]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input151_I (.I(itasegm[235]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1520_I (.I(itasel[661]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1521_I (.I(itasel[662]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1522_I (.I(itasel[663]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1523_I (.I(itasel[664]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1524_I (.I(itasel[665]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1525_I (.I(itasel[666]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1526_I (.I(itasel[667]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1527_I (.I(itasel[668]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1528_I (.I(itasel[669]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1529_I (.I(itasel[66]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input152_I (.I(itasegm[236]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1530_I (.I(itasel[670]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1531_I (.I(itasel[671]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1532_I (.I(itasel[672]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1533_I (.I(itasel[673]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1534_I (.I(itasel[674]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1535_I (.I(itasel[675]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1536_I (.I(itasel[676]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1537_I (.I(itasel[677]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1538_I (.I(itasel[678]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1539_I (.I(itasel[679]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input153_I (.I(itasegm[237]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1540_I (.I(itasel[67]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1541_I (.I(itasel[680]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1542_I (.I(itasel[681]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1543_I (.I(itasel[682]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1544_I (.I(itasel[683]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1545_I (.I(itasel[684]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1546_I (.I(itasel[685]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1547_I (.I(itasel[686]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1548_I (.I(itasel[687]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1549_I (.I(itasel[688]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input154_I (.I(itasegm[238]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1550_I (.I(itasel[689]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1551_I (.I(itasel[68]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1552_I (.I(itasel[690]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1553_I (.I(itasel[691]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1554_I (.I(itasel[692]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1555_I (.I(itasel[693]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1556_I (.I(itasel[694]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1557_I (.I(itasel[695]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1558_I (.I(itasel[696]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1559_I (.I(itasel[697]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input155_I (.I(itasegm[239]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1560_I (.I(itasel[698]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1561_I (.I(itasel[699]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1562_I (.I(itasel[69]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1563_I (.I(itasel[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1564_I (.I(itasel[700]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1565_I (.I(itasel[701]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1566_I (.I(itasel[702]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1567_I (.I(itasel[703]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1568_I (.I(itasel[704]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1569_I (.I(itasel[705]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input156_I (.I(itasegm[23]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1570_I (.I(itasel[706]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1571_I (.I(itasel[707]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1572_I (.I(itasel[708]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1573_I (.I(itasel[709]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1574_I (.I(itasel[70]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1575_I (.I(itasel[710]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1576_I (.I(itasel[711]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1577_I (.I(itasel[712]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1578_I (.I(itasel[713]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1579_I (.I(itasel[714]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input157_I (.I(itasegm[240]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1580_I (.I(itasel[715]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1581_I (.I(itasel[716]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1582_I (.I(itasel[717]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1583_I (.I(itasel[718]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1584_I (.I(itasel[719]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1585_I (.I(itasel[71]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1586_I (.I(itasel[720]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1587_I (.I(itasel[721]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1588_I (.I(itasel[722]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1589_I (.I(itasel[723]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input158_I (.I(itasegm[241]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1590_I (.I(itasel[724]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1591_I (.I(itasel[725]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1592_I (.I(itasel[726]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1593_I (.I(itasel[727]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1594_I (.I(itasel[728]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1595_I (.I(itasel[729]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1596_I (.I(itasel[72]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1597_I (.I(itasel[730]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1598_I (.I(itasel[731]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1599_I (.I(itasel[732]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input159_I (.I(itasegm[242]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input15_I (.I(itasegm[112]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1600_I (.I(itasel[733]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1601_I (.I(itasel[734]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1602_I (.I(itasel[735]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1603_I (.I(itasel[736]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1604_I (.I(itasel[737]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1605_I (.I(itasel[738]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1606_I (.I(itasel[739]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1607_I (.I(itasel[73]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1608_I (.I(itasel[740]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1609_I (.I(itasel[741]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input160_I (.I(itasegm[243]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1610_I (.I(itasel[742]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1611_I (.I(itasel[743]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1612_I (.I(itasel[744]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1613_I (.I(itasel[745]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1614_I (.I(itasel[746]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1615_I (.I(itasel[747]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1616_I (.I(itasel[748]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1617_I (.I(itasel[749]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1618_I (.I(itasel[74]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1619_I (.I(itasel[750]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input161_I (.I(itasegm[244]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1620_I (.I(itasel[751]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1621_I (.I(itasel[752]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1622_I (.I(itasel[753]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1623_I (.I(itasel[754]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1624_I (.I(itasel[755]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1625_I (.I(itasel[756]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1626_I (.I(itasel[757]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1627_I (.I(itasel[758]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1628_I (.I(itasel[759]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1629_I (.I(itasel[75]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input162_I (.I(itasegm[245]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1630_I (.I(itasel[760]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1631_I (.I(itasel[761]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1632_I (.I(itasel[762]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1633_I (.I(itasel[763]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1634_I (.I(itasel[764]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1635_I (.I(itasel[765]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1636_I (.I(itasel[766]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1637_I (.I(itasel[767]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1638_I (.I(itasel[76]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1639_I (.I(itasel[77]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input163_I (.I(itasegm[246]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1640_I (.I(itasel[78]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1641_I (.I(itasel[79]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1642_I (.I(itasel[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1643_I (.I(itasel[80]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1644_I (.I(itasel[81]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1645_I (.I(itasel[82]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1646_I (.I(itasel[83]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1647_I (.I(itasel[84]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1648_I (.I(itasel[85]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1649_I (.I(itasel[86]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input164_I (.I(itasegm[247]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1650_I (.I(itasel[87]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1651_I (.I(itasel[88]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1652_I (.I(itasel[89]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1653_I (.I(itasel[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1654_I (.I(itasel[90]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1655_I (.I(itasel[91]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1656_I (.I(itasel[92]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1657_I (.I(itasel[93]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1658_I (.I(itasel[94]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1659_I (.I(itasel[95]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input165_I (.I(itasegm[248]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1660_I (.I(itasel[96]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1661_I (.I(itasel[97]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1662_I (.I(itasel[98]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1663_I (.I(itasel[99]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1664_I (.I(itasel[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1665_I (.I(nsel[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1666_I (.I(nsel[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1667_I (.I(nsel[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1668_I (.I(nsel[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1669_I (.I(nsel[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input166_I (.I(itasegm[249]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1670_I (.I(nsel[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input167_I (.I(itasegm[24]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input168_I (.I(itasegm[250]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input169_I (.I(itasegm[251]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input16_I (.I(itasegm[113]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input170_I (.I(itasegm[252]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input171_I (.I(itasegm[253]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input172_I (.I(itasegm[254]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input173_I (.I(itasegm[255]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input174_I (.I(itasegm[256]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input175_I (.I(itasegm[257]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input176_I (.I(itasegm[258]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input177_I (.I(itasegm[259]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input178_I (.I(itasegm[25]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input179_I (.I(itasegm[260]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input17_I (.I(itasegm[114]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input180_I (.I(itasegm[261]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input181_I (.I(itasegm[262]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input182_I (.I(itasegm[263]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input183_I (.I(itasegm[264]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input184_I (.I(itasegm[265]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input185_I (.I(itasegm[266]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input186_I (.I(itasegm[267]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input187_I (.I(itasegm[268]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input188_I (.I(itasegm[269]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input189_I (.I(itasegm[26]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input18_I (.I(itasegm[115]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input190_I (.I(itasegm[270]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input191_I (.I(itasegm[271]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input192_I (.I(itasegm[272]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input193_I (.I(itasegm[273]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input194_I (.I(itasegm[274]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input195_I (.I(itasegm[275]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input196_I (.I(itasegm[276]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input197_I (.I(itasegm[277]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input198_I (.I(itasegm[278]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input199_I (.I(itasegm[279]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input19_I (.I(itasegm[116]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(itasegm[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input200_I (.I(itasegm[27]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input201_I (.I(itasegm[280]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input202_I (.I(itasegm[281]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input203_I (.I(itasegm[282]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input204_I (.I(itasegm[283]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input205_I (.I(itasegm[284]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input206_I (.I(itasegm[285]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input207_I (.I(itasegm[286]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input208_I (.I(itasegm[287]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input209_I (.I(itasegm[288]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input20_I (.I(itasegm[117]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input210_I (.I(itasegm[289]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input211_I (.I(itasegm[28]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input212_I (.I(itasegm[290]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input213_I (.I(itasegm[291]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input214_I (.I(itasegm[292]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input215_I (.I(itasegm[293]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input216_I (.I(itasegm[294]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input217_I (.I(itasegm[295]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input218_I (.I(itasegm[296]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input219_I (.I(itasegm[297]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input21_I (.I(itasegm[118]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input220_I (.I(itasegm[298]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input221_I (.I(itasegm[299]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input222_I (.I(itasegm[29]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input223_I (.I(itasegm[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input224_I (.I(itasegm[300]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input225_I (.I(itasegm[301]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input226_I (.I(itasegm[302]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input227_I (.I(itasegm[303]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input228_I (.I(itasegm[304]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input229_I (.I(itasegm[305]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input22_I (.I(itasegm[119]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input230_I (.I(itasegm[306]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input231_I (.I(itasegm[307]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input232_I (.I(itasegm[308]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input233_I (.I(itasegm[309]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input234_I (.I(itasegm[30]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input235_I (.I(itasegm[310]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input236_I (.I(itasegm[311]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input237_I (.I(itasegm[312]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input238_I (.I(itasegm[313]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input239_I (.I(itasegm[314]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input23_I (.I(itasegm[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input240_I (.I(itasegm[315]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input241_I (.I(itasegm[316]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input242_I (.I(itasegm[317]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input243_I (.I(itasegm[318]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input244_I (.I(itasegm[319]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input245_I (.I(itasegm[31]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input246_I (.I(itasegm[320]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input247_I (.I(itasegm[321]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input248_I (.I(itasegm[322]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input249_I (.I(itasegm[323]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input24_I (.I(itasegm[120]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input250_I (.I(itasegm[324]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input251_I (.I(itasegm[325]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input252_I (.I(itasegm[326]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input253_I (.I(itasegm[327]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input254_I (.I(itasegm[328]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input255_I (.I(itasegm[329]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input256_I (.I(itasegm[32]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input257_I (.I(itasegm[330]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input258_I (.I(itasegm[331]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input259_I (.I(itasegm[332]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input25_I (.I(itasegm[121]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input260_I (.I(itasegm[333]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input261_I (.I(itasegm[334]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input262_I (.I(itasegm[335]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input263_I (.I(itasegm[336]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input264_I (.I(itasegm[337]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input265_I (.I(itasegm[338]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input266_I (.I(itasegm[339]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input267_I (.I(itasegm[33]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input268_I (.I(itasegm[340]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input269_I (.I(itasegm[341]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input26_I (.I(itasegm[122]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input270_I (.I(itasegm[342]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input271_I (.I(itasegm[343]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input272_I (.I(itasegm[344]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input273_I (.I(itasegm[345]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input274_I (.I(itasegm[346]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input275_I (.I(itasegm[347]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input276_I (.I(itasegm[348]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input277_I (.I(itasegm[349]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input278_I (.I(itasegm[34]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input279_I (.I(itasegm[350]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input27_I (.I(itasegm[123]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input280_I (.I(itasegm[351]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input281_I (.I(itasegm[352]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input282_I (.I(itasegm[353]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input283_I (.I(itasegm[354]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input284_I (.I(itasegm[355]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input285_I (.I(itasegm[356]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input286_I (.I(itasegm[357]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input287_I (.I(itasegm[358]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input288_I (.I(itasegm[359]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input289_I (.I(itasegm[35]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input28_I (.I(itasegm[124]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input290_I (.I(itasegm[360]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input291_I (.I(itasegm[361]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input292_I (.I(itasegm[362]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input293_I (.I(itasegm[363]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input294_I (.I(itasegm[364]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input295_I (.I(itasegm[365]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input296_I (.I(itasegm[366]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input297_I (.I(itasegm[367]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input298_I (.I(itasegm[368]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input299_I (.I(itasegm[369]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input29_I (.I(itasegm[125]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(itasegm[100]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input300_I (.I(itasegm[36]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input301_I (.I(itasegm[370]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input302_I (.I(itasegm[371]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input303_I (.I(itasegm[372]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input304_I (.I(itasegm[373]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input305_I (.I(itasegm[374]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input306_I (.I(itasegm[375]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input307_I (.I(itasegm[376]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input308_I (.I(itasegm[377]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input309_I (.I(itasegm[378]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input30_I (.I(itasegm[126]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input310_I (.I(itasegm[379]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input311_I (.I(itasegm[37]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input312_I (.I(itasegm[380]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input313_I (.I(itasegm[381]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input314_I (.I(itasegm[382]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input315_I (.I(itasegm[383]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input316_I (.I(itasegm[384]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input317_I (.I(itasegm[385]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input318_I (.I(itasegm[386]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input319_I (.I(itasegm[387]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input31_I (.I(itasegm[127]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input320_I (.I(itasegm[388]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input321_I (.I(itasegm[389]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input322_I (.I(itasegm[38]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input323_I (.I(itasegm[390]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input324_I (.I(itasegm[391]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input325_I (.I(itasegm[392]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input326_I (.I(itasegm[393]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input327_I (.I(itasegm[394]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input328_I (.I(itasegm[395]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input329_I (.I(itasegm[396]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input32_I (.I(itasegm[128]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input330_I (.I(itasegm[397]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input331_I (.I(itasegm[398]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input332_I (.I(itasegm[399]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input333_I (.I(itasegm[39]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input334_I (.I(itasegm[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input335_I (.I(itasegm[400]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input336_I (.I(itasegm[401]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input337_I (.I(itasegm[402]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input338_I (.I(itasegm[403]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input339_I (.I(itasegm[404]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input33_I (.I(itasegm[129]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input340_I (.I(itasegm[405]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input341_I (.I(itasegm[406]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input342_I (.I(itasegm[407]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input343_I (.I(itasegm[408]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input344_I (.I(itasegm[409]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input345_I (.I(itasegm[40]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input346_I (.I(itasegm[410]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input347_I (.I(itasegm[411]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input348_I (.I(itasegm[412]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input349_I (.I(itasegm[413]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input34_I (.I(itasegm[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input350_I (.I(itasegm[414]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input351_I (.I(itasegm[415]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input352_I (.I(itasegm[416]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input353_I (.I(itasegm[417]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input354_I (.I(itasegm[418]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input355_I (.I(itasegm[419]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input356_I (.I(itasegm[41]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input357_I (.I(itasegm[420]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input358_I (.I(itasegm[421]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input359_I (.I(itasegm[422]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input35_I (.I(itasegm[130]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input360_I (.I(itasegm[423]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input361_I (.I(itasegm[424]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input362_I (.I(itasegm[425]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input363_I (.I(itasegm[426]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input364_I (.I(itasegm[427]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input365_I (.I(itasegm[428]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input366_I (.I(itasegm[429]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input367_I (.I(itasegm[42]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input368_I (.I(itasegm[430]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input369_I (.I(itasegm[431]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input36_I (.I(itasegm[131]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input370_I (.I(itasegm[432]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input371_I (.I(itasegm[433]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input372_I (.I(itasegm[434]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input373_I (.I(itasegm[435]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input374_I (.I(itasegm[436]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input375_I (.I(itasegm[437]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input376_I (.I(itasegm[438]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input377_I (.I(itasegm[439]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input378_I (.I(itasegm[43]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input379_I (.I(itasegm[440]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input37_I (.I(itasegm[132]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input380_I (.I(itasegm[441]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input381_I (.I(itasegm[442]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input382_I (.I(itasegm[443]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input383_I (.I(itasegm[444]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input384_I (.I(itasegm[445]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input385_I (.I(itasegm[446]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input386_I (.I(itasegm[447]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input387_I (.I(itasegm[448]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input388_I (.I(itasegm[449]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input389_I (.I(itasegm[44]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input38_I (.I(itasegm[133]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input390_I (.I(itasegm[450]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input391_I (.I(itasegm[451]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input392_I (.I(itasegm[452]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input393_I (.I(itasegm[453]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input394_I (.I(itasegm[454]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input395_I (.I(itasegm[455]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input396_I (.I(itasegm[456]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input397_I (.I(itasegm[457]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input398_I (.I(itasegm[458]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input399_I (.I(itasegm[459]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input39_I (.I(itasegm[134]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(itasegm[101]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input400_I (.I(itasegm[45]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input401_I (.I(itasegm[460]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input402_I (.I(itasegm[461]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input403_I (.I(itasegm[462]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input404_I (.I(itasegm[463]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input405_I (.I(itasegm[464]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input406_I (.I(itasegm[465]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input407_I (.I(itasegm[466]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input408_I (.I(itasegm[467]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input409_I (.I(itasegm[468]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input40_I (.I(itasegm[135]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input410_I (.I(itasegm[469]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input411_I (.I(itasegm[46]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input412_I (.I(itasegm[470]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input413_I (.I(itasegm[471]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input414_I (.I(itasegm[472]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input415_I (.I(itasegm[473]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input416_I (.I(itasegm[474]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input417_I (.I(itasegm[475]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input418_I (.I(itasegm[476]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input419_I (.I(itasegm[477]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input41_I (.I(itasegm[136]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input420_I (.I(itasegm[478]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input421_I (.I(itasegm[479]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input422_I (.I(itasegm[47]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input423_I (.I(itasegm[480]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input424_I (.I(itasegm[481]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input425_I (.I(itasegm[482]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input426_I (.I(itasegm[483]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input427_I (.I(itasegm[484]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input428_I (.I(itasegm[485]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input429_I (.I(itasegm[486]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input42_I (.I(itasegm[137]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input430_I (.I(itasegm[487]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input431_I (.I(itasegm[488]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input432_I (.I(itasegm[489]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input433_I (.I(itasegm[48]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input434_I (.I(itasegm[490]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input435_I (.I(itasegm[491]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input436_I (.I(itasegm[492]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input437_I (.I(itasegm[493]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input438_I (.I(itasegm[494]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input439_I (.I(itasegm[495]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input43_I (.I(itasegm[138]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input440_I (.I(itasegm[496]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input441_I (.I(itasegm[497]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input442_I (.I(itasegm[498]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input443_I (.I(itasegm[499]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input444_I (.I(itasegm[49]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input445_I (.I(itasegm[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input446_I (.I(itasegm[500]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input447_I (.I(itasegm[501]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input448_I (.I(itasegm[502]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input449_I (.I(itasegm[503]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input44_I (.I(itasegm[139]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input450_I (.I(itasegm[504]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input451_I (.I(itasegm[505]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input452_I (.I(itasegm[506]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input453_I (.I(itasegm[507]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input454_I (.I(itasegm[508]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input455_I (.I(itasegm[509]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input456_I (.I(itasegm[50]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input457_I (.I(itasegm[510]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input458_I (.I(itasegm[511]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input459_I (.I(itasegm[512]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input45_I (.I(itasegm[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input460_I (.I(itasegm[513]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input461_I (.I(itasegm[514]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input462_I (.I(itasegm[515]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input463_I (.I(itasegm[516]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input464_I (.I(itasegm[517]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input465_I (.I(itasegm[518]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input466_I (.I(itasegm[519]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input467_I (.I(itasegm[51]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input468_I (.I(itasegm[520]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input469_I (.I(itasegm[521]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input46_I (.I(itasegm[140]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input470_I (.I(itasegm[522]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input471_I (.I(itasegm[523]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input472_I (.I(itasegm[524]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input473_I (.I(itasegm[525]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input474_I (.I(itasegm[526]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input475_I (.I(itasegm[527]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input476_I (.I(itasegm[528]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input477_I (.I(itasegm[529]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input478_I (.I(itasegm[52]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input479_I (.I(itasegm[530]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input47_I (.I(itasegm[141]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input480_I (.I(itasegm[531]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input481_I (.I(itasegm[532]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input482_I (.I(itasegm[533]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input483_I (.I(itasegm[534]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input484_I (.I(itasegm[535]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input485_I (.I(itasegm[536]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input486_I (.I(itasegm[537]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input487_I (.I(itasegm[538]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input488_I (.I(itasegm[539]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input489_I (.I(itasegm[53]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input48_I (.I(itasegm[142]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input490_I (.I(itasegm[540]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input491_I (.I(itasegm[541]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input492_I (.I(itasegm[542]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input493_I (.I(itasegm[543]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input494_I (.I(itasegm[544]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input495_I (.I(itasegm[545]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input496_I (.I(itasegm[546]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input497_I (.I(itasegm[547]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input498_I (.I(itasegm[548]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input499_I (.I(itasegm[549]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input49_I (.I(itasegm[143]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(itasegm[102]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input500_I (.I(itasegm[54]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input501_I (.I(itasegm[550]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input502_I (.I(itasegm[551]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input503_I (.I(itasegm[552]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input504_I (.I(itasegm[553]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input505_I (.I(itasegm[554]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input506_I (.I(itasegm[555]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input507_I (.I(itasegm[556]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input508_I (.I(itasegm[557]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input509_I (.I(itasegm[558]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input50_I (.I(itasegm[144]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input510_I (.I(itasegm[559]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input511_I (.I(itasegm[55]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input512_I (.I(itasegm[560]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input513_I (.I(itasegm[561]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input514_I (.I(itasegm[562]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input515_I (.I(itasegm[563]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input516_I (.I(itasegm[564]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input517_I (.I(itasegm[565]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input518_I (.I(itasegm[566]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input519_I (.I(itasegm[567]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input51_I (.I(itasegm[145]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input520_I (.I(itasegm[568]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input521_I (.I(itasegm[569]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input522_I (.I(itasegm[56]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input523_I (.I(itasegm[570]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input524_I (.I(itasegm[571]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input525_I (.I(itasegm[572]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input526_I (.I(itasegm[573]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input527_I (.I(itasegm[574]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input528_I (.I(itasegm[575]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input529_I (.I(itasegm[576]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input52_I (.I(itasegm[146]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input530_I (.I(itasegm[577]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input531_I (.I(itasegm[578]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input532_I (.I(itasegm[579]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input533_I (.I(itasegm[57]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input534_I (.I(itasegm[580]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input535_I (.I(itasegm[581]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input536_I (.I(itasegm[582]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input537_I (.I(itasegm[583]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input538_I (.I(itasegm[584]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input539_I (.I(itasegm[585]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input53_I (.I(itasegm[147]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input540_I (.I(itasegm[586]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input541_I (.I(itasegm[587]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input542_I (.I(itasegm[588]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input543_I (.I(itasegm[589]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input544_I (.I(itasegm[58]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input545_I (.I(itasegm[590]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input546_I (.I(itasegm[591]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input547_I (.I(itasegm[592]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input548_I (.I(itasegm[593]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input549_I (.I(itasegm[594]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input54_I (.I(itasegm[148]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input550_I (.I(itasegm[595]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input551_I (.I(itasegm[596]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input552_I (.I(itasegm[597]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input553_I (.I(itasegm[598]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input554_I (.I(itasegm[599]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input555_I (.I(itasegm[59]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input556_I (.I(itasegm[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input557_I (.I(itasegm[600]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input558_I (.I(itasegm[601]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input559_I (.I(itasegm[602]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input55_I (.I(itasegm[149]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input560_I (.I(itasegm[603]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input561_I (.I(itasegm[604]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input562_I (.I(itasegm[605]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input563_I (.I(itasegm[606]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input564_I (.I(itasegm[607]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input565_I (.I(itasegm[608]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input566_I (.I(itasegm[609]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input567_I (.I(itasegm[60]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input568_I (.I(itasegm[610]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input569_I (.I(itasegm[611]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input56_I (.I(itasegm[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input570_I (.I(itasegm[612]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input571_I (.I(itasegm[613]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input572_I (.I(itasegm[614]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input573_I (.I(itasegm[615]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input574_I (.I(itasegm[616]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input575_I (.I(itasegm[617]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input576_I (.I(itasegm[618]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input577_I (.I(itasegm[619]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input578_I (.I(itasegm[61]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input579_I (.I(itasegm[620]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input57_I (.I(itasegm[150]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input580_I (.I(itasegm[621]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input581_I (.I(itasegm[622]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input582_I (.I(itasegm[623]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input583_I (.I(itasegm[624]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input584_I (.I(itasegm[625]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input585_I (.I(itasegm[626]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input586_I (.I(itasegm[627]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input587_I (.I(itasegm[628]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input588_I (.I(itasegm[629]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input589_I (.I(itasegm[62]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input58_I (.I(itasegm[151]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input590_I (.I(itasegm[630]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input591_I (.I(itasegm[631]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input592_I (.I(itasegm[632]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input593_I (.I(itasegm[633]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input594_I (.I(itasegm[634]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input595_I (.I(itasegm[635]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input596_I (.I(itasegm[636]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input597_I (.I(itasegm[637]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input598_I (.I(itasegm[638]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input599_I (.I(itasegm[639]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input59_I (.I(itasegm[152]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(itasegm[103]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input600_I (.I(itasegm[63]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input601_I (.I(itasegm[640]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input602_I (.I(itasegm[641]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input603_I (.I(itasegm[642]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input604_I (.I(itasegm[643]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input605_I (.I(itasegm[644]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input606_I (.I(itasegm[645]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input607_I (.I(itasegm[646]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input608_I (.I(itasegm[647]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input609_I (.I(itasegm[648]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input60_I (.I(itasegm[153]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input610_I (.I(itasegm[649]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input611_I (.I(itasegm[64]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input612_I (.I(itasegm[650]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input613_I (.I(itasegm[651]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input614_I (.I(itasegm[652]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input615_I (.I(itasegm[653]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input616_I (.I(itasegm[654]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input617_I (.I(itasegm[655]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input618_I (.I(itasegm[656]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input619_I (.I(itasegm[657]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input61_I (.I(itasegm[154]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input620_I (.I(itasegm[658]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input621_I (.I(itasegm[659]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input622_I (.I(itasegm[65]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input623_I (.I(itasegm[660]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input624_I (.I(itasegm[661]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input625_I (.I(itasegm[662]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input626_I (.I(itasegm[663]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input627_I (.I(itasegm[664]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input628_I (.I(itasegm[665]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input629_I (.I(itasegm[666]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input62_I (.I(itasegm[155]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input630_I (.I(itasegm[667]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input631_I (.I(itasegm[668]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input632_I (.I(itasegm[669]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input633_I (.I(itasegm[66]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input634_I (.I(itasegm[670]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input635_I (.I(itasegm[671]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input636_I (.I(itasegm[672]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input637_I (.I(itasegm[673]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input638_I (.I(itasegm[674]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input639_I (.I(itasegm[675]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input63_I (.I(itasegm[156]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input640_I (.I(itasegm[676]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input641_I (.I(itasegm[677]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input642_I (.I(itasegm[678]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input643_I (.I(itasegm[679]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input644_I (.I(itasegm[67]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input645_I (.I(itasegm[680]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input646_I (.I(itasegm[681]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input647_I (.I(itasegm[682]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input648_I (.I(itasegm[683]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input649_I (.I(itasegm[684]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input64_I (.I(itasegm[157]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input650_I (.I(itasegm[685]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input651_I (.I(itasegm[686]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input652_I (.I(itasegm[687]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input653_I (.I(itasegm[688]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input654_I (.I(itasegm[689]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input655_I (.I(itasegm[68]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input656_I (.I(itasegm[690]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input657_I (.I(itasegm[691]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input658_I (.I(itasegm[692]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input659_I (.I(itasegm[693]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input65_I (.I(itasegm[158]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input660_I (.I(itasegm[694]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input661_I (.I(itasegm[695]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input662_I (.I(itasegm[696]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input663_I (.I(itasegm[697]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input664_I (.I(itasegm[698]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input665_I (.I(itasegm[699]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input666_I (.I(itasegm[69]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input667_I (.I(itasegm[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input668_I (.I(itasegm[700]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input669_I (.I(itasegm[701]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input66_I (.I(itasegm[159]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input670_I (.I(itasegm[702]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input671_I (.I(itasegm[703]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input672_I (.I(itasegm[704]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input673_I (.I(itasegm[705]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input674_I (.I(itasegm[706]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input675_I (.I(itasegm[707]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input676_I (.I(itasegm[708]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input677_I (.I(itasegm[709]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input678_I (.I(itasegm[70]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input679_I (.I(itasegm[710]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input67_I (.I(itasegm[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input680_I (.I(itasegm[711]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input681_I (.I(itasegm[712]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input682_I (.I(itasegm[713]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input683_I (.I(itasegm[714]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input684_I (.I(itasegm[715]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input685_I (.I(itasegm[716]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input686_I (.I(itasegm[717]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input687_I (.I(itasegm[718]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input688_I (.I(itasegm[719]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input689_I (.I(itasegm[71]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input68_I (.I(itasegm[160]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input690_I (.I(itasegm[720]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input691_I (.I(itasegm[721]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input692_I (.I(itasegm[722]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input693_I (.I(itasegm[723]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input694_I (.I(itasegm[724]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input695_I (.I(itasegm[725]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input696_I (.I(itasegm[726]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input697_I (.I(itasegm[727]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input698_I (.I(itasegm[728]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input699_I (.I(itasegm[729]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input69_I (.I(itasegm[161]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(itasegm[104]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input700_I (.I(itasegm[72]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input701_I (.I(itasegm[730]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input702_I (.I(itasegm[731]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input703_I (.I(itasegm[732]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input704_I (.I(itasegm[733]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input705_I (.I(itasegm[734]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input706_I (.I(itasegm[735]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input707_I (.I(itasegm[736]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input708_I (.I(itasegm[737]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input709_I (.I(itasegm[738]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input70_I (.I(itasegm[162]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input710_I (.I(itasegm[739]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input711_I (.I(itasegm[73]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input712_I (.I(itasegm[740]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input713_I (.I(itasegm[741]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input714_I (.I(itasegm[742]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input715_I (.I(itasegm[743]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input716_I (.I(itasegm[744]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input717_I (.I(itasegm[745]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input718_I (.I(itasegm[746]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input719_I (.I(itasegm[747]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input71_I (.I(itasegm[163]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input720_I (.I(itasegm[748]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input721_I (.I(itasegm[749]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input722_I (.I(itasegm[74]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input723_I (.I(itasegm[750]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input724_I (.I(itasegm[751]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input725_I (.I(itasegm[752]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input726_I (.I(itasegm[753]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input727_I (.I(itasegm[754]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input728_I (.I(itasegm[755]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input729_I (.I(itasegm[756]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input72_I (.I(itasegm[164]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input730_I (.I(itasegm[757]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input731_I (.I(itasegm[758]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input732_I (.I(itasegm[759]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input733_I (.I(itasegm[75]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input734_I (.I(itasegm[760]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input735_I (.I(itasegm[761]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input736_I (.I(itasegm[762]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input737_I (.I(itasegm[763]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input738_I (.I(itasegm[764]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input739_I (.I(itasegm[765]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input73_I (.I(itasegm[165]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input740_I (.I(itasegm[766]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input741_I (.I(itasegm[767]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input742_I (.I(itasegm[768]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input743_I (.I(itasegm[769]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input744_I (.I(itasegm[76]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input745_I (.I(itasegm[770]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input746_I (.I(itasegm[771]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input747_I (.I(itasegm[772]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input748_I (.I(itasegm[773]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input749_I (.I(itasegm[774]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input74_I (.I(itasegm[166]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input750_I (.I(itasegm[775]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input751_I (.I(itasegm[776]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input752_I (.I(itasegm[777]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input753_I (.I(itasegm[778]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input754_I (.I(itasegm[779]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input755_I (.I(itasegm[77]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input756_I (.I(itasegm[780]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input757_I (.I(itasegm[781]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input758_I (.I(itasegm[782]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input759_I (.I(itasegm[783]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input75_I (.I(itasegm[167]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input760_I (.I(itasegm[784]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input761_I (.I(itasegm[785]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input762_I (.I(itasegm[786]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input763_I (.I(itasegm[787]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input764_I (.I(itasegm[788]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input765_I (.I(itasegm[789]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input766_I (.I(itasegm[78]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input767_I (.I(itasegm[790]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input768_I (.I(itasegm[791]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input769_I (.I(itasegm[792]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input76_I (.I(itasegm[168]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input770_I (.I(itasegm[793]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input771_I (.I(itasegm[794]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input772_I (.I(itasegm[795]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input773_I (.I(itasegm[796]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input774_I (.I(itasegm[797]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input775_I (.I(itasegm[798]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input776_I (.I(itasegm[799]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input777_I (.I(itasegm[79]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input778_I (.I(itasegm[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input779_I (.I(itasegm[800]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input77_I (.I(itasegm[169]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input780_I (.I(itasegm[801]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input781_I (.I(itasegm[802]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input782_I (.I(itasegm[803]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input783_I (.I(itasegm[804]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input784_I (.I(itasegm[805]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input785_I (.I(itasegm[806]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input786_I (.I(itasegm[807]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input787_I (.I(itasegm[808]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input788_I (.I(itasegm[809]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input789_I (.I(itasegm[80]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input78_I (.I(itasegm[16]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input790_I (.I(itasegm[810]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input791_I (.I(itasegm[811]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input792_I (.I(itasegm[812]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input793_I (.I(itasegm[813]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input794_I (.I(itasegm[814]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input795_I (.I(itasegm[815]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input796_I (.I(itasegm[816]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input797_I (.I(itasegm[817]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input798_I (.I(itasegm[818]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input799_I (.I(itasegm[819]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input79_I (.I(itasegm[170]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input7_I (.I(itasegm[105]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input800_I (.I(itasegm[81]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input801_I (.I(itasegm[820]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input802_I (.I(itasegm[821]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input803_I (.I(itasegm[822]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input804_I (.I(itasegm[823]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input805_I (.I(itasegm[824]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input806_I (.I(itasegm[825]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input807_I (.I(itasegm[826]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input808_I (.I(itasegm[827]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input809_I (.I(itasegm[828]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input80_I (.I(itasegm[171]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input810_I (.I(itasegm[829]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input811_I (.I(itasegm[82]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input812_I (.I(itasegm[830]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input813_I (.I(itasegm[831]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input814_I (.I(itasegm[832]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input815_I (.I(itasegm[833]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input816_I (.I(itasegm[834]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input817_I (.I(itasegm[835]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input818_I (.I(itasegm[836]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input819_I (.I(itasegm[837]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input81_I (.I(itasegm[172]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input820_I (.I(itasegm[838]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input821_I (.I(itasegm[839]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input822_I (.I(itasegm[83]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input823_I (.I(itasegm[840]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input824_I (.I(itasegm[841]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input825_I (.I(itasegm[842]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input826_I (.I(itasegm[843]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input827_I (.I(itasegm[844]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input828_I (.I(itasegm[845]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input829_I (.I(itasegm[846]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input82_I (.I(itasegm[173]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input830_I (.I(itasegm[847]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input831_I (.I(itasegm[848]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input832_I (.I(itasegm[849]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input833_I (.I(itasegm[84]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input834_I (.I(itasegm[850]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input835_I (.I(itasegm[851]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input836_I (.I(itasegm[852]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input837_I (.I(itasegm[853]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input838_I (.I(itasegm[854]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input839_I (.I(itasegm[855]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input83_I (.I(itasegm[174]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input840_I (.I(itasegm[856]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input841_I (.I(itasegm[857]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input842_I (.I(itasegm[858]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input843_I (.I(itasegm[859]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input844_I (.I(itasegm[85]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input845_I (.I(itasegm[860]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input846_I (.I(itasegm[861]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input847_I (.I(itasegm[862]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input848_I (.I(itasegm[863]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input849_I (.I(itasegm[864]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input84_I (.I(itasegm[175]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input850_I (.I(itasegm[865]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input851_I (.I(itasegm[866]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input852_I (.I(itasegm[867]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input853_I (.I(itasegm[868]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input854_I (.I(itasegm[869]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input855_I (.I(itasegm[86]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input856_I (.I(itasegm[870]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input857_I (.I(itasegm[871]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input858_I (.I(itasegm[872]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input859_I (.I(itasegm[873]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input85_I (.I(itasegm[176]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input860_I (.I(itasegm[874]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input861_I (.I(itasegm[875]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input862_I (.I(itasegm[876]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input863_I (.I(itasegm[877]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input864_I (.I(itasegm[878]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input865_I (.I(itasegm[879]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input866_I (.I(itasegm[87]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input867_I (.I(itasegm[880]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input868_I (.I(itasegm[881]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input869_I (.I(itasegm[882]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input86_I (.I(itasegm[177]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input870_I (.I(itasegm[883]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input871_I (.I(itasegm[884]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input872_I (.I(itasegm[885]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input873_I (.I(itasegm[886]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input874_I (.I(itasegm[887]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input875_I (.I(itasegm[888]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input876_I (.I(itasegm[889]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input877_I (.I(itasegm[88]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input878_I (.I(itasegm[890]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input879_I (.I(itasegm[891]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input87_I (.I(itasegm[178]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input880_I (.I(itasegm[892]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input881_I (.I(itasegm[893]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input882_I (.I(itasegm[894]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input883_I (.I(itasegm[895]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input884_I (.I(itasegm[89]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input885_I (.I(itasegm[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input886_I (.I(itasegm[90]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input887_I (.I(itasegm[91]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input888_I (.I(itasegm[92]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input889_I (.I(itasegm[93]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input88_I (.I(itasegm[179]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input890_I (.I(itasegm[94]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input891_I (.I(itasegm[95]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input892_I (.I(itasegm[96]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input893_I (.I(itasegm[97]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input894_I (.I(itasegm[98]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input895_I (.I(itasegm[99]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input896_I (.I(itasegm[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input897_I (.I(itasel[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input898_I (.I(itasel[100]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input899_I (.I(itasel[101]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input89_I (.I(itasegm[17]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input8_I (.I(itasegm[106]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input900_I (.I(itasel[102]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input901_I (.I(itasel[103]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input902_I (.I(itasel[104]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input903_I (.I(itasel[105]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input904_I (.I(itasel[106]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input905_I (.I(itasel[107]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input906_I (.I(itasel[108]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input907_I (.I(itasel[109]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input908_I (.I(itasel[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input909_I (.I(itasel[110]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input90_I (.I(itasegm[180]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input910_I (.I(itasel[111]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input911_I (.I(itasel[112]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input912_I (.I(itasel[113]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input913_I (.I(itasel[114]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input914_I (.I(itasel[115]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input915_I (.I(itasel[116]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input916_I (.I(itasel[117]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input917_I (.I(itasel[118]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input918_I (.I(itasel[119]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input919_I (.I(itasel[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input91_I (.I(itasegm[181]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input920_I (.I(itasel[120]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input921_I (.I(itasel[121]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input922_I (.I(itasel[122]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input923_I (.I(itasel[123]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input924_I (.I(itasel[124]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input925_I (.I(itasel[125]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input926_I (.I(itasel[126]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input927_I (.I(itasel[127]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input928_I (.I(itasel[128]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input929_I (.I(itasel[129]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input92_I (.I(itasegm[182]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input930_I (.I(itasel[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input931_I (.I(itasel[130]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input932_I (.I(itasel[131]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input933_I (.I(itasel[132]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input934_I (.I(itasel[133]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input935_I (.I(itasel[134]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input936_I (.I(itasel[135]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input937_I (.I(itasel[136]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input938_I (.I(itasel[137]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input939_I (.I(itasel[138]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input93_I (.I(itasegm[183]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input940_I (.I(itasel[139]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input941_I (.I(itasel[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input942_I (.I(itasel[140]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input943_I (.I(itasel[141]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input944_I (.I(itasel[142]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input945_I (.I(itasel[143]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input946_I (.I(itasel[144]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input947_I (.I(itasel[145]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input948_I (.I(itasel[146]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input949_I (.I(itasel[147]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input94_I (.I(itasegm[184]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input950_I (.I(itasel[148]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input951_I (.I(itasel[149]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input952_I (.I(itasel[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input953_I (.I(itasel[150]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input954_I (.I(itasel[151]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input955_I (.I(itasel[152]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input956_I (.I(itasel[153]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input957_I (.I(itasel[154]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input958_I (.I(itasel[155]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input959_I (.I(itasel[156]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input95_I (.I(itasegm[185]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input960_I (.I(itasel[157]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input961_I (.I(itasel[158]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input962_I (.I(itasel[159]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input963_I (.I(itasel[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input964_I (.I(itasel[160]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input965_I (.I(itasel[161]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input966_I (.I(itasel[162]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input967_I (.I(itasel[163]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input968_I (.I(itasel[164]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input969_I (.I(itasel[165]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input96_I (.I(itasegm[186]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input970_I (.I(itasel[166]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input971_I (.I(itasel[167]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input972_I (.I(itasel[168]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input973_I (.I(itasel[169]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input974_I (.I(itasel[16]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input975_I (.I(itasel[170]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input976_I (.I(itasel[171]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input977_I (.I(itasel[172]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input978_I (.I(itasel[173]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input979_I (.I(itasel[174]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input97_I (.I(itasegm[187]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input980_I (.I(itasel[175]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input981_I (.I(itasel[176]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input982_I (.I(itasel[177]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input983_I (.I(itasel[178]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input984_I (.I(itasel[179]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input985_I (.I(itasel[17]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input986_I (.I(itasel[180]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input987_I (.I(itasel[181]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input988_I (.I(itasel[182]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input989_I (.I(itasel[183]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input98_I (.I(itasegm[188]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input990_I (.I(itasel[184]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input991_I (.I(itasel[185]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input992_I (.I(itasel[186]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input993_I (.I(itasel[187]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input994_I (.I(itasel[188]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input995_I (.I(itasel[189]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input996_I (.I(itasel[18]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input997_I (.I(itasel[190]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input998_I (.I(itasel[191]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input999_I (.I(itasel[192]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input99_I (.I(itasegm[189]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input9_I (.I(itasegm[107]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output1673_I (.I(net1673));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output1674_I (.I(net1674));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output1675_I (.I(net1675));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output1682_I (.I(net1682));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output1684_I (.I(net1684));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output1685_I (.I(net1685));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output1686_I (.I(net1686));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output1687_I (.I(net1687));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output1688_I (.I(net1688));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output1689_I (.I(net1689));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output1690_I (.I(net1690));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output1691_I (.I(net1691));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output1692_I (.I(net1692));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output1693_I (.I(net1693));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output1694_I (.I(net1694));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output1695_I (.I(net1695));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output1696_I (.I(net1696));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1699_I (.I(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1700_I (.I(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1704_I (.I(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1706_I (.I(net1707));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1707_I (.I(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1708_I (.I(net1709));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1709_I (.I(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1710_I (.I(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1712_I (.I(net1713));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1713_I (.I(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1714_I (.I(net1715));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1715_I (.I(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1716_I (.I(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1717_I (.I(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1718_I (.I(net1719));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1719_I (.I(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1720_I (.I(net1721));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1721_I (.I(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1722_I (.I(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1724_I (.I(net1725));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1725_I (.I(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1726_I (.I(net1727));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1727_I (.I(_0606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1728_I (.I(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1729_I (.I(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1730_I (.I(net1731));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1731_I (.I(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1732_I (.I(net1733));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1733_I (.I(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1734_I (.I(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1735_I (.I(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1736_I (.I(net1737));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1737_I (.I(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1738_I (.I(net1739));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1739_I (.I(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1740_I (.I(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1742_I (.I(net1743));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1743_I (.I(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1744_I (.I(net1745));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1745_I (.I(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1746_I (.I(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1747_I (.I(_0276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1748_I (.I(net1749));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1749_I (.I(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1750_I (.I(net1751));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1751_I (.I(_0225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1752_I (.I(_0144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1753_I (.I(_2174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1754_I (.I(_2166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1755_I (.I(_2162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1756_I (.I(_2113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1757_I (.I(_2105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1758_I (.I(_2100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1759_I (.I(_2048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1760_I (.I(_2040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1761_I (.I(_2036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1762_I (.I(_1971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1763_I (.I(_1955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1764_I (.I(_1947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1765_I (.I(_1856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1766_I (.I(_1848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1767_I (.I(_1844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1768_I (.I(_1795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1769_I (.I(_1787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1770_I (.I(_1782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1771_I (.I(_1730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1772_I (.I(_1722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1773_I (.I(_1718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1774_I (.I(_1694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1776_I (.I(_1653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1777_I (.I(_1637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1778_I (.I(_1629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1779_I (.I(net1780));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1780_I (.I(_1530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1781_I (.I(net1782));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1782_I (.I(_1526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1783_I (.I(_1502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1784_I (.I(_1498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1785_I (.I(net1786));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1786_I (.I(_1469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1787_I (.I(net1788));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1788_I (.I(_1464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1789_I (.I(_1438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1790_I (.I(_1434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1791_I (.I(net1792));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1792_I (.I(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1793_I (.I(net1794));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1794_I (.I(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1795_I (.I(net1796));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1796_I (.I(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1797_I (.I(net1798));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1798_I (.I(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1799_I (.I(net1800));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1800_I (.I(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1801_I (.I(net1802));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1802_I (.I(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1803_I (.I(net1804));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1804_I (.I(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1805_I (.I(net1806));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1806_I (.I(_1145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1807_I (.I(net1808));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1808_I (.I(_1085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1809_I (.I(net1810));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1810_I (.I(_1081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1811_I (.I(net1812));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1812_I (.I(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1813_I (.I(net1814));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1814_I (.I(_0964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1815_I (.I(_2296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1816_I (.I(_2288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1817_I (.I(_2284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1818_I (.I(_2270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1820_I (.I(_2227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1821_I (.I(_2223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1822_I (.I(_2209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1824_I (.I(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1825_I (.I(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1826_I (.I(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_100_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_100_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_100_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_100_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_100_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_100_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_101_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_101_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_101_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_101_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_101_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_101_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_102_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_102_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_102_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_102_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_103_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_103_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_103_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_103_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_103_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_103_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_104_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_104_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_104_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_104_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_104_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_104_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_104_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_105_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_105_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_105_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_105_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_105_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_106_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_106_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_106_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_106_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_106_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_107_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_107_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_107_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_107_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_108_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_108_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_108_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_108_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_108_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_108_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_108_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_109_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_109_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_109_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_109_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_109_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_110_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_110_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_110_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_110_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_111_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_111_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_111_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_111_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_111_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_111_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_112_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_112_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_112_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_112_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_112_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_112_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_113_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_113_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_113_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_113_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_113_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_114_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_114_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_114_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_115_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_115_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_115_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_115_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_116_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_116_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_116_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_116_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_116_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_116_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_117_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_117_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_117_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_117_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_117_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_117_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_118_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_118_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_118_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_118_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_118_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_118_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_119_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_119_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_119_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_119_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_119_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_119_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_119_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_120_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_120_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_120_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_120_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_121_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_121_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_121_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_121_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_121_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_121_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_122_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_122_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_122_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_122_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_122_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_123_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_123_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_123_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_123_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_123_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_123_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_123_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_123_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_123_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_124_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_124_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_124_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_124_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_124_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_125_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_125_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_125_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_125_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_125_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_126_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_126_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_126_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_126_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_127_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_127_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_127_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_127_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_127_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_128_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_128_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_128_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_128_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_128_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_128_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_129_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_129_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_129_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_129_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_129_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_129_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_129_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_130_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_130_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_130_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_130_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_130_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_130_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_130_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_131_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_131_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_131_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_131_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_131_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_131_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_131_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_132_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_132_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_132_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_132_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_132_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_133_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_133_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_133_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_133_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_133_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_133_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_134_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_134_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_134_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_134_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_134_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_134_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_134_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_134_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_135_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_135_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_135_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_135_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_135_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_135_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_135_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_135_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_135_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_135_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_136_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_136_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_136_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_137_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_137_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_138_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_138_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_138_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_138_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_138_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_139_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_139_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_139_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_139_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_13_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_140_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_140_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_140_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_140_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_140_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_141_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_141_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_141_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_141_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_142_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_142_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_142_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_142_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_142_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_143_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_143_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_143_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_144_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_144_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_144_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_144_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_144_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_144_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_144_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_145_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_145_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_145_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_145_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_145_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_145_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_146_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_146_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_146_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_146_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_146_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_146_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_146_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_146_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_146_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_147_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_147_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_147_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_147_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_147_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_147_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_147_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_147_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_148_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_148_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_148_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_148_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_148_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_148_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_148_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_148_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_148_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_148_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_149_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_149_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_149_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_149_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_149_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_149_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_149_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_150_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_150_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_151_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_151_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_151_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_151_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_151_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_151_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_151_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_152_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_152_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_152_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_152_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_152_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_152_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_153_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_153_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_153_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_153_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_153_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_153_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_153_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_153_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_153_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_153_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_153_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_153_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_153_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_153_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_153_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_154_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_154_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_154_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_154_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_154_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_154_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_154_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_154_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_154_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_154_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_155_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_155_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_155_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_156_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_156_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_156_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_156_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_156_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_157_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_157_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_157_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_157_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_157_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_157_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_158_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_158_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_158_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_158_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_158_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_158_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_158_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_159_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_159_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_159_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_159_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_159_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_159_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_159_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_15_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_15_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_160_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_160_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_160_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_160_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_160_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_160_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_160_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_161_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_161_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_161_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_161_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_162_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_162_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_162_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_162_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_162_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_162_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_162_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_162_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_162_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_163_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_163_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_163_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_163_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_163_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_163_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_163_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_163_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_163_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_163_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_163_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_163_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_163_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_163_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_163_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_163_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_164_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_164_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_164_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_164_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_164_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_164_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_164_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_164_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_164_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_164_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_164_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_164_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_164_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_165_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_165_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_165_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_165_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_165_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_165_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_165_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_165_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_165_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_165_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_165_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_165_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_165_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_165_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_165_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_165_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_165_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_165_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_166_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_166_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_166_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_166_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_166_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_166_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_166_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_166_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_166_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_166_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_166_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_166_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_166_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_166_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_166_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_166_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_167_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_167_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_167_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_167_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_167_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_167_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_167_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_167_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_167_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_167_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_167_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_167_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_168_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_169_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_169_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_169_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_169_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_169_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_169_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_169_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_169_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_169_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_16_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_16_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_170_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_170_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_170_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_170_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_170_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_170_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_170_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_170_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_170_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_170_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_170_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_170_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_170_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_170_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_170_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_170_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_170_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_171_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_171_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_171_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_171_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_171_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_171_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_171_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_171_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_171_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_171_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_171_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_171_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_171_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_171_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_172_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_172_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_172_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_172_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_172_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_172_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_172_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_172_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_172_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_172_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_172_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_172_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_172_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_172_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_172_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_172_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_173_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_173_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_173_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_173_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_173_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_173_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_173_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_173_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_173_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_173_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_173_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_173_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_173_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_173_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_173_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_173_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_173_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_173_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_173_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_173_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_173_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_173_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_174_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_174_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_174_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_174_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_174_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_174_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_174_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_174_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_174_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_174_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_174_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_174_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_174_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_174_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_174_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_174_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_175_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_175_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_175_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_175_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_175_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_175_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_175_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_175_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_175_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_175_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_175_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_175_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_175_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_175_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_175_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_175_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_175_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_175_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_175_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_175_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_175_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_175_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_175_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_175_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_175_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_175_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_175_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_175_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_175_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_176_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_176_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_176_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_176_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_176_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_176_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_176_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_176_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_176_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_176_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_176_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_176_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_176_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_176_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_176_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_177_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_177_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_177_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_177_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_177_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_177_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_177_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_177_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_177_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_177_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_177_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_177_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_177_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_177_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_178_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_178_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_178_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_178_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_178_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_178_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_178_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_178_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_178_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_178_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_178_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_178_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_178_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_178_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_178_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_178_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_179_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_179_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_179_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_179_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_179_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_179_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_179_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_179_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_179_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_179_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_179_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_179_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_179_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_179_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_179_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_179_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_179_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_179_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_180_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_180_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_180_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_180_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_180_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_180_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_180_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_180_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_180_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_180_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_180_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_180_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_180_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_181_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_181_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_181_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_181_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_181_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_181_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_181_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_181_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_181_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_181_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_181_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_181_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_181_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_181_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_181_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_181_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_181_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_181_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_181_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_181_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_181_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_181_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_182_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_182_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_182_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_182_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_182_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_182_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_182_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_182_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_182_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_182_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_182_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_182_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_182_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_182_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_182_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_182_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_183_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_183_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_183_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_183_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_183_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_183_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_183_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_183_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_183_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_183_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_183_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_183_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_183_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_183_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_183_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_183_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_183_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_183_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_183_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_183_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_183_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_183_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_183_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_183_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_183_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_183_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_183_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_183_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_183_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_183_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_183_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_183_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_183_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_183_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_183_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_183_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_183_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_183_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_183_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_183_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_183_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_183_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_183_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_183_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_183_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_184_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_184_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_184_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_184_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_184_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_184_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_184_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_184_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_184_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_184_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_184_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_184_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_184_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_184_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_184_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_184_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_184_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_184_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_184_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_184_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_184_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_184_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_184_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_184_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_184_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_184_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_184_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_184_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_184_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_184_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_184_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_184_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_184_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_184_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_184_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_184_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_184_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_184_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_184_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_184_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_184_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_184_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_184_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_184_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_184_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_185_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_185_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_185_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_185_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_185_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_185_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_185_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_185_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_185_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_185_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_185_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_185_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_185_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_185_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_185_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_185_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_185_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_185_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_185_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_185_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_185_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_185_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_185_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_185_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_185_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_185_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_185_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_185_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_185_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_185_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_185_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_185_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_185_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_185_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_186_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_186_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_186_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_186_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_186_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_186_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_186_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_186_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_186_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_186_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_186_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_186_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_186_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_186_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_186_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_186_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_186_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_186_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_186_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_186_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_186_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_186_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_186_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_186_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_186_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_186_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_186_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_186_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_186_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_186_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_186_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_186_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_186_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_186_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_186_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_186_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_186_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_186_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_187_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_187_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_187_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_187_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_187_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_187_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_187_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_187_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_187_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_187_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_187_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_187_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_187_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_187_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_187_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_187_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_187_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_187_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_187_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_187_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_187_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_187_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_187_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_187_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_187_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_187_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_187_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_187_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_187_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_187_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_188_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_188_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_188_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_188_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_188_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_188_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_188_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_188_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_188_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_188_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_188_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_188_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_188_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_188_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_188_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_188_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_188_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_188_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_188_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_188_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_189_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_189_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_189_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_189_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_189_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_189_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_189_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_189_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_189_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_189_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_189_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_189_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_189_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_189_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_189_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_189_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_189_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_189_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_189_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_189_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_189_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_189_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_189_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_190_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_190_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_190_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_190_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_190_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_190_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_190_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_190_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_190_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_190_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_190_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_190_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_190_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_190_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_190_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_190_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_190_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_190_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_190_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_190_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_190_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_190_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_190_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_190_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_191_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_191_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_191_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_191_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_191_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_191_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_191_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_191_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_191_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_191_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_191_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_191_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_191_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_191_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_191_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_191_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_191_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_191_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_191_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_191_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_191_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_191_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_191_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_191_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_191_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_191_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_191_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_191_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_191_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_192_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_192_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_192_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_192_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_192_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_192_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_192_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_192_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_192_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_192_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_192_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_192_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_192_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_192_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_192_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_192_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_192_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_192_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_192_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_192_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_192_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_192_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_192_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_192_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_192_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_192_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_192_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_193_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_193_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_193_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_193_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_193_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_193_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_193_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_193_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_193_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_193_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_193_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_193_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_193_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_193_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_193_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_193_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_193_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_193_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_193_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_193_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_193_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_193_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_193_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_193_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_193_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_193_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_193_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_193_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_193_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_193_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_193_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_193_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_193_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_193_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_193_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_193_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_193_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_193_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_193_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_193_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_193_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_193_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_193_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_193_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_193_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_194_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_194_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_194_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_194_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_194_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_194_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_194_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_194_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_194_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_194_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_194_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_194_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_194_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_194_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_194_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_194_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_194_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_194_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_194_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_194_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_194_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_194_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_194_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_194_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_195_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_195_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_195_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_195_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_195_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_195_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_195_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_195_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_195_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_195_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_196_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_196_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_196_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_196_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_196_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_196_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_196_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_196_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_196_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_196_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_196_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_196_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_196_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_196_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_196_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_196_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_196_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_196_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_196_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_196_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_196_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_196_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_196_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_196_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_196_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_196_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_196_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_196_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_196_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_196_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_196_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_196_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_196_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_196_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_196_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_196_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_196_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_196_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_196_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_197_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_197_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_197_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_197_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_197_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_197_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_197_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_197_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_197_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_197_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_197_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_197_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_197_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_197_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_197_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_197_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_197_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_197_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_197_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_197_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_197_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_197_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_197_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_197_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_197_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_197_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_197_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_197_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_197_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_197_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_198_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_198_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_198_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_198_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_198_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_198_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_198_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_198_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_198_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_198_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_198_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_198_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_198_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_198_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_198_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_198_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_198_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_198_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_198_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_198_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_198_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_198_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_198_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_198_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_198_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_198_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_198_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_199_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_199_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_199_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_199_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_199_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_199_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_199_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_199_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_199_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_199_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_199_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_199_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_199_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_199_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_199_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_199_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_199_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_199_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_199_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_199_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_199_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_199_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_199_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_199_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_199_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_199_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_199_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_199_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_199_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_19_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_200_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_200_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_200_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_200_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_200_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_200_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_200_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_200_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_200_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_200_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_200_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_200_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_200_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_200_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_200_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_200_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_200_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_200_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_200_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_200_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_200_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_200_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_200_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_200_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_200_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_200_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_200_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_200_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_200_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_200_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_200_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_200_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_201_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_201_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_201_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_201_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_201_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_201_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_201_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_201_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_201_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_201_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_201_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_201_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_201_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_201_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_201_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_201_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_201_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_201_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_201_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_201_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_201_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_201_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_201_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_201_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_201_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_201_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_202_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_202_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_202_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_202_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_202_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_202_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_202_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_202_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_202_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_202_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_202_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_202_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_202_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_202_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_202_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_202_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_202_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_202_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_202_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_202_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_202_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_202_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_202_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_202_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_202_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_202_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_202_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_202_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_202_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_202_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_202_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_202_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_202_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_202_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_202_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_202_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_202_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_202_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_202_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_202_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_202_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_202_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_202_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_202_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_202_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_202_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_203_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_203_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_203_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_203_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_203_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_203_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_203_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_203_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_203_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_203_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_203_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_203_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_203_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_203_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_203_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_203_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_203_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_203_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_203_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_203_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_203_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_203_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_203_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_203_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_203_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_203_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_203_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_203_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_203_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_203_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_203_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_203_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_203_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_203_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_204_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_204_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_204_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_204_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_204_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_204_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_204_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_204_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_204_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_204_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_204_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_204_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_204_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_204_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_204_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_204_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_204_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_204_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_204_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_204_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_204_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_204_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_204_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_204_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_204_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_204_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_204_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_204_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_204_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_204_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_204_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_204_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_204_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_204_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_204_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_204_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_205_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_205_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_205_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_205_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_205_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_205_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_205_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_205_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_205_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_205_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_205_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_205_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_205_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_205_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_205_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_205_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_205_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_205_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_205_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_205_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_205_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_205_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_205_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_205_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_205_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_205_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_205_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_205_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_205_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_205_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_205_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_205_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_205_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_205_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_205_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_205_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_205_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_205_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_205_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_205_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_205_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_206_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_206_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_206_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_206_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_206_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_206_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_206_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_206_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_206_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_206_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_206_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_206_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_206_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_206_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_206_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_206_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_206_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_206_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_206_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_206_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_206_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_206_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_206_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_206_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_206_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_206_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_206_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_206_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_206_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_206_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_206_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_206_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_207_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_207_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_207_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_207_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_207_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_207_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_207_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_207_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_207_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_207_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_207_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_207_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_207_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_207_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_207_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_207_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_207_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_207_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_207_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_207_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_207_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_207_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_207_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_207_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_207_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_207_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_207_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_207_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_207_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_207_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_207_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_207_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_207_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_207_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_207_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_207_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_207_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_208_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_208_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_208_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_208_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_208_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_208_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_208_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_208_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_208_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_208_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_208_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_208_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_208_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_208_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_208_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_208_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_208_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_208_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_208_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_208_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_208_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_208_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_208_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_209_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_209_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_209_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_209_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_209_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_209_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_209_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_209_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_209_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_209_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_209_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_209_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_209_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_209_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_209_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_209_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_209_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_209_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_209_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_209_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_209_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_209_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_209_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_209_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_209_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_209_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_209_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_209_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_209_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_209_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_210_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_210_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_210_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_210_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_210_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_210_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_210_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_210_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_210_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_210_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_210_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_210_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_210_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_210_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_210_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_210_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_210_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_210_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_210_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_210_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_210_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_210_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_210_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_210_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_210_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_210_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_210_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_210_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_211_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_211_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_211_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_211_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_211_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_211_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_211_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_211_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_211_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_211_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_211_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_211_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_211_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_211_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_211_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_211_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_211_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_211_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_211_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_211_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_211_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_211_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_211_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_211_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_211_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_211_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_211_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_211_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_211_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_211_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_211_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_212_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_212_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_212_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_212_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_212_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_212_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_212_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_212_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_212_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_212_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_212_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_212_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_212_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_212_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_212_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_212_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_212_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_212_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_212_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_212_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_212_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_212_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_212_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_212_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_212_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_212_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_212_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_212_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_212_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_212_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_212_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_212_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_212_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_212_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_212_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_212_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_212_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_212_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_212_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_213_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_213_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_213_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_213_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_213_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_213_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_213_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_213_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_213_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_213_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_213_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_213_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_213_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_213_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_213_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_213_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_213_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_213_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_213_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_213_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_213_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_213_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_213_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_213_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_213_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_213_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_213_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_213_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_213_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_213_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_213_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_214_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_214_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_214_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_214_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_214_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_214_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_214_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_214_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_214_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_214_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_214_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_214_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_214_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_214_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_214_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_214_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_214_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_214_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_214_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_214_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_214_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_214_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_214_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_214_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_214_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_214_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_214_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_214_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_214_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_214_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_214_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_214_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_214_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_214_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_214_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_214_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_214_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_214_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_214_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_214_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_215_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_215_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_215_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_215_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_215_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_215_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_215_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_215_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_215_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_215_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_215_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_215_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_215_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_215_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_215_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_215_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_215_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_215_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_215_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_215_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_215_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_215_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_215_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_215_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_215_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_215_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_215_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_215_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_215_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_216_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_216_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_216_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_216_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_216_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_216_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_216_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_216_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_216_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_216_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_216_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_216_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_216_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_216_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_216_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_216_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_216_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_216_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_216_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_216_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_216_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_216_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_216_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_216_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_216_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_216_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_216_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_216_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_216_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_216_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_216_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_216_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_216_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_216_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_216_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_216_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_217_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_217_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_217_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_217_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_217_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_217_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_217_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_217_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_217_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_217_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_217_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_217_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_217_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_217_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_217_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_217_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_217_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_217_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_217_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_217_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_217_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_217_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_217_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_217_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_217_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_217_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_217_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_217_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_217_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_217_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_217_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_217_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_217_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_217_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_218_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_218_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_218_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_218_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_218_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_218_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_218_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_218_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_218_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_218_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_218_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_218_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_218_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_218_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_218_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_218_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_218_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_218_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_218_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_218_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_218_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_218_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_218_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_218_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_218_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_218_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_218_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_218_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_218_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_218_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_218_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_218_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_218_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_218_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_218_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_218_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_218_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_219_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_219_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_219_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_219_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_219_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_219_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_219_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_219_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_219_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_219_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_219_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_219_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_219_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_219_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_219_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_219_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_219_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_219_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_219_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_219_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_219_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_21_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_220_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_220_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_220_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_220_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_220_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_220_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_220_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_220_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_220_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_220_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_220_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_220_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_220_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_220_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_220_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_220_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_220_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_220_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_220_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_220_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_220_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_220_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_221_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_221_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_221_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_221_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_221_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_221_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_221_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_221_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_221_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_221_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_221_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_221_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_221_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_221_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_221_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_221_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_221_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_221_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_221_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_221_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_221_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_221_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_221_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_221_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_221_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_221_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_221_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_221_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_221_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_221_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_221_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_221_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_221_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_221_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_221_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_221_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_221_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_221_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_222_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_222_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_222_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_222_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_222_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_222_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_222_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_222_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_222_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_222_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_222_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_222_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_222_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_222_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_222_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_222_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_222_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_222_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_222_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_222_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_222_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_222_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_222_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_222_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_222_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_222_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_222_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_222_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_222_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_222_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_222_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_222_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_222_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_222_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_223_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_223_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_223_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_223_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_223_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_223_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_223_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_223_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_223_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_223_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_223_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_223_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_223_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_223_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_223_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_223_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_223_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_223_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_223_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_223_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_223_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_223_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_223_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_223_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_223_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_223_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_223_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_223_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_223_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_223_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_223_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_223_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_223_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_223_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_223_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_223_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_223_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_223_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_224_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_224_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_224_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_224_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_224_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_224_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_224_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_224_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_224_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_224_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_224_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_224_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_224_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_224_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_224_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_224_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_224_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_224_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_224_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_224_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_224_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_224_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_224_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_224_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_224_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_224_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_224_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_224_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_224_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_224_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_224_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_224_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_224_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_224_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_224_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_224_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_225_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_225_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_225_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_225_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_225_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_225_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_225_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_225_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_225_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_225_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_225_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_225_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_225_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_225_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_225_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_225_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_225_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_225_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_225_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_225_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_225_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_225_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_225_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_225_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_225_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_225_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_225_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_225_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_225_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_225_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_225_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_225_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_225_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_226_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_226_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_226_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_226_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_226_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_226_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_226_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_226_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_226_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_226_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_226_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_226_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_226_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_226_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_226_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_226_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_226_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_226_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_226_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_226_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_226_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_226_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_226_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_226_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_226_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_226_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_226_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_226_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_226_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_226_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_226_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_226_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_226_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_227_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_227_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_227_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_227_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_227_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_227_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_227_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_227_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_227_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_227_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_227_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_227_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_227_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_227_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_227_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_227_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_227_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_227_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_227_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_227_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_227_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_227_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_227_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_227_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_227_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_227_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_227_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_227_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_227_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_227_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_227_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_227_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_227_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_227_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_227_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_227_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_227_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_227_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_227_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_227_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_228_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_228_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_228_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_228_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_228_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_228_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_228_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_228_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_228_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_228_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_228_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_228_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_228_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_228_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_228_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_228_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_228_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_228_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_228_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_228_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_228_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_228_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_228_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_228_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_228_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_228_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_228_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_228_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_228_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_228_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_229_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_229_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_229_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_229_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_229_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_229_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_229_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_229_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_229_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_229_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_229_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_229_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_229_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_229_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_229_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_229_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_229_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_229_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_229_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_229_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_229_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_229_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_229_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_229_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_229_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_229_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_229_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_229_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_229_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_229_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_229_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_229_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_229_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_229_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_229_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_229_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_229_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_229_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_230_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_230_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_230_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_230_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_230_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_230_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_230_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_230_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_230_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_230_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_230_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_230_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_230_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_230_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_230_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_230_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_230_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_230_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_230_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_230_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_230_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_230_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_230_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_230_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_230_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_230_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_230_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_230_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_230_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_230_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_231_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_231_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_231_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_231_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_231_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_231_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_231_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_231_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_231_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_231_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_231_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_231_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_231_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_231_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_231_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_231_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_231_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_231_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_231_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_231_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_231_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_231_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_231_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_231_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_231_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_231_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_231_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_231_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_231_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_231_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_231_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_231_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_232_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_232_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_232_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_232_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_232_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_232_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_232_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_232_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_232_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_232_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_232_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_232_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_232_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_232_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_232_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_232_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_232_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_232_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_232_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_232_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_232_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_232_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_232_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_232_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_232_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_232_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_232_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_232_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_232_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_232_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_233_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_233_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_233_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_233_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_233_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_233_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_233_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_233_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_233_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_233_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_233_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_233_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_233_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_233_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_233_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_233_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_233_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_233_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_233_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_233_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_233_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_233_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_233_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_233_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_233_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_233_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_233_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_233_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_233_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_233_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_233_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_233_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_233_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_233_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_233_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_234_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_234_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_234_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_234_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_234_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_234_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_234_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_234_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_234_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_234_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_234_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_234_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_234_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_234_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_234_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_234_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_234_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_234_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_234_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_234_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_234_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_234_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_234_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_234_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_234_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_234_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_234_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_234_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_234_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_234_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_234_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_235_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_235_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_235_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_235_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_235_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_235_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_235_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_235_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_235_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_235_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_235_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_235_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_235_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_235_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_235_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_235_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_235_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_235_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_235_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_235_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_235_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_235_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_235_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_235_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_235_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_235_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_235_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_235_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_235_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_235_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_235_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_235_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_235_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_235_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_235_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_235_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_235_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_235_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_236_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_236_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_236_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_236_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_236_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_236_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_236_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_236_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_236_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_236_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_236_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_236_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_236_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_236_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_236_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_236_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_236_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_236_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_236_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_236_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_236_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_236_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_236_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_236_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_236_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_236_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_236_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_236_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_236_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_236_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_236_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_236_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_236_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_236_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_236_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_237_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_237_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_237_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_237_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_237_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_237_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_237_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_237_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_237_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_237_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_237_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_237_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_237_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_237_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_237_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_237_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_237_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_237_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_237_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_237_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_237_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_237_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_237_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_237_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_237_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_237_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_237_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_237_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_237_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_237_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_237_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_237_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_237_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_237_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_237_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_237_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_237_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_237_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_238_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_238_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_238_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_238_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_238_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_238_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_238_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_238_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_238_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_238_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_238_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_238_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_238_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_238_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_238_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_238_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_238_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_238_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_238_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_238_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_238_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_238_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_238_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_238_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_238_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_239_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_239_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_239_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_239_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_239_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_239_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_239_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_239_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_239_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_239_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_239_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_239_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_239_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_239_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_239_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_239_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_239_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_239_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_239_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_239_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_239_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_239_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_239_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_239_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_239_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_239_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_239_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_239_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_239_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_239_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_239_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_239_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_239_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_23_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_240_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_240_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_240_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_240_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_240_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_240_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_240_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_240_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_240_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_240_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_240_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_240_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_240_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_240_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_240_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_240_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_240_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_240_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_240_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_240_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_240_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_240_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_240_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_240_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_240_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_240_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_240_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_240_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_241_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_241_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_241_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_241_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_241_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_241_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_241_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_241_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_241_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_241_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_241_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_241_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_241_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_241_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_241_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_241_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_241_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_241_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_241_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_241_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_241_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_241_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_241_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_242_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_242_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_242_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_242_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_242_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_242_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_242_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_242_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_242_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_242_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_242_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_242_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_242_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_242_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_242_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_242_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_242_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_242_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_242_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_242_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_242_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_242_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_242_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_242_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_242_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_242_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_242_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_242_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_242_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_242_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_242_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_242_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_242_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_242_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_242_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_242_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_243_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_243_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_243_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_243_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_243_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_243_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_243_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_243_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_243_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_243_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_243_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_243_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_243_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_243_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_243_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_243_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_243_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_243_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_243_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_243_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_243_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_243_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_243_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_243_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_243_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_243_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_243_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_243_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_243_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_243_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_243_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_244_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_244_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_244_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_244_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_244_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_244_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_244_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_244_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_244_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_244_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_244_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_244_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_244_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_244_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_244_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_244_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_244_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_244_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_244_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_244_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_244_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_244_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_244_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_244_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_244_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_244_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_244_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_244_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_244_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_244_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_244_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_244_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_244_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_244_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_244_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_244_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_244_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_244_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_244_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_244_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_244_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_245_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_245_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_245_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_245_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_245_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_245_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_245_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_245_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_245_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_245_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_245_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_245_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_245_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_245_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_245_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_245_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_245_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_245_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_245_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_245_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_245_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_245_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_245_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_245_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_245_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_245_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_245_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_245_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_245_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_245_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_245_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_245_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_245_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_245_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_245_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_245_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_245_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_245_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_245_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_246_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_246_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_246_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_246_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_246_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_246_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_246_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_246_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_246_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_246_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_246_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_246_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_246_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_246_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_246_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_246_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_246_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_246_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_246_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_246_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_246_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_246_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_246_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_246_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_246_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_246_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_246_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_246_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_246_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_246_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_246_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_246_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_246_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_246_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_246_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_246_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_246_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_246_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_246_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_246_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_246_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_246_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_247_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_247_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_247_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_247_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_247_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_247_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_247_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_247_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_247_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_247_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_247_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_247_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_247_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_247_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_247_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_247_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_247_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_247_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_247_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_247_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_247_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_247_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_247_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_247_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_247_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_247_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_247_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_247_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_247_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_247_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_247_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_247_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_247_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_247_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_247_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_247_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_247_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_247_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_248_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_248_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_248_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_248_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_248_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_248_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_248_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_248_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_248_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_248_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_248_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_248_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_248_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_248_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_248_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_248_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_248_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_248_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_248_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_248_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_248_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_248_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_248_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_248_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_248_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_248_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_248_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_248_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_248_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_249_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_249_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_249_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_249_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_249_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_249_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_249_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_249_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_249_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_249_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_249_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_249_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_249_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_249_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_249_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_249_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_249_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_249_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_249_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_249_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_249_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_249_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_249_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_249_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_249_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_249_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_249_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_249_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_249_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_249_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_250_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_250_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_250_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_250_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_250_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_250_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_250_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_250_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_250_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_250_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_250_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_250_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_250_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_250_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_250_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_250_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_250_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_250_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_250_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_250_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_250_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_250_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_250_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_250_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_250_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_250_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_250_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_250_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_251_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_251_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_251_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_251_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_251_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_251_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_251_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_251_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_251_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_251_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_251_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_251_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_251_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_251_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_251_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_251_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_251_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_251_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_251_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_251_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_251_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_251_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_251_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_251_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_251_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_251_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_251_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_251_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_251_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_251_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_251_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_251_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_251_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_251_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_251_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_251_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_251_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_252_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_252_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_252_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_252_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_252_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_252_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_252_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_252_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_252_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_252_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_252_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_252_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_252_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_252_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_252_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_252_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_252_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_252_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_252_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_252_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_252_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_252_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_252_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_252_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_252_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_252_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_252_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_252_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_252_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_252_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_252_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_252_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_252_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_252_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_252_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_252_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_252_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_252_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_252_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_252_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_253_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_253_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_253_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_253_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_253_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_253_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_253_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_253_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_253_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_253_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_253_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_253_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_253_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_253_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_253_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_253_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_253_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_253_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_253_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_253_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_253_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_253_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_253_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_253_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_253_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_253_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_253_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_253_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_253_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_253_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_253_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_253_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_253_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_253_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_253_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_253_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_253_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_253_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_253_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_253_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_253_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_253_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_253_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_253_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_254_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_254_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_254_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_254_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_254_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_254_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_254_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_254_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_254_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_254_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_254_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_254_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_254_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_254_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_254_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_254_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_254_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_254_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_254_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_254_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_254_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_254_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_254_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_254_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_254_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_254_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_254_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_254_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_254_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_254_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_254_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_254_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_254_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_254_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_255_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_255_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_255_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_255_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_255_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_255_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_255_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_255_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_255_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_255_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_255_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_255_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_255_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_255_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_255_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_255_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_255_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_255_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_255_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_255_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_255_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_255_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_255_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_255_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_255_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_255_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_255_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_255_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_255_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_255_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_255_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_255_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_256_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_256_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_256_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_256_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_256_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_256_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_256_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_256_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_256_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_256_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_256_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_256_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_256_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_256_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_256_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_256_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_256_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_256_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_256_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_256_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_256_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_256_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_256_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_256_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_256_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_256_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_256_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_256_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_256_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_256_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_257_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_257_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_257_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_257_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_257_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_257_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_257_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_257_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_257_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_257_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_257_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_257_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_257_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_257_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_257_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_257_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_257_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_257_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_257_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_257_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_257_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_257_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_257_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_257_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_258_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_258_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_258_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_258_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_258_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_258_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_258_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_258_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_258_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_258_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_258_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_258_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_258_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_258_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_258_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_258_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_258_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_258_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_258_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_258_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_258_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_258_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_258_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_258_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_258_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_258_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_258_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_258_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_258_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_258_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_258_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_258_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_258_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_258_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_258_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_258_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_258_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_258_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_258_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_258_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_258_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_258_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_259_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_259_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_259_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_259_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_259_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_259_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_259_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_259_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_259_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_259_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_259_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_259_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_259_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_259_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_259_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_259_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_259_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_259_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_259_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_259_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_259_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_259_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_259_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_259_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_259_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_259_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_259_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_259_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_259_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_259_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_259_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_259_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_259_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_259_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_259_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_259_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_259_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_259_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_259_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_259_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_259_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_25_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_25_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_260_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_260_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_260_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_260_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_260_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_260_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_260_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_260_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_260_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_260_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_260_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_260_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_260_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_260_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_260_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_260_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_260_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_260_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_260_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_260_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_260_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_260_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_260_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_260_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_261_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_261_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_261_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_261_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_261_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_261_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_261_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_261_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_261_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_261_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_261_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_261_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_261_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_261_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_261_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_261_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_261_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_261_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_261_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_261_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_261_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_261_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_261_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_261_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_261_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_261_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_261_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_261_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_262_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_262_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_262_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_262_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_262_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_262_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_262_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_262_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_262_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_262_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_262_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_262_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_262_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_262_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_262_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_262_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_262_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_262_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_262_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_262_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_262_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_262_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_262_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_262_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_262_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_262_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_262_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_262_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_262_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_262_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_262_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_262_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_262_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_262_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_262_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_262_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_262_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_262_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_262_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_262_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_262_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_262_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_262_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_262_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_262_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_262_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_262_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_263_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_263_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_263_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_263_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_263_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_263_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_263_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_263_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_263_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_263_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_263_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_263_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_263_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_263_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_263_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_263_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_263_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_263_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_263_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_263_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_263_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_263_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_263_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_263_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_263_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_263_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_263_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_263_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_263_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_263_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_263_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_263_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_263_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_263_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_263_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_264_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_264_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_264_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_264_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_264_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_264_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_264_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_264_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_264_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_264_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_264_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_264_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_264_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_264_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_264_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_264_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_264_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_264_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_264_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_264_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_264_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_264_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_264_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_264_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_264_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_264_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_264_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_264_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_264_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_264_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_264_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_264_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_264_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_265_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_265_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_265_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_265_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_265_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_265_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_265_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_265_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_265_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_265_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_265_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_265_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_265_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_265_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_265_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_265_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_265_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_265_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_265_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_265_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_265_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_265_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_265_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_265_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_265_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_265_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_265_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_265_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_265_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_265_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_265_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_265_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_265_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_265_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_265_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_265_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_265_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_265_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_265_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_265_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_265_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_265_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_266_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_266_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_266_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_266_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_266_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_266_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_266_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_266_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_266_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_266_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_266_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_266_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_266_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_266_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_266_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_266_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_266_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_266_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_266_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_266_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_266_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_266_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_266_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_266_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_266_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_266_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_266_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_266_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_266_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_266_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_266_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_266_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_266_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_266_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_267_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_267_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_267_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_267_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_267_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_267_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_267_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_267_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_267_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_267_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_267_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_267_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_267_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_267_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_267_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_267_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_267_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_267_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_267_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_267_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_267_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_267_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_267_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_267_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_267_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_267_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_267_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_267_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_267_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_267_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_267_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_268_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_268_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_268_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_268_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_268_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_268_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_268_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_268_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_268_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_268_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_268_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_268_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_268_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_268_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_268_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_268_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_268_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_268_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_268_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_268_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_268_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_268_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_268_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_268_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_268_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_268_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_268_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_268_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_268_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_268_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_269_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_269_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_269_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_269_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_269_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_269_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_269_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_269_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_269_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_269_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_269_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_269_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_269_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_269_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_269_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_269_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_269_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_269_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_269_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_269_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_269_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_269_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_269_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_269_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_269_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_269_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_269_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_269_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_269_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_269_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_269_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_269_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_269_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_269_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_269_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_269_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_269_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_269_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_269_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_269_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_269_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_26_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_270_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_270_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_270_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_270_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_270_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_270_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_270_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_270_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_270_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_270_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_270_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_270_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_270_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_270_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_270_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_270_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_270_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_270_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_270_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_270_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_270_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_270_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_270_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_270_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_270_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_270_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_270_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_270_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_270_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_270_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_271_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_271_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_271_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_271_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_271_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_271_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_271_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_271_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_271_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_271_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_271_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_271_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_271_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_271_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_271_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_271_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_271_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_271_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_271_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_271_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_271_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_271_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_271_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_271_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_271_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_271_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_271_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_271_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_271_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_271_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_271_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_271_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_272_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_272_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_272_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_272_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_272_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_272_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_272_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_272_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_272_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_272_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_272_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_272_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_272_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_272_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_272_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_272_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_272_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_272_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_272_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_272_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_272_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_272_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_272_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_272_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_272_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_272_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_272_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_273_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_273_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_273_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_273_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_273_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_273_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_273_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_273_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_273_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_273_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_273_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_273_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_273_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_273_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_273_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_273_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_273_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_273_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_273_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_273_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_273_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_273_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_273_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_273_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_273_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_273_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_273_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_273_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_273_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_273_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_273_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_273_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_273_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_273_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_273_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_273_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_273_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_273_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_273_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_273_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_273_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_273_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_273_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_273_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_273_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_273_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_274_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_274_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_274_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_274_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_274_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_274_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_274_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_274_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_274_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_274_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_274_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_274_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_274_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_274_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_274_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_274_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_274_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_274_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_274_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_274_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_274_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_274_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_274_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_274_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_274_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_274_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_274_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_274_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_274_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_274_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_274_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_274_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_275_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_275_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_275_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_275_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_275_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_275_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_275_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_275_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_275_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_275_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_275_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_275_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_275_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_275_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_275_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_275_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_275_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_275_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_275_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_275_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_275_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_275_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_275_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_275_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_275_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_275_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_275_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_275_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_276_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_276_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_276_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_276_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_276_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_276_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_276_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_276_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_276_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_276_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_276_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_276_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_276_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_276_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_276_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_276_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_276_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_276_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_276_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_276_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_276_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_276_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_276_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_276_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_276_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_276_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_276_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_276_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_276_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_276_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_276_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_276_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_276_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_276_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_276_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_276_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_276_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_276_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_276_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_276_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_276_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_276_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_276_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_277_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_277_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_277_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_277_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_277_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_277_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_277_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_277_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_277_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_277_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_277_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_277_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_277_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_277_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_277_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_277_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_277_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_277_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_277_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_277_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_277_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_277_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_277_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_277_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_277_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_277_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_277_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_277_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_277_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_277_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_277_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_277_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_277_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_277_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_277_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_277_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_277_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_277_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_277_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_277_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_277_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_277_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_277_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_277_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_277_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_277_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_277_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_277_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_277_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_278_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_278_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_278_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_278_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_278_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_278_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_278_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_278_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_278_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_278_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_278_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_278_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_278_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_278_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_278_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_278_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_278_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_278_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_278_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_278_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_278_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_278_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_278_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_278_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_278_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_278_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_278_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_278_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_278_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_279_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_279_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_279_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_279_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_279_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_279_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_279_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_279_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_279_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_279_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_279_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_279_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_279_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_279_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_279_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_279_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_279_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_279_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_279_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_279_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_279_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_279_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_279_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_279_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_279_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_279_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_279_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_279_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_279_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_279_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_279_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_279_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_279_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_279_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_279_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_279_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_279_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_279_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_27_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_280_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_280_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_280_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_280_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_280_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_280_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_280_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_280_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_280_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_280_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_280_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_280_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_280_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_280_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_280_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_280_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_280_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_280_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_280_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_280_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_280_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_280_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_280_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_280_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_280_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_280_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_280_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_280_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_280_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_280_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_280_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_281_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_281_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_281_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_281_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_281_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_281_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_281_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_281_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_281_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_281_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_281_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_281_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_281_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_281_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_281_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_281_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_281_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_281_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_281_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_281_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_281_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_281_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_281_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_281_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_282_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_282_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_282_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_282_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_282_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_282_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_282_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_282_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_282_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_282_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_282_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_282_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_282_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_282_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_282_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_282_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_282_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_282_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_282_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_282_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_282_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_282_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_282_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_282_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_282_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_282_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_282_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_282_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_282_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_282_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_282_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_282_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_282_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_283_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_283_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_283_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_283_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_283_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_283_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_283_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_283_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_283_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_283_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_283_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_283_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_283_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_283_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_283_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_283_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_283_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_283_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_283_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_283_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_283_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_284_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_284_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_284_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_284_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_284_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_284_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_284_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_284_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_284_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_284_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_284_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_284_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_284_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_284_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_284_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_284_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_284_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_284_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_284_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_284_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_284_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_284_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_284_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_284_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_284_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_284_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_284_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_284_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_284_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_284_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_284_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_284_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_284_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_284_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_284_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_284_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_284_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_284_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_284_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_284_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_285_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_285_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_285_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_285_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_285_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_285_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_285_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_285_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_285_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_285_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_285_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_285_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_285_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_285_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_285_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_285_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_285_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_285_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_285_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_285_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_285_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_285_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_285_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_285_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_285_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_285_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_285_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_285_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_285_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_285_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_285_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_285_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_285_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_285_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_285_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_285_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_285_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_286_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_286_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_286_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_286_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_286_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_286_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_286_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_286_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_286_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_286_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_286_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_286_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_286_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_286_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_286_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_286_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_286_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_286_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_286_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_286_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_286_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_286_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_286_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_286_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_286_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_286_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_286_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_286_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_286_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_286_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_286_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_286_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_286_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_287_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_287_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_287_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_287_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_287_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_287_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_287_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_287_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_287_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_287_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_287_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_287_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_287_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_287_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_287_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_287_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_287_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_287_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_287_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_287_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_287_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_287_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_287_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_287_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_287_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_287_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_287_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_287_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_287_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_287_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_287_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_287_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_287_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_287_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_287_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_287_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_287_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_287_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_287_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_288_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_288_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_288_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_288_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_288_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_288_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_288_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_288_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_288_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_288_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_288_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_288_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_288_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_288_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_288_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_288_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_288_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_288_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_288_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_288_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_288_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_288_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_288_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_288_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_289_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_289_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_289_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_289_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_289_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_289_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_289_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_289_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_289_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_289_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_289_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_289_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_289_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_289_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_289_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_289_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_289_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_289_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_289_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_289_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_289_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_289_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_289_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_289_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_289_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_289_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_289_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_289_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_290_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_290_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_290_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_290_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_290_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_290_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_290_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_290_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_290_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_290_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_290_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_290_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_290_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_290_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_290_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_290_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_290_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_290_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_290_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_290_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_290_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_290_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_290_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_290_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_290_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_290_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_290_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_291_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_291_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_291_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_291_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_291_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_291_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_291_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_291_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_291_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_291_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_291_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_291_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_291_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_291_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_291_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_291_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_291_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_291_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_291_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_291_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_291_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_291_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_291_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_291_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_291_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_291_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_291_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_291_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_291_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_291_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_292_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_292_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_292_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_292_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_292_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_292_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_292_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_292_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_292_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_292_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_292_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_292_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_292_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_292_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_292_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_292_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_292_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_292_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_292_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_292_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_292_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_292_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_293_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_293_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_293_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_293_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_293_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_293_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_293_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_293_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_293_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_293_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_293_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_293_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_293_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_293_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_293_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_293_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_293_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_293_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_293_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_293_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_294_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_294_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_294_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_294_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_294_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_294_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_294_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_294_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_294_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_294_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_294_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_294_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_294_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_294_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_294_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_294_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_294_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_294_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_294_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_294_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_294_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_294_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_294_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_294_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_294_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_294_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_294_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_294_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_294_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_294_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_294_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_294_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_294_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_294_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_294_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_294_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_294_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_294_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_294_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_294_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_295_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_295_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_295_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_295_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_295_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_295_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_295_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_295_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_295_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_295_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_295_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_295_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_295_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_295_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_295_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_295_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_295_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_295_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_295_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_295_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_295_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_295_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_295_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_295_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_295_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_295_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_295_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_295_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_295_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_295_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_295_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_295_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_295_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_295_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_295_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_295_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_295_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_295_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_295_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_295_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_295_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_296_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_296_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_296_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_296_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_296_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_296_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_296_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_296_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_296_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_296_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_296_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_296_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_296_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_296_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_296_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_296_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_296_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_296_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_296_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_296_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_296_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_296_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_296_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_296_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_296_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_296_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_296_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_296_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_296_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_296_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_296_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_296_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_296_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_297_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_297_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_297_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_297_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_297_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_297_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_297_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_297_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_297_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_297_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_297_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_297_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_297_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_297_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_297_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_297_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_297_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_297_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_297_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_297_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_297_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_297_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_297_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_297_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_297_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_297_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_297_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_297_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_297_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_297_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_297_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_297_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_297_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_297_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_297_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_297_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_297_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_298_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_298_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_298_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_298_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_298_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_298_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_298_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_298_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_298_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_298_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_298_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_298_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_298_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_298_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_298_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_298_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_298_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_298_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_298_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_298_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_298_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_298_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_298_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_298_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_298_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_298_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_298_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_298_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_298_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_298_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_298_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_298_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_298_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_298_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_298_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_298_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_298_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_298_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_299_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_299_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_299_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_299_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_299_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_299_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_299_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_299_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_299_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_299_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_299_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_299_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_299_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_299_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_299_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_299_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_299_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_299_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_299_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_299_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_299_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_299_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_299_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_299_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_299_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_299_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_299_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_299_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_299_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_299_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_299_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_299_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_299_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_299_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_299_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_299_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_299_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_299_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_299_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_299_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_299_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_29_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_300_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_300_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_300_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_300_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_300_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_300_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_300_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_300_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_300_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_300_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_300_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_300_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_300_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_300_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_300_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_300_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_300_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_300_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_300_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_300_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_300_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_300_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_300_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_300_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_300_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_300_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_300_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_300_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_300_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_300_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_300_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_300_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_300_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_300_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_300_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_300_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_300_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_300_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_301_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_301_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_301_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_301_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_301_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_301_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_301_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_301_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_301_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_301_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_301_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_301_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_301_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_301_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_301_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_301_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_301_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_301_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_301_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_301_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_301_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_301_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_301_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_301_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_301_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_301_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_301_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_301_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_302_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_302_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_302_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_302_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_302_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_302_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_302_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_302_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_302_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_302_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_302_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_302_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_302_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_302_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_302_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_302_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_302_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_302_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_302_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_302_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_302_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_302_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_302_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_302_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_302_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_302_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_303_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_303_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_303_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_303_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_303_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_303_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_303_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_303_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_303_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_303_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_303_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_303_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_303_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_303_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_303_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_303_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_303_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_303_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_303_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_303_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_303_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_303_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_303_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_303_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_303_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_303_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_303_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_303_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_304_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_304_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_304_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_304_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_304_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_304_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_304_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_304_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_304_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_304_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_304_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_304_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_304_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_304_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_304_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_304_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_304_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_304_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_304_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_304_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_304_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_304_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_304_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_304_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_304_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_304_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_304_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_304_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_304_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_304_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_304_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_304_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_305_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_305_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_305_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_305_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_305_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_305_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_305_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_305_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_305_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_305_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_305_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_305_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_305_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_305_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_305_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_305_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_305_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_305_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_305_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_305_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_305_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_305_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_305_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_305_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_305_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_305_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_305_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_305_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_305_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_305_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_305_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_305_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_306_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_306_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_306_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_306_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_306_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_306_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_306_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_306_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_306_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_306_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_306_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_306_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_306_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_306_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_306_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_306_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_306_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_306_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_306_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_306_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_306_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_306_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_306_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_306_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_306_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_306_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_306_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_306_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_306_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_306_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_306_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_306_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_306_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_307_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_307_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_307_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_307_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_307_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_307_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_307_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_307_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_307_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_307_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_307_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_307_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_307_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_307_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_307_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_307_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_307_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_307_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_307_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_307_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_307_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_307_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_307_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_307_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_307_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_307_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_307_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_307_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_307_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_307_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_307_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_307_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_307_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_307_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_307_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_307_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_307_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_307_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_307_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_307_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_307_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_308_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_308_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_308_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_308_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_308_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_308_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_308_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_308_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_308_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_308_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_308_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_308_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_308_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_308_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_308_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_308_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_308_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_308_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_308_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_308_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_308_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_308_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_308_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_308_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_308_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_308_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_308_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_308_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_308_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_308_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_308_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_308_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_308_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_308_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_308_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_308_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_308_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_308_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_308_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_308_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_308_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_308_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_308_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_308_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_308_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_309_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_309_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_309_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_309_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_309_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_309_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_309_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_309_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_309_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_309_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_309_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_309_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_309_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_309_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_309_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_309_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_309_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_309_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_309_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_309_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_309_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_309_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_309_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_309_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_309_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_309_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_309_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_309_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_309_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_309_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_309_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_309_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_309_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_309_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_309_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_309_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_309_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_309_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_309_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_309_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_309_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_309_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_309_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_310_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_310_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_310_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_310_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_310_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_310_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_310_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_310_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_310_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_310_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_310_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_310_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_310_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_310_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_310_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_310_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_310_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_310_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_310_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_310_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_310_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_310_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_310_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_310_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_310_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_310_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_310_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_310_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_310_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_310_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_311_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_311_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_311_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_311_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_311_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_311_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_311_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_311_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_311_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_311_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_311_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_311_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_311_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_311_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_311_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_311_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_311_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_311_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_311_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_311_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_311_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_311_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_311_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_311_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_311_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_311_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_311_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_311_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_311_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_311_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_312_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_312_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_312_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_312_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_312_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_312_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_312_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_312_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_312_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_312_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_312_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_312_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_312_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_312_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_312_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_312_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_312_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_312_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_312_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_312_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_312_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_312_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_312_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_312_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_312_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_312_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_312_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_312_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_312_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_313_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_313_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_313_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_313_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_313_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_313_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_313_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_313_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_313_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_313_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_313_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_313_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_313_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_313_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_313_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_313_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_313_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_313_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_313_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_313_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_313_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_313_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_313_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_313_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_313_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_313_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_313_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_313_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_313_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_313_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_313_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_314_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_314_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_314_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_314_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_314_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_314_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_314_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_314_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_314_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_314_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_314_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_314_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_314_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_314_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_314_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_314_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_314_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_314_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_314_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_314_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_314_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_314_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_314_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_314_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_314_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_314_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_314_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_314_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_314_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_314_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_314_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_315_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_315_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_315_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_315_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_315_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_315_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_315_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_315_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_315_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_315_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_315_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_315_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_315_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_315_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_315_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_315_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_315_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_315_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_315_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_315_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_315_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_315_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_315_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_315_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_315_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_315_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_315_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_315_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_315_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_315_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_315_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_315_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_315_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_316_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_316_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_316_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_316_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_316_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_316_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_316_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_316_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_316_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_316_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_316_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_316_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_316_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_316_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_316_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_316_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_316_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_316_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_316_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_316_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_316_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_316_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_316_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_316_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_316_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_317_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_317_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_317_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_317_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_317_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_317_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_317_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_317_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_317_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_317_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_317_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_317_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_317_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_317_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_317_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_317_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_317_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_317_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_317_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_317_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_317_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_317_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_317_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_317_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_317_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_317_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_317_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_317_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_317_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_317_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_317_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_317_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_317_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_317_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_317_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_318_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_318_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_318_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_318_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_318_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_318_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_318_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_318_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_318_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_318_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_318_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_318_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_318_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_318_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_318_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_318_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_318_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_318_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_318_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_318_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_318_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_318_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_318_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_318_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_318_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_318_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_318_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_318_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_318_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_318_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_319_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_319_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_319_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_319_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_319_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_319_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_319_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_319_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_319_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_319_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_319_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_319_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_319_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_319_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_319_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_319_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_319_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_319_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_319_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_319_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_319_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_319_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_319_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_319_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_319_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_319_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_31_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_320_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_320_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_320_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_320_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_320_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_320_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_320_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_320_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_320_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_320_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_320_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_320_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_320_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_320_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_320_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_320_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_320_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_320_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_320_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_320_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_320_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_320_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_320_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_320_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_320_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_320_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_320_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_320_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_320_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_320_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_320_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_320_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_320_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_320_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_320_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_320_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_320_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_320_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_320_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_320_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_321_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_321_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_321_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_321_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_321_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_321_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_321_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_321_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_321_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_321_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_321_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_321_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_321_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_321_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_321_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_321_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_321_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_321_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_321_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_321_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_321_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_321_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_321_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_321_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_321_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_321_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_321_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_321_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_321_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_321_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_321_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_322_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_322_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_322_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_322_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_322_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_322_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_322_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_322_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_322_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_322_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_322_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_322_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_322_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_322_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_322_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_322_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_322_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_322_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_322_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_322_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_322_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_322_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_322_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_322_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_322_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_322_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_322_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_322_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_322_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_322_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_323_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_323_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_323_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_323_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_323_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_323_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_323_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_323_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_323_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_323_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_323_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_323_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_323_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_323_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_323_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_323_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_323_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_323_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_323_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_323_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_323_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_323_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_323_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_323_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_323_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_323_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_323_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_323_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_324_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_324_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_324_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_324_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_324_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_324_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_324_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_324_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_324_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_324_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_324_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_324_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_324_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_324_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_324_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_324_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_324_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_324_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_324_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_324_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_324_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_324_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_324_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_324_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_324_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_325_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_325_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_325_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_325_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_325_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_325_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_325_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_325_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_325_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_325_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_325_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_325_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_325_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_325_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_325_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_325_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_325_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_325_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_325_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_325_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_325_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_325_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_325_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_325_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_325_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_325_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_325_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_325_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_325_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_325_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_325_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_325_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_325_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_325_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_325_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_325_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_325_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_325_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_326_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_326_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_326_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_326_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_326_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_326_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_326_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_326_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_326_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_326_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_326_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_326_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_326_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_326_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_326_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_326_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_326_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_326_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_326_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_326_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_326_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_326_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_326_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_326_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_326_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_326_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_326_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_326_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_326_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_326_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_326_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_327_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_327_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_327_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_327_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_327_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_327_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_327_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_327_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_327_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_327_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_327_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_327_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_327_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_327_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_327_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_327_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_327_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_327_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_327_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_327_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_327_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_327_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_327_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_327_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_327_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_327_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_327_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_327_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_327_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_327_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_327_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_327_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_327_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_327_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_327_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_327_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_327_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_327_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_327_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_327_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_327_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_327_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_327_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_328_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_328_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_328_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_328_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_328_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_328_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_328_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_328_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_328_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_328_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_328_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_328_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_328_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_328_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_328_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_328_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_328_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_328_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_328_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_328_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_328_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_328_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_328_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_328_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_328_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_328_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_328_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_328_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_328_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_328_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_328_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_329_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_329_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_329_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_329_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_329_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_329_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_329_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_329_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_329_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_329_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_329_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_329_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_329_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_329_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_329_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_329_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_329_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_329_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_329_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_329_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_329_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_329_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_329_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_329_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_329_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_329_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_329_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_329_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_329_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_329_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_329_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_329_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_329_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_329_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_329_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_329_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_329_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_329_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_329_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_329_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_329_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_329_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_329_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_329_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_329_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_329_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_329_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_330_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_330_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_330_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_330_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_330_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_330_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_330_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_330_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_330_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_330_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_330_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_330_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_330_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_330_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_330_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_330_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_330_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_330_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_330_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_330_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_330_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_330_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_330_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_330_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_330_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_330_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_330_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_330_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_330_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_330_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_330_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_330_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_330_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_330_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_330_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_330_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_331_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_331_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_331_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_331_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_331_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_331_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_331_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_331_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_331_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_331_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_331_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_331_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_331_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_331_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_331_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_331_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_331_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_331_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_331_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_331_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_331_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_331_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_331_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_331_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_331_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_331_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_331_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_331_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_331_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_331_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_331_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_331_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_331_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_331_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_331_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_331_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_331_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_332_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_332_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_332_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_332_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_332_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_332_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_332_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_332_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_332_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_332_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_332_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_332_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_332_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_332_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_332_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_332_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_332_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_332_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_332_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_332_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_332_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_332_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_332_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_332_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_332_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_332_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_332_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_332_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_332_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_332_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_333_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_333_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_333_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_333_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_333_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_333_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_333_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_333_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_333_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_333_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_333_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_333_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_333_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_333_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_333_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_333_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_333_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_333_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_333_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_333_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_333_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_333_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_333_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_333_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_333_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_333_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_333_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_333_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_333_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_333_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_333_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_333_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_333_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_333_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_333_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_333_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_333_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_334_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_334_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_334_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_334_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_334_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_334_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_334_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_334_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_334_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_334_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_334_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_334_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_334_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_334_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_334_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_334_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_334_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_334_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_334_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_334_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_334_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_334_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_334_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_334_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_334_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_334_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_334_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_334_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_334_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_335_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_335_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_335_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_335_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_335_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_335_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_335_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_335_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_335_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_335_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_335_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_335_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_335_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_335_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_335_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_335_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_335_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_335_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_335_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_335_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_335_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_335_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_335_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_335_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_335_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_335_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_335_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_335_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_335_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_335_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_335_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_335_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_335_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_335_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_335_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_335_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_335_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_336_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_336_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_336_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_336_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_336_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_336_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_336_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_336_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_336_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_336_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_336_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_336_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_336_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_336_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_336_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_336_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_336_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_336_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_336_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_336_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_336_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_336_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_336_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_336_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_336_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_336_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_336_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_336_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_336_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_336_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_336_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_336_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_336_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_336_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_337_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_337_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_337_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_337_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_337_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_337_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_337_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_337_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_337_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_337_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_337_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_337_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_337_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_337_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_337_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_337_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_337_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_337_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_337_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_337_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_337_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_337_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_337_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_337_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_337_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_337_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_338_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_338_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_338_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_338_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_338_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_338_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_338_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_338_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_338_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_338_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_338_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_338_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_338_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_338_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_338_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_338_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_338_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_338_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_338_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_338_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_338_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_338_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_338_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_338_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_338_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_338_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_338_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_339_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_339_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_339_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_339_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_339_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_339_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_339_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_339_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_339_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_339_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_339_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_339_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_339_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_339_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_339_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_339_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_339_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_339_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_339_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_339_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_339_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_339_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_339_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_339_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_339_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_339_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_339_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_339_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_339_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_339_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_33_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_340_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_340_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_340_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_340_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_340_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_340_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_340_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_340_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_340_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_340_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_340_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_340_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_340_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_340_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_340_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_340_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_340_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_340_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_340_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_340_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_340_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_340_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_340_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_340_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_340_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_340_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_341_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_341_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_341_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_341_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_341_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_341_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_341_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_341_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_341_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_341_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_341_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_341_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_341_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_341_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_341_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_341_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_341_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_341_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_341_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_341_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_341_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_341_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_341_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_341_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_341_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_341_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_341_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_341_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_341_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_341_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_341_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_341_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_341_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_341_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_341_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_341_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_342_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_342_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_342_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_342_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_342_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_342_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_342_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_342_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_342_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_342_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_342_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_342_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_342_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_342_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_342_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_342_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_342_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_342_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_342_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_342_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_342_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_342_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_342_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_342_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_342_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_342_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_342_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_342_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_342_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_342_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_342_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_342_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_342_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_342_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_342_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_342_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_342_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_342_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_342_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_342_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_343_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_343_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_343_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_343_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_343_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_343_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_343_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_343_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_343_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_343_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_343_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_343_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_343_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_343_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_343_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_343_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_343_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_343_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_343_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_343_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_343_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_343_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_343_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_343_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_343_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_343_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_343_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_343_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_344_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_344_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_344_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_344_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_344_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_344_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_344_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_344_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_344_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_344_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_344_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_344_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_344_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_344_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_344_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_344_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_344_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_344_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_344_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_344_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_344_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_344_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_344_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_344_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_344_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_344_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_344_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_344_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_344_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_344_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_344_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_344_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_344_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_344_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_344_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_344_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_344_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_344_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_345_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_345_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_345_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_345_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_345_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_345_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_345_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_345_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_345_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_345_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_345_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_345_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_345_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_345_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_345_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_345_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_345_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_345_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_345_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_345_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_345_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_345_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_345_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_345_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_345_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_345_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_345_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_345_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_345_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_345_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_345_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_345_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_345_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_345_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_345_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_345_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_345_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_345_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_345_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_345_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_345_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_345_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_346_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_346_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_346_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_346_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_346_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_346_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_346_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_346_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_346_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_346_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_346_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_346_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_346_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_346_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_346_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_346_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_346_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_346_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_346_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_346_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_346_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_346_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_346_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_346_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_346_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_346_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_346_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_346_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_346_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_346_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_346_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_347_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_347_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_347_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_347_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_347_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_347_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_347_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_347_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_347_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_347_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_347_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_347_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_347_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_347_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_347_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_347_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_347_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_347_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_347_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_347_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_347_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_347_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_347_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_347_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_347_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_347_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_347_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_347_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_347_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_347_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_347_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_348_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_348_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_348_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_348_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_348_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_348_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_348_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_348_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_348_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_348_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_348_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_348_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_348_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_348_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_348_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_348_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_348_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_348_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_348_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_348_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_348_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_348_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_348_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_348_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_348_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_348_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_348_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_349_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_349_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_349_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_349_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_349_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_349_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_349_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_349_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_349_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_349_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_349_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_349_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_349_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_349_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_349_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_349_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_349_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_349_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_349_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_349_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_349_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_349_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_349_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_349_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_349_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_349_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_349_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_349_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_349_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_349_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_349_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_349_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_349_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_349_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_350_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_350_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_350_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_350_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_350_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_350_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_350_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_350_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_350_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_350_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_350_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_350_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_350_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_350_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_350_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_350_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_350_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_350_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_350_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_350_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_350_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_350_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_350_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_350_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_350_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_350_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_350_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_350_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_351_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_351_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_351_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_351_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_351_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_351_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_351_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_351_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_351_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_351_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_351_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_351_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_351_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_351_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_351_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_351_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_351_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_351_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_351_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_351_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_351_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_351_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_351_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_351_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_351_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_351_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_351_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_351_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_351_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_351_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_351_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_351_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_351_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_351_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_351_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_351_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_351_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_351_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_352_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_352_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_352_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_352_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_352_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_352_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_352_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_352_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_352_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_352_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_352_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_352_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_352_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_352_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_352_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_352_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_352_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_352_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_352_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_352_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_352_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_352_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_352_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_352_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_352_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_353_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_353_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_353_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_353_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_353_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_353_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_353_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_353_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_353_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_353_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_353_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_353_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_353_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_353_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_353_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_353_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_353_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_353_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_353_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_353_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_353_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_353_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_353_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_353_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_353_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_353_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_353_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_353_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_353_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_353_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_353_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_353_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_353_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_353_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_353_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_354_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_354_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_354_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_354_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_354_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_354_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_354_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_354_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_354_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_354_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_354_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_354_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_354_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_354_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_354_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_354_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_354_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_354_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_354_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_354_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_354_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_354_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_354_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_354_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_354_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_354_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_354_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_354_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_354_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_354_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_354_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_354_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_354_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_355_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_355_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_355_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_355_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_355_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_355_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_355_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_355_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_355_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_355_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_355_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_355_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_355_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_355_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_355_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_355_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_355_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_355_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_355_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_355_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_355_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_355_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_355_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_355_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_355_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_355_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_355_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_355_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_355_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_355_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_355_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_355_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_355_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_355_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_355_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_355_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_355_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_355_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_356_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_356_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_356_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_356_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_356_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_356_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_356_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_356_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_356_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_356_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_356_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_356_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_356_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_356_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_356_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_356_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_356_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_356_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_356_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_356_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_356_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_356_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_356_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_356_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_357_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_357_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_357_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_357_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_357_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_357_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_357_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_357_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_357_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_357_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_357_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_357_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_357_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_357_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_357_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_357_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_357_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_357_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_357_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_357_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_357_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_357_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_357_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_357_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_357_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_358_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_358_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_358_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_358_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_358_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_358_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_358_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_358_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_358_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_358_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_358_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_358_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_358_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_358_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_358_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_358_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_358_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_358_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_358_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_358_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_358_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_358_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_358_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_358_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_358_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_358_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_358_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_358_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_358_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_358_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_358_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_358_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_359_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_359_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_359_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_359_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_359_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_359_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_359_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_359_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_359_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_359_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_359_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_359_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_359_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_359_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_359_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_359_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_359_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_359_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_359_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_359_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_359_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_359_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_359_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_359_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_359_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_359_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_359_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_359_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_359_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_359_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_359_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_359_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_359_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_359_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_359_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_359_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_359_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_359_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_35_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_360_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_360_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_360_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_360_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_360_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_360_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_360_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_360_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_360_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_360_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_360_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_360_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_360_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_360_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_360_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_360_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_360_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_360_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_360_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_360_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_360_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_360_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_360_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_360_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_360_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_360_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_360_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_360_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_360_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_360_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_360_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_360_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_360_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_360_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_360_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_360_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_360_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_360_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_360_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_361_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_361_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_361_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_361_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_361_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_361_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_361_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_361_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_361_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_361_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_361_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_361_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_361_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_361_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_361_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_361_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_361_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_361_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_361_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_361_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_361_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_361_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_361_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_361_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_361_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_361_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_361_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_361_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_361_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_361_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_361_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_361_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_361_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_362_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_362_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_362_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_362_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_362_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_362_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_362_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_362_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_362_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_362_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_362_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_362_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_362_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_362_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_362_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_362_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_362_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_362_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_362_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_362_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_362_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_362_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_362_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_362_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_362_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_362_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_362_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_362_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_362_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_362_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_362_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_362_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_362_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_362_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_362_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_362_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_362_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_362_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_362_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_363_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_363_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_363_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_363_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_363_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_363_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_363_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_363_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_363_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_363_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_363_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_363_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_363_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_363_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_363_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_363_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_363_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_363_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_363_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_363_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_363_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_363_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_363_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_363_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_363_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_363_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_363_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_363_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_363_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_363_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_363_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_363_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_363_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_363_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_363_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_363_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_363_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_364_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_364_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_364_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_364_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_364_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_364_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_364_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_364_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_364_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_364_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_364_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_364_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_364_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_364_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_364_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_364_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_364_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_364_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_364_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_364_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_364_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_364_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_364_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_364_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_364_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_364_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_364_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_364_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_364_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_364_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_364_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_364_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_364_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_364_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_364_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_364_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_364_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_364_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_364_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_364_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_365_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_365_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_365_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_365_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_365_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_365_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_365_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_365_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_365_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_365_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_365_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_365_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_365_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_365_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_365_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_365_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_365_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_365_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_365_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_365_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_365_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_365_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_365_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_365_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_365_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_365_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_365_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_365_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_365_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_365_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_366_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_366_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_366_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_366_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_366_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_366_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_366_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_366_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_366_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_366_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_366_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_366_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_366_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_366_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_366_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_366_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_366_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_366_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_366_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_366_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_366_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_366_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_366_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_366_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_366_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_366_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_366_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_366_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_366_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_366_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_366_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_366_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_366_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_366_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_366_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_366_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_366_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_367_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_367_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_367_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_367_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_367_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_367_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_367_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_367_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_367_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_367_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_367_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_367_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_367_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_367_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_367_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_367_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_367_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_367_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_367_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_367_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_367_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_367_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_367_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_367_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_367_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_367_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_367_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_367_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_367_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_367_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_367_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_367_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_367_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_367_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_367_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_368_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_368_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_368_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_368_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_368_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_368_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_368_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_368_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_368_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_368_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_368_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_368_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_368_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_368_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_368_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_368_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_368_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_368_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_368_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_368_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_368_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_368_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_368_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_368_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_368_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_368_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_368_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_369_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_369_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_369_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_369_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_369_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_369_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_369_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_369_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_369_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_369_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_369_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_369_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_369_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_369_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_369_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_369_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_369_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_369_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_369_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_369_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_369_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_369_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_369_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_369_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_369_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_369_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_369_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_369_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_369_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_369_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_370_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_370_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_370_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_370_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_370_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_370_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_370_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_370_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_370_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_370_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_370_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_370_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_370_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_370_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_370_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_370_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_370_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_370_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_370_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_370_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_370_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_370_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_370_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_370_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_370_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_370_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_370_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_370_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_370_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_370_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_370_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_370_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_370_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_371_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_371_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_371_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_371_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_371_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_371_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_371_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_371_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_371_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_371_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_371_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_371_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_371_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_371_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_371_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_371_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_371_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_371_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_371_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_371_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_371_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_371_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_371_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_371_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_371_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_371_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_371_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_371_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_371_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_371_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_371_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_371_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_371_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_371_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_371_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_371_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_371_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_372_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_372_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_372_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_372_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_372_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_372_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_372_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_372_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_372_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_372_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_372_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_372_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_372_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_372_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_372_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_372_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_372_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_372_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_372_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_372_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_372_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_372_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_372_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_372_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_372_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_372_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_372_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_372_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_372_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_372_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_372_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_372_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_372_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_372_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_372_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_372_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_372_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_373_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_373_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_373_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_373_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_373_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_373_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_373_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_373_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_373_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_373_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_373_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_373_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_373_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_373_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_373_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_373_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_373_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_373_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_373_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_373_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_373_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_373_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_373_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_373_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_373_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_373_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_373_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_373_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_374_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_374_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_374_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_374_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_374_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_374_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_374_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_374_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_374_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_374_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_374_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_374_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_374_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_374_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_374_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_374_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_374_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_374_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_374_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_374_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_374_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_374_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_374_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_374_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_374_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_374_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_374_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_375_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_375_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_375_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_375_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_375_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_375_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_375_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_375_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_375_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_375_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_375_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_375_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_375_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_375_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_375_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_375_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_375_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_375_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_375_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_375_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_375_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_375_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_375_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_375_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_375_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_375_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_375_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_375_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_376_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_376_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_376_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_376_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_376_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_376_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_376_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_376_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_376_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_376_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_376_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_376_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_376_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_376_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_376_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_376_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_376_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_376_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_376_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_376_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_376_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_376_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_376_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_376_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_376_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_376_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_376_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_376_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_376_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_376_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_376_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_376_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_376_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_376_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_377_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_377_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_377_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_377_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_377_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_377_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_377_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_377_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_377_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_377_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_377_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_377_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_377_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_377_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_377_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_377_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_377_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_377_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_377_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_377_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_377_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_377_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_377_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_377_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_377_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_377_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_377_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_377_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_377_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_377_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_377_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_377_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_377_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_377_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_378_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_378_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_378_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_378_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_378_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_378_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_378_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_378_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_378_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_378_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_378_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_378_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_378_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_378_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_378_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_378_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_378_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_378_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_378_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_378_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_378_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_378_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_378_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_378_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_378_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_378_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_378_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_378_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_378_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_378_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_378_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_378_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_378_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_378_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_378_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_378_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_378_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_378_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_379_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_379_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_379_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_379_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_379_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_379_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_379_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_379_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_379_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_379_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_379_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_379_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_379_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_379_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_379_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_379_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_379_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_379_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_379_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_379_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_379_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_379_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_379_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_379_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_379_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_379_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_379_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_379_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_379_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_379_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_379_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_379_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_379_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_379_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_379_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_379_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_379_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_379_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_380_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_380_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_380_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_380_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_380_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_380_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_380_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_380_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_380_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_380_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_380_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_380_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_380_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_380_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_380_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_380_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_380_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_380_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_380_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_380_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_380_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_380_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_380_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_380_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_380_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_380_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_380_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_380_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_380_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_380_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_380_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_381_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_381_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_381_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_381_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_381_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_381_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_381_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_381_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_381_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_381_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_381_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_381_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_381_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_381_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_381_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_381_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_381_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_381_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_381_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_381_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_381_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_381_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_381_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_381_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_381_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_381_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_381_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_381_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_381_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_381_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_382_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_382_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_382_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_382_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_382_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_382_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_382_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_382_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_382_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_382_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_382_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_382_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_382_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_382_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_382_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_382_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_382_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_382_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_382_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_382_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_382_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_382_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_382_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_382_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_382_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_382_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_382_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_382_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_382_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_382_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_383_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_383_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_383_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_383_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_383_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_383_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_383_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_383_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_383_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_383_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_383_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_383_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_383_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_383_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_383_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_383_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_383_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_383_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_383_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_383_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_383_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_383_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_383_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_383_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_383_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_383_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_383_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_383_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_383_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_383_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_383_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_383_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_384_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_384_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_384_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_384_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_384_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_384_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_384_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_384_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_384_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_384_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_384_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_384_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_384_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_384_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_384_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_384_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_384_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_384_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_384_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_384_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_384_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_384_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_384_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_384_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_384_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_384_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_384_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_384_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_384_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_384_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_384_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_384_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_384_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_384_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_384_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_384_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_384_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_384_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_384_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_384_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_384_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_384_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_384_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_385_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_385_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_385_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_385_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_385_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_385_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_385_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_385_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_385_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_385_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_385_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_385_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_385_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_385_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_385_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_385_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_385_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_385_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_385_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_385_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_385_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_385_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_385_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_385_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_385_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_385_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_385_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_385_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_385_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_385_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_386_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_386_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_386_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_386_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_386_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_386_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_386_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_386_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_386_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_386_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_386_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_386_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_386_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_386_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_386_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_386_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_386_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_386_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_386_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_386_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_386_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_386_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_386_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_386_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_386_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_386_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_386_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_386_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_386_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_386_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_386_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_386_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_386_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_386_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_386_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_386_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_386_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_386_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_386_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_386_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_386_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_386_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_386_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_386_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_386_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_386_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_386_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_387_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_387_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_387_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_387_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_387_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_387_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_387_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_387_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_387_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_387_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_387_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_387_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_387_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_387_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_387_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_387_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_387_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_387_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_387_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_387_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_387_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_387_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_387_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_387_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_387_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_387_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_387_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_387_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_387_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_387_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_388_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_388_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_388_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_388_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_388_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_388_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_388_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_388_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_388_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_388_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_388_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_388_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_388_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_388_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_388_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_388_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_388_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_388_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_388_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_388_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_388_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_388_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_388_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_388_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_389_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_389_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_389_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_389_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_389_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_389_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_389_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_389_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_389_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_389_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_389_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_389_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_389_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_389_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_389_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_389_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_389_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_389_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_389_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_389_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_389_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_389_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_389_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_389_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_389_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_389_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_389_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_389_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_390_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_390_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_390_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_390_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_390_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_390_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_390_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_390_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_390_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_390_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_390_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_390_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_390_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_390_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_390_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_390_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_390_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_390_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_390_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_390_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_390_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_390_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_390_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_390_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_390_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_390_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_390_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_390_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_391_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_391_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_391_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_391_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_391_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_391_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_391_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_391_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_391_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_391_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_391_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_391_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_391_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_391_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_391_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_391_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_391_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_391_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_391_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_391_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_391_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_391_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_391_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_391_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_391_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_391_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_391_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_391_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_391_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_391_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_391_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_392_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_392_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_392_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_392_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_392_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_392_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_392_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_392_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_392_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_392_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_392_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_392_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_392_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_392_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_392_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_392_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_392_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_392_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_392_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_392_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_392_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_392_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_392_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_392_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_392_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_392_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_392_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_392_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_392_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_392_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_392_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_392_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_392_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_392_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_392_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_392_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_392_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_392_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_393_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_393_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_393_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_393_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_393_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_393_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_393_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_393_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_393_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_393_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_393_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_393_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_393_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_393_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_393_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_393_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_393_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_393_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_393_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_393_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_393_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_393_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_393_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_393_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_393_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_393_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_393_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_393_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_393_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_393_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_393_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_393_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_393_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_393_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_393_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_394_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_394_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_394_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_394_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_394_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_394_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_394_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_394_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_394_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_394_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_394_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_394_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_394_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_394_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_394_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_394_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_394_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_394_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_394_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_394_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_394_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_394_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_394_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_394_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_394_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_394_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_394_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_394_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_394_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_394_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_394_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_394_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_394_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_394_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_394_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_394_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_394_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_394_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_394_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_395_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_395_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_395_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_395_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_395_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_395_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_395_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_395_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_395_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_395_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_395_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_395_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_395_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_395_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_395_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_395_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_395_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_395_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_395_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_395_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_395_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_395_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_395_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_395_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_395_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_395_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_395_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_395_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_395_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_395_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_395_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_395_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_395_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_395_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_395_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_395_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_395_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_395_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_395_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_395_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_395_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_396_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_396_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_396_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_396_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_396_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_396_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_396_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_396_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_396_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_396_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_396_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_396_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_396_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_396_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_396_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_396_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_396_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_396_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_396_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_396_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_396_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_396_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_396_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_396_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_396_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_396_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_396_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_396_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_396_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_397_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_397_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_397_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_397_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_397_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_397_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_397_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_397_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_397_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_397_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_397_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_397_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_397_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_397_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_397_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_397_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_397_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_397_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_397_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_397_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_397_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_397_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_397_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_397_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_397_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_397_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_397_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_397_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_397_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_397_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_397_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_397_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_397_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_398_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_398_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_398_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_398_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_398_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_398_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_398_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_398_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_398_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_398_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_398_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_398_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_398_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_398_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_398_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_398_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_398_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_398_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_398_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_398_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_398_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_398_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_398_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_398_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_398_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_398_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_398_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_398_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_398_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_398_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_398_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_398_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_398_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_398_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_398_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_398_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_399_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_399_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_399_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_399_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_399_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_399_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_399_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_399_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_399_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_399_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_399_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_399_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_399_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_399_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_399_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_399_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_399_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_399_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_399_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_399_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_399_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_399_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_399_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_399_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_399_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_399_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_399_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_39_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_3_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_400_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_400_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_400_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_400_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_400_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_400_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_400_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_400_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_400_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_400_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_400_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_400_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_400_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_400_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_400_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_400_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_400_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_400_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_400_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_400_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_401_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_401_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_401_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_401_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_401_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_401_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_401_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_401_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_401_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_401_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_401_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_401_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_401_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_401_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_401_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_401_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_401_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_401_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_401_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_401_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_401_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_401_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_401_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_401_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_401_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_401_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_401_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_401_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_401_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_401_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_401_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_401_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_401_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_401_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_401_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_401_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_401_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_401_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_401_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_402_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_402_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_402_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_402_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_402_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_402_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_402_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_402_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_402_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_402_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_402_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_402_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_402_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_402_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_402_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_402_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_402_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_402_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_402_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_402_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_402_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_402_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_402_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_402_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_402_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_402_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_402_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_402_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_402_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_402_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_402_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_402_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_402_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_402_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_402_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_402_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_402_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_402_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_403_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_403_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_403_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_403_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_403_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_403_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_403_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_403_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_403_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_403_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_403_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_403_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_403_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_403_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_403_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_403_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_403_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_403_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_403_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_403_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_403_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_403_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_403_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_403_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_403_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_403_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_403_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_403_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_403_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_403_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_403_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_404_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_404_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_404_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_404_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_404_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_404_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_404_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_404_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_404_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_404_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_404_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_404_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_404_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_404_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_404_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_404_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_404_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_404_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_404_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_404_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_404_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_404_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_404_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_404_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_404_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_404_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_404_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_404_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_404_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_404_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_404_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_404_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_404_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_404_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_404_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_404_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_404_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_404_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_404_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_405_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_405_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_405_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_405_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_405_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_405_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_405_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_405_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_405_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_405_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_405_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_405_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_405_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_405_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_405_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_405_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_405_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_405_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_405_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_405_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_405_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_405_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_405_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_405_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_405_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_405_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_405_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_405_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_405_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_405_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_405_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_405_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_405_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_405_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_405_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_405_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_406_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_406_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_406_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_406_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_406_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_406_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_406_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_406_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_406_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_406_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_406_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_406_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_406_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_406_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_406_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_406_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_406_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_406_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_406_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_406_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_406_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_406_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_406_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_406_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_406_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_406_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_406_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_406_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_406_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_406_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_406_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_406_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_406_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_406_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_406_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_406_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_406_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_406_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_406_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_406_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_406_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_407_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_407_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_407_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_407_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_407_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_407_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_407_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_407_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_407_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_407_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_407_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_407_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_407_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_407_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_407_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_407_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_407_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_407_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_407_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_407_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_407_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_407_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_408_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_408_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_408_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_408_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_408_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_408_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_408_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_408_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_408_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_408_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_408_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_408_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_408_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_408_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_408_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_408_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_408_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_408_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_409_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_409_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_409_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_409_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_409_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_409_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_409_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_409_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_409_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_409_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_409_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_409_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_409_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_409_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_409_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_409_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_409_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_409_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_409_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_409_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_409_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_409_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_409_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_409_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_409_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_409_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_409_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_409_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_410_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_410_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_410_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_410_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_410_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_410_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_410_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_410_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_410_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_410_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_410_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_410_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_410_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_410_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_410_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_410_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_410_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_410_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_410_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_410_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_410_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_410_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_410_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_410_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_410_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_410_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_410_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_411_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_411_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_411_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_411_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_411_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_411_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_411_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_411_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_411_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_411_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_411_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_411_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_411_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_411_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_411_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_411_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_411_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_411_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_411_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_411_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_411_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_411_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_411_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_411_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_411_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_411_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_411_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_411_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_411_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_411_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_411_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_411_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_411_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_411_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_411_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_411_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_411_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_411_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_411_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_411_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_411_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_412_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_412_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_412_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_412_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_412_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_412_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_412_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_412_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_412_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_412_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_412_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_412_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_412_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_412_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_412_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_412_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_412_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_412_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_412_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_412_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_412_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_412_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_412_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_412_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_412_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_412_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_412_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_412_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_412_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_412_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_412_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_412_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_412_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_412_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_412_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_412_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_412_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_412_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_412_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_412_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_413_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_413_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_413_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_413_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_413_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_413_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_413_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_413_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_413_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_413_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_413_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_413_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_413_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_413_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_413_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_413_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_413_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_413_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_413_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_413_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_413_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_413_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_413_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_413_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_413_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_413_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_413_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_413_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_413_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_413_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_413_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_413_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_413_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_414_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_414_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_414_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_414_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_414_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_414_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_414_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_414_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_414_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_414_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_414_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_414_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_414_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_414_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_414_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_414_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_414_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_414_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_414_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_414_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_414_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_414_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_414_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_414_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_414_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_414_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_414_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_414_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_414_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_414_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_415_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_415_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_415_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_415_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_415_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_415_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_415_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_415_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_415_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_415_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_415_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_415_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_415_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_415_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_415_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_415_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_415_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_415_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_415_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_415_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_415_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_415_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_415_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_415_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_416_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_416_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_416_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_416_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_416_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_416_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_416_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_416_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_416_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_416_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_416_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_416_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_416_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_416_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_416_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_416_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_416_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_416_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_416_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_416_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_416_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_416_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_416_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_416_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_416_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_416_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_416_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_416_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_416_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_416_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_416_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_417_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_417_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_417_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_417_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_417_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_417_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_417_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_417_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_417_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_417_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_417_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_417_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_417_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_417_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_417_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_417_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_417_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_417_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_417_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_417_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_417_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_417_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_417_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_417_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_417_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_417_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_417_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_417_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_417_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_417_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_417_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_417_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_418_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_418_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_418_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_418_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_418_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_418_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_418_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_418_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_418_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_418_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_418_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_418_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_418_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_418_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_418_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_418_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_418_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_418_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_418_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_418_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_418_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_418_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_418_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_418_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_418_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_419_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_419_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_419_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_419_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_419_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_419_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_419_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_419_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_419_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_419_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_419_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_419_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_419_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_419_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_419_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_419_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_419_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_419_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_419_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_419_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_419_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_419_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_419_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_419_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_41_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_420_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_420_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_420_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_420_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_420_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_420_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_420_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_420_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_420_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_420_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_420_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_420_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_420_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_420_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_420_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_420_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_420_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_420_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_420_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_420_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_420_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_420_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_420_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_420_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_420_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_420_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_420_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_420_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_421_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_421_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_421_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_421_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_421_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_421_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_421_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_421_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_421_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_421_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_421_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_421_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_421_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_421_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_421_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_421_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_421_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_421_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_421_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_421_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_421_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_421_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_421_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_421_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_421_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_421_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_421_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_421_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_421_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_421_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_421_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_421_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_421_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_421_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_421_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_421_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_421_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_421_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_422_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_422_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_422_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_422_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_422_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_422_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_422_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_422_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_422_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_422_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_422_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_422_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_422_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_422_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_422_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_422_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_422_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_422_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_422_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_422_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_422_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_422_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_422_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_422_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_422_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_422_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_422_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_422_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_422_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_422_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_422_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_422_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_422_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_422_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_422_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_422_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_422_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_422_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_422_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_422_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_422_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_422_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_422_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_422_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_422_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_423_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_423_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_423_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_423_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_423_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_423_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_423_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_423_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_423_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_423_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_423_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_423_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_423_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_423_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_423_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_423_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_423_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_423_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_423_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_423_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_423_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_423_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_423_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_423_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_423_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_424_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_424_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_424_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_424_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_424_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_424_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_424_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_424_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_424_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_424_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_424_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_424_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_424_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_424_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_424_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_424_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_424_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_424_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_424_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_424_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_424_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_424_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_424_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_424_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_424_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_424_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_424_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_424_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_424_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_424_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_425_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_425_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_425_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_425_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_425_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_425_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_425_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_425_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_425_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_425_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_425_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_425_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_425_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_425_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_425_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_425_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_425_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_425_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_425_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_425_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_425_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_425_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_425_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_425_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_425_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_425_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_425_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_425_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_425_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_425_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_426_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_426_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_426_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_426_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_426_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_426_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_426_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_426_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_426_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_426_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_426_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_426_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_426_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_426_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_426_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_426_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_426_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_426_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_426_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_426_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_426_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_426_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_426_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_426_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_426_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_426_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_426_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_426_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_426_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_426_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_426_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_427_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_427_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_427_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_427_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_427_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_427_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_427_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_427_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_427_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_427_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_427_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_427_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_427_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_427_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_427_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_427_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_427_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_427_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_427_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_427_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_427_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_427_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_427_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_427_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_427_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_427_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_427_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_427_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_427_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_427_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_427_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_427_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_428_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_428_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_428_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_428_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_428_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_428_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_428_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_428_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_428_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_428_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_428_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_428_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_428_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_428_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_428_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_428_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_428_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_428_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_428_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_428_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_428_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_428_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_428_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_428_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_428_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_428_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_428_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_428_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_428_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_428_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_428_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_428_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_428_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_429_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_429_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_429_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_429_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_429_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_429_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_429_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_429_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_429_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_429_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_429_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_429_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_429_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_429_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_429_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_429_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_429_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_429_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_429_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_429_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_429_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_429_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_429_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_429_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_429_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_429_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_429_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_429_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_429_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_429_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_429_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_429_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_429_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_429_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_429_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_429_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_429_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_429_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_430_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_430_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_430_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_430_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_430_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_430_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_430_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_430_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_430_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_430_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_430_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_430_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_430_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_430_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_430_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_430_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_430_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_430_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_430_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_430_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_430_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_430_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_430_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_430_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_430_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_430_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_430_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_430_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_430_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_430_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_430_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_430_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_430_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_431_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_431_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_431_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_431_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_431_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_431_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_431_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_431_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_431_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_431_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_431_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_431_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_431_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_431_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_431_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_431_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_431_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_431_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_431_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_431_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_431_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_431_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_431_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_431_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_431_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_431_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_431_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_431_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_431_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_431_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_431_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_431_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_431_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_431_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_431_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_431_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_431_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_431_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_431_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_431_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_431_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_431_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_431_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_432_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_432_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_432_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_432_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_432_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_432_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_432_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_432_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_432_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_432_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_432_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_432_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_432_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_432_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_432_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_432_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_432_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_432_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_432_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_432_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_432_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_432_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_432_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_432_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_432_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_432_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_432_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_432_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_432_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_432_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_433_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_433_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_433_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_433_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_433_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_433_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_433_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_433_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_433_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_433_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_433_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_433_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_433_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_433_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_433_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_433_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_433_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_433_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_433_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_433_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_433_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_433_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_433_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_433_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_433_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_433_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_433_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_433_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_433_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_433_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_433_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_433_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_433_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_433_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_433_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_433_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_434_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_434_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_434_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_434_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_434_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_434_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_434_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_434_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_434_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_434_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_434_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_434_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_434_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_434_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_434_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_434_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_434_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_434_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_434_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_434_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_434_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_434_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_434_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_434_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_434_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_434_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_434_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_434_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_434_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_434_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_434_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_434_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_434_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_434_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_434_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_434_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_435_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_435_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_435_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_435_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_435_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_435_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_435_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_435_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_435_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_435_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_435_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_435_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_435_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_435_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_435_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_435_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_435_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_435_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_435_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_435_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_435_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_435_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_435_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_435_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_435_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_435_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_435_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_436_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_436_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_436_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_436_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_436_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_436_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_436_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_436_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_436_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_436_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_436_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_436_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_436_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_436_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_436_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_436_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_436_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_436_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_436_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_436_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_436_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_436_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_436_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_436_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_436_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_436_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_436_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_436_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_436_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_437_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_437_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_437_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_437_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_437_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_437_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_437_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_437_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_437_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_437_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_437_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_437_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_437_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_437_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_437_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_437_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_437_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_437_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_437_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_437_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_437_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_437_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_437_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_437_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_437_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_437_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_437_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_437_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_437_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_437_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_437_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_437_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_437_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_437_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_437_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_437_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_437_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_437_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_437_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_437_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_438_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_438_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_438_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_438_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_438_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_438_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_438_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_438_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_438_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_438_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_438_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_438_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_438_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_438_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_438_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_438_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_438_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_438_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_438_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_438_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_438_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_438_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_438_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_438_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_438_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_438_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_438_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_438_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_438_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_438_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_438_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_438_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_438_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_438_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_438_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_438_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_438_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_438_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_438_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_439_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_439_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_439_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_439_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_439_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_439_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_439_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_439_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_439_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_439_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_439_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_439_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_439_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_439_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_439_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_439_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_439_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_439_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_439_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_439_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_439_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_439_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_439_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_439_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_439_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_439_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_439_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_439_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_439_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_439_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_439_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_439_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_439_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_439_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_439_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_43_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_440_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_440_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_440_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_440_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_440_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_440_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_440_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_440_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_440_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_440_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_440_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_440_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_440_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_440_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_440_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_440_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_440_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_440_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_440_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_440_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_440_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_440_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_440_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_440_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_440_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_440_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_440_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_440_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_441_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_441_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_441_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_441_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_441_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_441_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_441_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_441_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_441_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_441_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_441_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_441_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_441_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_441_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_441_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_441_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_441_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_441_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_441_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_441_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_441_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_441_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_441_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_441_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_441_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_441_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_441_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_441_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_441_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_441_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_441_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_441_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_442_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_442_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_442_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_442_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_442_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_442_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_442_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_442_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_442_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_442_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_442_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_442_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_442_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_442_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_442_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_442_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_442_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_442_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_442_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_442_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_442_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_442_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_442_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_442_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_442_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_442_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_442_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_442_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_442_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_443_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_443_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_443_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_443_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_443_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_443_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_443_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_443_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_443_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_443_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_443_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_443_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_443_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_443_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_443_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_443_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_443_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_443_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_443_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_444_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_444_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_444_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_444_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_444_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_444_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_444_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_444_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_444_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_444_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_444_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_444_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_444_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_444_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_444_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_444_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_444_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_444_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_444_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_444_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_444_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_444_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_444_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_444_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_444_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_444_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_444_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_444_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_444_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_444_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_444_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_444_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_444_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_444_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_445_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_445_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_445_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_445_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_445_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_445_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_445_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_445_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_445_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_445_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_445_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_445_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_445_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_445_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_445_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_445_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_445_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_445_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_445_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_445_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_445_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_445_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_445_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_445_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_445_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_445_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_445_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_445_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_445_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_445_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_445_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_445_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_445_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_446_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_446_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_446_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_446_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_446_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_446_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_446_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_446_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_446_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_446_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_446_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_446_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_446_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_446_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_446_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_446_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_446_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_446_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_446_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_446_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_446_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_446_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_446_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_446_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_446_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_446_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_446_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_446_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_446_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_446_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_446_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_446_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_446_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_446_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_446_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_446_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_446_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_446_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_446_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_446_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_446_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_447_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_447_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_447_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_447_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_447_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_447_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_447_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_447_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_447_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_447_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_447_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_447_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_447_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_447_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_447_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_447_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_447_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_447_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_447_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_447_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_447_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_447_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_447_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_447_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_447_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_447_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_447_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_447_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_447_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_447_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_447_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_447_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_447_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_447_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_447_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_447_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_447_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_447_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_447_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_447_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_448_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_448_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_448_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_448_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_448_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_448_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_448_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_448_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_448_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_448_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_448_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_448_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_448_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_448_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_448_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_448_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_448_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_448_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_448_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_448_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_448_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_448_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_448_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_448_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_448_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_448_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_448_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_448_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_448_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_448_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_448_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_448_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_449_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_449_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_449_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_449_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_449_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_449_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_449_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_449_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_449_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_449_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_449_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_449_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_449_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_449_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_449_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_449_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_449_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_449_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_449_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_449_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_449_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_449_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_449_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_449_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_449_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_449_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_449_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_450_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_450_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_450_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_450_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_450_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_450_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_450_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_450_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_450_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_450_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_450_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_450_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_450_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_450_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_450_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_450_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_450_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_450_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_450_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_450_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_450_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_450_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_450_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_450_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_450_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_450_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_450_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_451_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_451_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_451_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_451_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_451_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_451_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_451_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_451_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_451_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_451_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_451_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_451_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_451_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_451_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_451_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_451_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_451_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_451_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_451_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_451_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_451_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_451_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_451_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_451_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_451_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_451_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_451_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_451_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_451_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_451_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_451_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_451_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_451_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_451_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_451_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_452_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_452_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_452_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_452_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_452_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_452_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_452_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_452_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_452_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_452_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_452_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_452_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_452_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_452_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_452_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_452_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_452_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_452_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_452_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_452_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_452_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_452_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_452_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_452_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_452_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_452_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_452_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_452_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_452_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_452_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_452_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_452_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_452_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_452_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_452_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_452_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_453_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_453_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_453_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_453_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_453_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_453_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_453_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_453_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_453_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_453_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_453_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_453_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_453_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_453_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_453_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_453_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_453_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_453_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_453_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_453_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_453_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_453_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_453_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_453_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_453_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_453_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_453_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_453_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_453_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_454_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_454_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_454_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_454_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_454_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_454_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_454_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_454_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_454_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_454_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_454_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_454_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_454_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_454_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_454_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_454_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_454_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_454_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_454_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_454_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_454_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_454_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_454_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_454_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_454_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_454_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_454_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_454_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_454_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_454_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_454_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_454_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_454_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_454_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_454_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_454_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_454_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_454_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_454_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_454_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_454_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_454_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_454_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_454_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_454_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_454_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_454_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_454_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_454_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_454_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_455_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_455_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_455_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_455_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_455_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_455_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_455_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_455_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_455_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_455_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_455_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_455_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_455_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_455_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_455_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_455_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_455_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_455_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_455_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_455_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_455_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_455_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_455_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_455_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_455_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_455_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_455_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_455_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_455_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_455_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_455_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_455_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_455_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_455_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_455_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_455_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_455_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_455_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_455_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_455_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_455_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_455_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_456_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_456_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_456_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_456_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_456_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_456_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_456_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_456_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_456_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_456_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_456_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_456_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_456_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_456_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_456_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_456_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_456_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_456_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_456_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_456_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_456_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_456_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_456_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_456_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_456_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_456_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_456_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_456_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_456_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_456_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_456_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_456_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_456_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_456_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_456_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_456_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_456_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_456_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_456_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_456_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_456_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_456_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_457_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_457_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_457_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_457_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_457_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_457_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_457_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_457_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_457_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_457_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_457_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_457_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_457_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_457_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_457_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_457_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_457_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_457_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_457_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_457_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_457_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_457_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_457_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_457_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_457_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_457_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_457_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_457_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_457_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_457_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_457_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_457_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_457_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_457_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_457_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_457_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_457_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_457_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_457_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_457_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_457_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_458_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_458_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_458_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_458_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_458_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_458_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_458_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_458_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_458_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_458_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_458_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_458_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_458_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_458_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_458_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_458_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_458_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_458_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_458_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_458_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_458_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_458_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_458_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_458_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_458_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_458_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_458_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_458_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_458_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_458_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_458_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_459_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_459_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_459_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_459_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_459_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_459_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_459_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_459_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_459_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_459_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_459_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_459_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_459_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_459_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_459_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_459_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_459_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_459_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_459_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_459_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_459_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_459_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_459_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_459_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_459_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_459_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_459_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_459_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_459_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_460_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_460_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_460_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_460_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_460_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_460_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_460_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_460_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_460_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_460_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_460_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_460_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_460_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_460_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_460_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_460_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_460_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_460_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_460_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_460_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_460_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_460_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_460_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_460_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_460_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_460_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_460_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_461_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_461_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_461_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_461_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_461_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_461_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_461_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_461_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_461_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_461_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_461_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_461_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_461_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_461_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_461_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_461_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_461_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_461_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_461_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_461_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_461_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_461_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_461_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_461_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_461_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_461_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_461_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_461_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_461_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_461_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_461_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_461_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_461_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_461_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_461_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_461_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_461_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_461_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_461_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_462_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_462_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_462_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_462_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_462_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_462_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_462_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_462_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_462_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_462_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_462_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_462_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_462_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_462_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_462_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_462_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_462_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_462_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_462_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_462_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_462_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_462_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_462_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_462_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_462_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_462_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_462_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_462_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_462_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_462_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_462_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_462_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_462_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_462_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_462_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_462_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_462_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_462_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_462_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_463_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_463_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_463_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_463_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_463_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_463_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_463_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_463_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_463_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_463_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_463_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_463_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_463_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_463_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_463_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_463_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_463_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_463_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_463_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_463_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_463_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_463_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_463_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_463_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_463_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_463_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_463_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_463_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_463_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_463_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_463_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_464_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_464_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_464_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_464_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_464_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_464_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_464_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_464_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_464_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_464_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_464_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_464_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_464_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_464_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_464_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_464_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_464_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_464_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_464_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_464_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_464_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_464_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_464_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_464_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_464_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_464_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_464_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_465_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_465_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_465_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_465_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_465_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_465_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_465_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_465_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_465_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_465_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_465_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_465_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_465_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_465_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_465_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_465_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_465_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_465_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_465_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_465_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_465_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_465_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_465_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_465_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_465_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_465_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_465_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_465_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_465_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_465_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_465_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_466_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_466_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_466_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_466_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_466_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_466_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_466_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_466_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_466_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_466_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_466_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_466_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_466_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_466_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_466_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_466_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_466_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_466_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_466_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_466_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_466_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_466_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_466_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_466_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_466_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_466_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_466_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_466_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_466_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_466_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_466_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_466_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_466_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_466_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_466_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_466_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_466_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_467_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_467_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_467_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_467_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_467_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_467_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_467_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_467_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_467_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_467_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_467_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_467_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_467_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_467_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_467_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_467_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_467_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_467_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_467_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_467_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_467_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_467_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_467_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_467_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_467_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_467_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_467_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_468_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_468_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_468_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_468_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_468_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_468_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_468_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_468_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_468_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_468_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_468_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_468_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_468_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_468_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_468_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_468_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_468_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_468_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_468_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_468_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_468_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_468_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_469_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_469_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_469_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_469_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_469_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_469_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_469_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_469_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_469_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_469_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_469_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_469_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_469_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_469_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_469_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_469_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_469_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_469_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_469_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_469_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_469_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_469_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_469_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_469_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_469_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_469_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_469_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_469_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_469_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_469_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_469_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_469_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_469_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_470_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_470_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_470_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_470_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_470_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_470_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_470_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_470_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_470_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_470_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_470_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_470_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_470_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_470_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_470_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_470_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_470_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_470_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_470_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_470_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_470_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_470_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_470_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_470_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_470_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_470_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_470_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_470_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_470_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_470_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_470_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_471_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_471_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_471_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_471_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_471_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_471_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_471_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_471_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_471_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_471_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_471_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_471_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_471_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_471_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_471_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_471_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_471_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_471_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_471_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_471_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_471_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_471_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_471_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_471_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_471_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_471_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_471_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_471_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_471_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_472_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_472_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_472_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_472_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_472_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_472_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_472_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_472_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_472_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_472_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_472_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_472_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_472_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_472_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_472_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_472_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_472_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_472_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_472_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_472_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_472_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_472_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_472_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_472_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_472_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_472_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_472_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_472_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_472_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_473_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_473_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_473_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_473_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_473_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_473_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_473_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_473_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_473_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_473_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_473_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_473_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_473_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_473_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_473_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_473_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_473_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_473_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_473_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_473_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_473_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_473_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_473_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_473_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_473_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_473_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_473_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_473_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_473_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_473_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_473_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_473_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_473_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_473_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_474_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_474_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_474_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_474_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_474_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_474_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_474_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_474_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_474_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_474_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_474_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_474_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_474_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_474_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_474_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_474_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_474_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_474_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_474_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_474_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_474_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_474_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_474_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_474_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_474_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_474_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_474_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_474_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_474_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_474_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_474_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_474_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_474_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_474_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_474_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_474_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_474_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_474_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_474_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_474_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_474_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_474_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_475_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_475_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_475_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_475_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_475_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_475_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_475_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_475_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_475_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_475_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_475_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_475_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_475_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_475_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_475_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_475_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_475_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_475_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_475_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_475_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_475_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_475_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_475_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_475_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_475_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_475_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_475_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_475_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_475_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_475_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_475_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_475_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_475_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_475_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_475_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_476_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_476_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_476_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_476_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_476_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_476_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_476_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_476_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_476_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_476_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_476_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_476_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_476_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_476_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_476_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_476_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_476_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_476_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_476_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_476_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_476_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_476_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_476_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_476_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_476_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_476_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_476_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_476_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_476_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_476_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_476_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_476_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_476_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_476_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_477_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_477_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_477_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_477_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_477_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_477_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_477_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_477_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_477_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_477_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_477_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_477_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_477_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_477_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_477_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_477_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_477_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_477_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_477_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_477_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_477_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_477_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_477_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_477_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_477_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_477_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_477_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_477_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_477_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_477_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_477_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_477_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_477_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_477_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_477_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_477_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_477_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_477_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_477_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_478_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_478_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_478_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_478_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_478_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_478_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_478_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_478_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_478_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_478_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_478_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_478_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_478_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_478_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_478_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_478_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_478_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_478_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_478_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_478_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_478_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_478_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_478_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_478_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_478_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_478_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_478_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_478_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_478_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_478_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_478_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_478_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_479_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_479_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_479_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_479_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_479_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_479_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_479_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_479_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_479_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_479_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_479_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_479_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_479_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_479_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_479_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_479_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_479_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_479_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_479_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_479_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_479_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_479_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_479_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_479_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_479_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_47_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_47_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_480_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_480_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_480_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_480_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_480_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_480_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_480_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_480_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_480_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_480_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_480_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_480_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_480_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_480_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_480_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_480_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_480_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_480_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_480_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_480_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_481_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_481_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_481_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_481_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_481_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_481_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_481_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_481_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_481_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_481_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_481_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_481_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_481_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_481_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_481_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_481_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_481_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_481_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_481_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_481_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_481_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_481_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_481_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_481_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_481_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_481_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_481_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_481_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_481_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_482_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_482_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_482_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_482_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_482_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_482_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_482_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_482_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_482_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_482_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_482_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_482_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_482_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_482_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_482_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_482_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_482_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_482_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_482_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_482_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_482_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_482_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_482_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_482_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_482_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_482_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_482_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_482_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_482_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_483_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_483_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_483_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_483_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_483_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_483_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_483_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_483_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_483_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_483_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_483_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_483_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_483_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_483_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_483_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_483_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_483_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_483_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_483_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_483_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_483_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_483_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_483_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_483_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_483_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_483_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_483_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_483_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_483_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_483_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_483_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_483_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_483_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_483_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_483_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_483_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_483_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_484_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_484_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_484_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_484_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_484_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_484_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_484_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_484_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_484_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_484_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_484_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_484_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_484_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_484_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_484_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_484_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_484_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_484_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_484_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_484_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_484_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_484_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_484_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_484_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_484_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_484_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_484_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_484_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_484_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_484_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_484_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_484_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_484_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_484_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_484_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_485_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_485_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_485_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_485_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_485_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_485_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_485_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_485_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_485_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_485_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_485_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_485_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_485_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_485_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_485_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_485_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_485_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_485_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_485_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_485_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_485_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_485_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_485_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_485_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_485_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_485_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_485_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_485_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_485_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_485_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_485_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_486_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_486_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_486_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_486_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_486_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_486_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_486_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_486_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_486_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_486_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_486_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_486_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_486_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_486_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_486_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_486_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_486_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_486_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_486_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_486_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_486_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_486_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_486_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_486_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_486_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_486_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_486_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_486_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_486_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_486_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_486_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_486_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_486_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_486_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_486_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_486_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_486_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_486_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_486_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_486_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_486_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_486_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_486_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_487_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_487_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_487_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_487_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_487_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_487_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_487_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_487_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_487_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_487_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_487_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_487_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_487_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_487_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_487_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_487_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_487_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_487_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_487_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_487_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_487_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_487_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_487_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_487_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_487_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_487_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_487_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_487_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_487_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_487_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_487_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_487_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_487_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_487_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_487_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_487_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_487_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_488_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_488_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_488_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_488_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_488_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_488_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_488_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_488_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_488_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_488_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_488_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_488_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_488_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_488_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_488_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_488_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_488_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_488_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_488_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_488_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_488_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_488_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_488_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_488_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_488_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_488_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_488_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_489_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_489_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_489_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_489_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_489_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_489_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_489_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_489_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_489_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_489_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_489_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_489_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_489_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_489_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_489_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_489_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_489_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_489_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_489_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_489_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_489_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_489_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_489_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_489_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_489_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_48_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_490_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_490_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_490_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_490_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_490_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_490_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_490_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_490_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_490_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_490_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_490_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_490_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_490_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_490_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_490_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_490_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_490_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_490_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_490_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_490_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_490_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_490_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_490_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_490_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_490_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_490_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_491_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_491_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_491_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_491_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_491_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_491_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_491_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_491_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_491_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_491_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_491_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_491_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_491_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_491_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_491_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_491_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_491_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_491_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_491_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_491_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_491_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_491_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_491_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_492_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_492_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_492_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_492_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_492_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_492_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_492_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_492_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_492_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_492_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_492_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_492_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_492_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_492_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_492_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_492_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_492_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_492_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_492_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_493_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_493_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_493_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_493_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_493_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_493_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_493_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_493_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_493_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_493_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_493_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_493_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_493_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_493_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_493_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_493_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_493_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_493_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_493_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_493_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_493_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_493_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_493_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_493_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_493_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_493_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_493_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_493_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_493_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_493_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_493_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_493_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_493_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_493_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_493_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_493_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_493_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_493_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_493_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_494_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_494_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_494_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_494_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_494_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_494_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_494_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_494_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_494_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_494_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_494_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_494_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_494_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_494_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_494_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_494_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_494_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_494_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_494_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_494_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_494_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_494_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_494_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_494_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_494_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_494_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_494_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_494_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_494_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_494_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_494_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_494_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_494_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_494_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_494_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_494_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_494_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_494_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_494_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_494_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_494_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_494_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_494_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_494_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_494_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_495_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_495_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_495_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_495_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_495_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_495_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_495_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_495_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_495_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_495_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_495_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_495_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_495_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_495_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_495_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_495_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_495_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_495_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_495_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_495_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_495_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_495_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_495_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_495_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_495_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_495_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_495_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_495_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_495_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_495_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_495_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_495_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_495_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_495_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_495_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_495_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_495_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_495_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_495_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_495_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_495_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_495_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_495_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_495_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_495_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_495_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_495_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_495_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_496_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_496_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_496_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_496_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_496_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_496_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_496_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_496_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_496_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_496_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_496_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_496_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_496_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_496_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_496_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_496_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_496_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_496_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_496_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_496_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_496_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_496_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_496_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_496_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_496_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_496_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_496_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_496_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_496_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_496_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_496_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_496_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_496_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_496_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_496_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_496_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_496_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_496_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_496_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_496_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_496_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_496_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_496_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_497_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_497_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_497_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_497_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_497_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_497_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_497_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_497_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_497_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_497_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_497_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_497_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_497_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_497_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_497_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_497_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_497_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_497_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_497_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_497_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_497_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_497_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_497_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_497_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_497_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_497_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_497_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_497_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_497_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_497_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_497_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_498_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_498_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_498_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_498_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_498_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_498_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_498_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_498_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_498_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_498_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_498_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_498_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_498_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_498_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_498_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_498_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_498_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_498_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_498_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_498_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_498_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_498_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_499_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_499_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_499_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_499_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_499_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_499_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_499_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_499_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_499_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_499_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_499_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_499_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_499_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_499_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_499_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_499_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_499_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_499_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_499_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_499_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_499_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_499_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_499_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_499_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_499_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_499_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_499_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_499_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_499_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_499_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_499_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_499_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_499_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_49_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_49_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_500_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_500_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_500_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_500_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_500_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_500_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_500_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_500_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_500_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_500_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_500_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_500_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_500_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_500_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_500_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_500_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_500_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_500_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_500_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_500_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_500_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_501_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_501_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_501_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_501_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_501_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_501_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_501_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_501_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_501_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_501_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_501_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_501_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_501_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_501_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_501_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_501_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_501_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_501_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_501_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_501_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_501_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_501_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_501_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_501_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_502_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_502_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_502_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_502_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_502_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_502_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_502_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_502_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_502_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_502_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_502_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_502_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_502_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_502_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_502_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_502_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_502_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_502_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_502_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_502_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_502_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_502_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_502_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_502_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_502_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_502_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_502_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_502_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_502_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_503_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_503_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_503_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_503_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_503_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_503_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_503_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_503_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_503_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_503_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_503_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_503_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_503_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_503_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_503_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_503_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_503_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_503_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_503_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_503_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_503_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_503_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_503_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_503_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_503_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_503_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_503_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_503_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_503_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_503_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_503_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_503_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_503_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_503_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_503_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_503_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_503_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_503_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_503_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_503_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_503_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_503_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_503_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_503_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_504_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_504_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_504_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_504_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_504_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_504_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_504_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_504_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_504_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_504_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_504_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_504_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_504_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_504_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_504_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_504_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_504_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_504_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_504_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_504_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_504_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_504_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_504_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_504_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_504_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_504_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_504_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_504_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_504_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_504_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_504_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_504_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_504_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_504_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_504_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_504_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_504_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_504_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_504_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_504_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_504_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_505_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_505_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_505_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_505_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_505_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_505_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_505_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_505_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_505_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_505_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_505_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_505_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_505_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_505_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_505_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_505_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_505_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_505_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_505_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_505_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_505_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_505_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_505_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_505_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_505_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_505_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_505_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_505_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_505_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_505_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_505_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_505_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_505_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_505_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_505_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_505_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_505_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_505_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_505_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_505_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_505_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_505_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_505_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_505_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_505_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_505_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_506_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_506_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_506_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_506_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_506_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_506_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_506_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_506_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_506_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_506_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_506_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_506_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_506_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_506_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_506_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_506_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_506_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_506_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_506_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_506_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_506_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_506_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_506_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_506_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_506_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_506_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_506_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_506_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_506_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_506_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_506_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_506_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_506_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_506_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_506_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_506_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_506_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_506_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_506_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_507_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_507_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_507_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_507_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_507_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_507_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_507_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_507_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_507_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_507_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_507_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_507_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_507_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_507_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_507_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_507_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_507_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_507_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_507_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_507_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_507_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_507_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_507_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_507_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_507_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_507_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_507_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_507_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_507_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_507_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_508_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_508_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_508_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_508_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_508_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_508_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_508_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_508_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_508_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_508_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_508_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_508_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_508_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_508_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_508_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_508_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_508_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_508_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_508_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_508_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_508_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_508_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_508_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_508_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_509_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_509_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_509_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_509_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_509_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_509_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_509_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_509_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_509_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_509_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_509_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_509_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_509_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_509_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_509_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_509_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_509_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_509_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_509_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_509_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_509_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_509_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_50_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_50_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_510_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_510_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_510_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_510_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_510_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_510_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_510_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_510_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_510_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_510_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_510_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_510_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_510_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_510_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_510_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_510_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_510_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_510_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_511_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_511_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_511_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_511_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_511_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_511_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_511_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_511_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_511_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_511_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_511_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_511_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_511_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_511_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_511_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_511_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_511_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_511_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_511_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_511_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_511_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_511_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_511_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_511_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_511_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_511_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_511_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_511_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_511_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_512_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_512_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_512_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_512_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_512_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_512_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_512_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_512_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_512_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_512_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_512_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_512_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_512_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_512_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_512_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_512_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_512_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_512_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_512_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_512_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_512_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_512_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_512_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_512_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_512_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_512_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_512_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_512_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_512_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_512_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_512_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_512_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_512_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_512_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_512_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_512_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_512_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_512_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_513_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_513_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_513_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_513_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_513_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_513_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_513_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_513_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_513_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_513_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_513_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_513_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_513_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_513_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_513_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_513_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_513_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_513_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_513_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_513_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_513_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_513_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_513_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_513_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_513_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_513_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_513_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_513_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_513_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_513_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_513_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_513_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_513_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_513_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_513_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_513_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_513_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_514_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_514_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_514_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_514_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_514_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_514_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_514_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_514_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_514_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_514_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_514_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_514_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_514_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_514_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_514_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_514_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_514_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_514_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_514_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_514_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_514_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_514_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_514_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_514_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_514_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_514_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_514_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_514_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_514_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_514_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_514_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_514_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_515_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_515_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_515_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_515_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_515_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_515_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_515_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_515_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_515_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_515_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_515_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_515_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_515_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_515_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_515_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_515_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_515_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_515_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_515_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_515_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_515_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_515_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_515_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_515_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_515_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_515_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_515_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_515_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_515_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_515_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_515_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_515_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_515_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_515_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_515_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_515_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_515_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_515_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_515_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_515_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_515_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_515_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_515_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_515_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_516_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_516_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_516_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_516_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_516_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_516_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_516_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_516_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_516_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_516_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_516_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_516_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_516_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_516_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_516_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_516_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_516_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_516_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_516_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_516_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_516_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_516_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_516_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_516_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_516_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_516_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_517_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_517_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_517_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_517_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_517_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_517_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_517_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_517_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_517_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_517_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_517_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_517_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_517_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_517_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_517_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_517_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_517_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_517_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_517_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_517_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_517_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_517_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_517_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_517_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_517_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_517_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_517_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_517_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_517_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_517_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_517_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_517_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_517_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_517_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_517_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_517_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_517_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_517_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_517_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_517_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_517_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_518_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_518_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_518_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_518_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_518_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_518_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_518_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_518_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_518_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_518_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_518_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_518_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_518_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_518_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_518_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_518_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_518_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_518_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_518_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_518_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_518_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_518_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_518_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_518_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_518_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_518_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_518_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_518_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_518_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_518_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_518_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_518_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_518_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_518_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_518_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_518_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_518_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_518_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_518_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_519_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_519_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_519_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_519_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_519_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_519_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_519_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_519_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_519_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_519_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_519_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_519_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_519_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_519_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_519_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_519_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_519_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_519_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_519_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_51_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_51_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_51_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_520_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_520_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_520_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_520_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_520_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_520_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_520_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_520_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_520_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_520_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_520_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_520_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_520_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_520_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_520_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_520_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_520_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_520_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_520_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_520_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_520_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_520_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_520_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_520_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_520_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_521_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_521_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_521_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_521_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_521_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_521_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_521_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_521_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_521_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_521_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_521_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_521_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_521_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_521_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_521_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_521_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_521_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_521_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_521_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_522_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_522_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_522_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_522_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_522_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_522_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_522_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_522_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_522_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_522_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_522_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_522_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_522_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_522_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_522_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_522_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_522_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_522_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_522_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_522_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_522_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_522_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_522_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_522_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_522_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_522_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_522_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_522_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_523_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_523_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_523_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_523_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_523_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_523_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_523_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_523_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_523_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_523_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_523_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_523_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_523_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_523_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_523_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_523_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_523_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_523_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_523_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_523_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_523_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_523_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_523_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_523_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_523_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_523_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_523_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_523_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_523_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_523_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_523_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_523_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_523_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_523_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_524_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_524_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_524_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_524_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_524_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_524_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_524_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_524_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_524_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_524_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_524_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_524_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_524_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_524_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_524_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_524_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_524_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_524_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_524_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_524_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_524_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_524_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_524_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_524_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_524_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_524_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_524_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_524_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_524_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_524_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_524_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_524_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_524_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_524_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_524_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_524_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_524_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_524_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_524_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_524_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_524_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_524_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_525_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_525_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_525_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_525_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_525_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_525_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_525_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_525_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_525_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_525_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_525_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_525_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_525_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_525_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_525_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_525_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_525_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_525_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_525_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_525_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_525_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_525_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_525_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_525_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_525_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_525_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_526_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_526_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_526_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_526_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_526_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_526_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_526_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_526_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_526_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_526_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_526_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_526_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_526_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_526_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_526_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_526_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_526_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_526_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_526_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_526_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_526_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_526_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_526_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_526_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_526_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_526_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_526_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_526_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_526_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_526_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_526_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_526_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_526_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_526_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_526_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_526_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_526_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_526_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_526_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_526_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_526_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_526_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_526_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_526_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_527_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_527_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_527_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_527_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_527_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_527_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_527_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_527_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_527_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_527_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_527_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_527_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_527_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_527_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_527_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_527_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_527_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_527_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_527_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_527_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_527_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_527_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_527_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_527_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_527_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_527_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_527_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_527_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_527_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_527_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_527_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_527_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_527_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_527_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_527_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_527_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_527_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_527_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_527_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_527_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_527_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_527_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_528_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_528_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_528_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_528_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_528_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_528_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_528_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_528_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_528_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_528_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_528_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_528_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_528_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_528_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_528_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_528_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_528_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_528_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_528_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_528_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_528_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_528_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_528_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_528_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_528_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_528_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_528_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_528_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_528_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_528_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_528_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_528_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_529_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_529_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_529_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_529_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_529_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_529_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_529_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_529_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_529_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_529_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_529_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_529_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_529_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_529_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_529_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_529_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_529_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_529_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_529_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_529_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_529_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_529_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_529_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_529_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_529_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_529_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_529_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_529_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_529_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_52_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_530_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_530_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_530_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_530_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_530_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_530_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_530_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_530_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_530_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_530_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_530_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_530_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_530_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_530_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_530_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_530_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_530_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_530_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_530_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_530_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_530_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_530_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_530_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_530_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_530_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_530_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_530_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_530_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_530_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_531_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_531_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_531_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_531_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_531_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_531_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_531_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_531_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_531_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_531_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_531_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_531_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_531_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_531_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_531_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_531_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_531_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_531_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_531_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_531_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_531_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_531_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_531_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_531_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_531_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_532_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_532_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_532_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_532_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_532_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_532_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_532_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_532_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_532_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_532_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_532_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_532_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_532_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_532_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_532_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_532_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_532_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_532_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_532_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_532_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_532_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_532_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_532_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_532_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_532_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_533_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_533_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_533_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_533_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_533_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_533_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_533_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_533_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_533_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_533_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_533_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_533_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_533_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_533_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_533_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_533_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_533_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_533_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_533_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_533_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_533_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_533_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_533_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_533_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_533_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_533_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_533_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_534_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_534_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_534_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_534_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_534_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_534_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_534_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_534_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_534_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_534_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_534_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_534_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_534_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_534_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_534_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_534_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_534_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_534_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_534_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_534_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_534_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_534_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_534_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_534_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_534_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_534_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_534_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_534_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_534_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_534_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_534_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_534_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_534_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_534_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_535_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_535_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_535_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_535_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_535_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_535_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_535_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_535_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_535_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_535_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_535_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_535_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_535_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_535_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_535_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_535_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_535_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_535_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_535_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_535_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_535_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_535_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_535_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_535_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_535_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_535_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_535_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_535_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_536_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_536_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_536_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_536_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_536_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_536_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_536_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_536_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_536_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_536_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_536_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_536_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_536_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_536_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_536_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_536_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_536_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_536_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_536_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_536_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_536_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_536_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_536_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_536_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_536_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_536_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_536_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_536_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_536_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_536_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_536_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_536_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_536_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_536_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_537_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_537_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_537_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_537_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_537_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_537_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_537_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_537_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_537_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_537_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_537_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_537_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_537_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_537_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_537_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_537_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_537_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_537_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_537_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_537_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_537_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_537_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_537_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_537_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_537_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_537_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_537_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_537_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_537_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_537_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_538_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_538_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_538_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_538_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_538_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_538_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_538_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_538_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_538_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_538_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_538_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_538_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_538_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_538_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_538_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_538_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_538_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_538_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_538_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_538_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_538_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_538_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_538_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_538_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_538_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_538_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_538_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_538_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_538_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_538_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_538_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_538_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_538_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_538_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_538_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_538_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_539_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_539_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_539_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_539_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_539_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_539_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_539_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_539_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_539_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_539_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_539_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_539_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_539_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_539_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_539_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_539_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_539_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_539_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_539_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_539_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_539_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_539_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_539_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_539_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_539_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_53_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_53_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_540_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_540_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_540_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_540_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_540_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_540_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_540_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_540_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_540_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_540_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_540_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_540_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_540_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_540_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_540_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_540_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_540_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_540_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_540_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_540_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_540_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_541_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_541_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_541_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_541_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_541_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_541_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_541_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_541_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_541_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_541_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_541_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_541_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_541_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_541_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_541_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_541_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_541_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_541_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_541_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_541_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_541_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_541_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_541_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_542_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_542_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_542_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_542_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_542_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_542_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_542_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_542_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_542_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_542_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_542_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_542_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_542_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_542_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_542_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_542_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_542_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_542_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_542_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_542_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_542_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_542_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_542_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_542_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_542_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_542_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_543_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_543_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_543_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_543_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_543_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_543_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_543_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_543_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_543_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_543_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_543_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_543_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_543_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_543_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_543_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_543_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_543_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_543_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_543_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_543_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_543_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_543_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_543_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_543_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_543_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_543_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_543_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_543_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_543_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_543_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_543_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_543_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_543_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_544_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_544_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_544_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_544_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_544_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_544_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_544_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_544_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_544_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_544_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_544_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_544_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_544_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_544_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_544_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_544_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_544_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_544_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_544_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_544_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_544_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_544_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_544_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_544_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_544_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_544_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_544_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_544_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_544_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_544_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_544_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_544_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_544_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_544_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_544_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_544_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_544_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_544_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_544_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_544_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_544_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_544_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_544_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_544_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_544_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_544_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_544_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_544_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_545_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_545_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_545_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_545_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_545_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_545_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_545_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_545_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_545_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_545_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_545_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_545_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_545_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_545_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_545_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_545_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_545_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_545_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_545_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_545_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_545_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_545_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_545_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_545_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_545_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_545_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_545_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_545_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_545_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_545_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_545_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_545_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_545_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_545_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_545_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_545_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_546_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_546_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_546_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_546_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_546_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_546_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_546_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_546_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_546_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_546_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_546_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_546_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_546_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_546_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_546_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_546_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_546_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_546_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_546_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_546_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_546_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_546_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_546_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_546_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_546_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_546_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_546_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_546_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_546_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_546_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_546_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_546_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_546_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_546_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_546_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_546_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_546_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_547_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_547_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_547_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_547_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_547_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_547_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_547_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_547_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_547_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_547_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_547_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_547_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_547_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_547_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_547_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_547_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_547_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_547_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_547_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_547_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_547_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_547_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_547_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_547_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_547_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_547_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_547_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_547_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_547_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_547_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_547_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_547_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_548_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_548_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_548_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_548_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_548_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_548_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_548_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_548_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_548_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_548_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_548_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_548_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_548_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_548_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_548_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_548_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_548_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_548_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_548_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_548_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_548_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_548_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_548_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_548_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_549_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_549_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_549_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_549_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_549_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_549_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_549_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_549_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_549_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_549_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_549_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_549_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_549_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_549_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_549_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_549_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_549_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_549_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_549_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_549_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_549_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_549_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_549_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_549_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_549_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_549_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_549_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_549_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_549_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_549_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_549_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_549_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_549_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_549_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_549_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_549_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_549_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_549_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_550_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_550_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_550_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_550_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_550_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_550_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_550_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_550_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_550_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_550_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_550_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_550_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_550_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_550_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_550_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_550_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_550_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_550_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_550_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_550_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_550_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_550_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_550_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_550_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_550_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_550_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_550_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_551_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_551_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_551_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_551_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_551_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_551_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_551_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_551_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_551_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_551_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_551_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_551_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_551_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_551_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_551_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_551_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_551_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_551_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_551_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_551_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_551_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_551_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_551_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_552_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_552_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_552_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_552_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_552_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_552_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_552_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_552_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_552_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_552_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_552_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_552_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_552_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_552_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_552_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_552_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_552_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_552_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_552_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_552_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_552_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_552_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_552_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_552_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_552_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_552_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_552_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_552_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_552_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_552_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_552_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_552_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_552_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_552_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_552_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_552_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_552_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_552_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_552_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_552_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_552_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_552_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_553_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_553_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_553_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_553_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_553_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_553_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_553_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_553_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_553_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_553_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_553_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_553_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_553_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_553_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_553_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_553_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_553_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_553_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_553_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_553_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_553_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_553_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_553_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_553_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_553_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_553_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_553_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_554_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_554_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_554_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_554_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_554_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_554_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_554_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_554_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_554_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_554_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_554_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_554_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_554_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_554_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_554_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_554_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_554_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_554_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_554_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_554_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_554_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_554_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_554_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_554_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_554_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_554_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_554_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_554_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_554_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_555_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_555_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_555_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_555_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_555_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_555_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_555_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_555_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_555_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_555_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_555_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_555_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_555_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_555_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_555_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_555_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_555_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_555_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_555_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_555_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_555_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_555_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_555_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_555_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_555_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_555_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_555_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_556_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_556_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_556_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_556_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_556_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_556_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_556_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_556_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_556_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_556_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_556_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_556_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_556_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_556_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_556_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_556_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_556_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_556_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_556_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_556_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_556_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_556_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_556_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_557_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_557_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_557_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_557_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_557_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_557_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_557_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_557_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_557_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_557_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_557_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_557_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_557_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_557_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_557_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_557_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_557_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_557_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_557_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_557_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_557_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_558_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_558_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_558_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_558_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_558_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_558_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_558_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_558_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_558_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_558_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_558_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_558_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_558_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_558_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_558_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_558_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_558_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_558_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_558_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_558_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_558_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_558_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_558_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_558_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_558_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_558_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_558_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_558_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_558_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_558_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_558_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_559_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_559_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_559_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_559_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_559_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_559_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_559_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_559_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_559_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_559_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_559_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_559_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_559_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_559_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_559_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_559_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_559_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_559_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_559_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_559_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_559_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_559_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_55_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_55_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_560_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_560_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_560_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_560_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_560_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_560_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_560_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_560_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_560_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_560_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_560_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_560_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_560_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_560_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_560_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_560_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_560_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_560_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_560_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_560_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_560_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_560_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_560_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_560_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_560_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_560_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_560_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_560_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_560_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_561_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_561_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_561_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_561_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_561_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_561_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_561_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_561_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_561_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_561_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_561_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_561_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_561_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_561_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_561_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_561_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_561_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_561_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_561_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_561_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_561_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_561_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_561_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_561_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_561_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_561_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_561_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_561_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_561_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_561_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_562_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_562_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_562_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_562_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_562_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_562_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_562_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_562_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_562_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_562_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_562_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_562_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_562_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_562_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_562_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_562_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_562_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_562_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_562_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_562_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_562_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_562_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_563_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_563_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_563_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_563_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_563_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_563_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_563_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_563_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_563_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_563_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_563_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_563_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_563_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_563_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_563_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_563_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_563_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_563_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_563_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_563_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_563_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_563_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_563_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_563_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_563_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_563_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_563_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_563_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_564_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_564_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_564_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_564_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_564_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_564_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_564_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_564_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_564_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_564_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_564_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_564_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_564_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_564_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_564_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_564_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_564_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_564_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_564_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_564_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_564_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_564_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_565_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_565_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_565_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_565_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_565_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_565_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_565_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_565_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_565_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_565_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_565_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_565_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_565_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_565_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_565_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_565_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_565_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_565_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_565_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_565_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_565_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_565_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_565_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_565_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_565_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_565_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_565_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_565_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_565_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_565_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_566_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_566_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_566_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_566_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_566_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_566_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_566_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_566_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_566_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_566_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_566_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_566_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_566_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_566_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_566_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_566_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_566_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_566_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_566_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_566_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_566_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_566_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_566_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_566_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_566_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_566_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_566_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_567_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_567_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_567_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_567_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_567_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_567_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_567_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_567_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_567_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_567_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_567_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_567_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_567_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_567_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_567_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_567_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_567_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_567_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_567_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_567_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_567_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_567_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_567_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_567_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_567_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_567_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_567_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_567_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_567_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_567_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_567_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_567_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_568_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_568_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_568_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_568_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_568_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_568_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_568_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_568_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_568_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_568_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_568_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_568_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_568_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_568_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_568_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_568_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_568_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_568_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_568_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_568_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_568_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_568_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_568_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_568_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_568_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_568_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_569_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_569_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_569_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_569_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_569_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_569_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_569_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_569_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_569_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_569_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_569_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_569_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_569_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_569_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_569_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_569_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_569_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_569_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_569_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_569_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_569_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_569_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_569_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_569_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_569_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_569_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_569_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_56_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_56_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_570_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_570_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_570_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_570_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_570_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_570_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_570_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_570_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_570_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_570_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_570_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_570_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_570_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_570_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_570_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_570_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_570_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_570_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_570_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_570_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_570_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_570_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_570_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_570_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_570_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_570_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_571_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_571_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_571_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_571_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_571_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_571_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_571_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_571_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_571_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_571_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_571_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_571_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_571_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_571_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_571_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_571_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_571_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_571_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_571_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_571_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_571_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_571_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_571_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_571_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_571_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_571_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_572_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_572_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_572_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_572_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_572_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_572_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_572_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_572_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_572_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_572_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_572_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_572_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_572_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_572_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_572_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_572_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_572_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_572_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_572_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_572_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_572_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_572_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_572_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_572_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_572_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_572_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_572_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_572_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_572_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_572_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_572_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_572_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_572_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_573_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_573_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_573_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_573_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_573_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_573_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_573_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_573_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_573_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_573_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_573_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_573_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_573_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_573_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_573_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_573_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_573_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_573_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_573_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_573_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_573_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_573_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_573_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_573_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_573_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_573_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_573_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_574_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_574_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_574_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_574_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_574_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_574_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_574_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_574_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_574_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_574_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_574_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_574_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_574_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_574_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_574_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_574_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_574_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_574_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_574_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_574_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_574_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_574_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_574_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_574_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_574_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_574_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_574_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_574_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_574_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_574_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_574_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_574_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_575_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_575_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_575_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_575_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_575_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_575_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_575_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_575_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_575_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_575_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_575_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_575_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_575_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_575_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_575_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_575_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_575_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_575_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_575_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_575_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_575_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_575_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_575_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_575_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_575_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_575_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_575_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_575_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_575_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_575_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_575_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_575_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_575_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_575_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_575_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_575_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_575_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_575_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_575_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_575_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_575_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_576_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_576_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_576_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_576_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_576_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_576_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_576_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_576_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_576_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_576_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_576_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_576_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_576_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_576_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_576_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_576_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_576_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_576_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_576_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_576_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_576_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_576_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_576_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_576_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_576_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_576_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_576_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_576_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_576_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_576_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_576_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_576_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_577_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_577_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_577_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_577_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_577_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_577_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_577_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_577_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_577_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_577_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_577_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_577_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_577_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_577_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_577_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_577_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_577_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_577_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_577_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_577_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_577_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_577_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_577_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_577_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_577_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_577_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_577_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_577_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_577_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_577_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_577_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_577_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_578_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_578_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_578_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_578_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_578_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_578_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_578_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_578_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_578_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_578_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_578_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_578_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_578_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_578_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_578_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_578_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_578_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_578_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_578_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_578_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_578_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_578_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_578_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_578_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_578_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_578_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_578_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_578_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_578_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_578_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_579_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_579_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_579_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_579_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_579_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_579_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_579_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_579_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_579_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_579_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_579_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_579_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_579_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_579_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_579_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_579_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_579_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_579_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_579_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_579_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_579_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_579_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_579_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_579_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_579_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_579_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_579_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_579_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_579_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_579_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_579_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_579_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_579_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_579_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_579_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_579_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_579_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_579_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_579_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_57_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_580_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_580_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_580_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_580_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_580_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_580_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_580_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_580_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_580_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_580_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_580_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_580_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_580_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_580_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_580_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_580_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_580_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_580_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_580_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_580_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_580_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_580_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_580_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_580_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_580_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_580_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_580_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_580_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_580_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_580_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_580_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_580_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_580_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_581_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_581_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_581_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_581_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_581_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_581_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_581_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_581_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_581_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_581_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_581_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_581_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_581_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_581_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_581_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_581_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_581_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_581_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_581_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_581_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_581_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_581_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_581_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_581_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_581_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_581_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_581_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_581_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_581_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_581_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_581_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_581_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_581_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_582_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_582_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_582_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_582_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_582_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_582_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_582_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_582_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_582_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_582_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_582_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_582_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_582_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_582_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_582_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_582_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_582_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_582_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_582_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_582_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_582_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_582_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_582_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_582_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_582_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_582_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_582_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_582_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_582_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_582_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_582_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_582_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_582_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_582_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_583_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_583_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_583_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_583_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_583_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_583_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_583_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_583_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_583_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_583_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_583_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_583_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_583_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_583_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_583_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_583_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_583_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_583_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_583_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_583_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_583_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_583_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_583_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_583_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_583_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_583_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_583_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_583_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_583_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_583_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_584_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_584_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_584_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_584_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_584_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_584_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_584_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_584_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_584_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_584_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_584_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_584_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_584_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_584_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_584_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_584_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_584_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_584_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_584_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_584_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_584_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_584_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_584_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_584_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_584_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_585_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_585_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_585_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_585_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_585_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_585_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_585_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_585_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_585_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_585_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_585_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_585_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_585_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_585_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_585_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_585_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_585_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_585_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_585_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_585_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_585_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_585_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_585_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_585_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_585_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_585_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_585_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_585_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_585_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_585_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_585_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_585_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_585_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_585_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_585_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_585_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_586_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_586_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_586_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_586_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_586_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_586_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_586_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_586_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_586_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_586_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_586_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_586_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_586_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_586_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_586_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_586_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_586_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_586_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_586_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_586_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_586_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_586_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_586_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_586_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_586_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_586_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_586_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_586_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_586_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_586_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_586_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_586_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_586_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_586_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_586_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_587_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_587_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_587_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_587_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_587_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_587_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_587_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_587_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_587_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_587_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_587_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_587_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_587_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_587_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_587_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_587_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_587_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_587_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_587_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_587_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_587_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_587_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_587_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_587_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_587_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_587_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_587_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_587_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_587_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_587_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_587_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_587_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_587_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_588_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_588_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_588_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_588_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_588_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_588_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_588_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_588_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_588_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_588_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_588_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_588_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_588_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_588_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_588_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_588_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_588_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_588_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_588_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_588_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_588_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_588_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_588_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_588_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_589_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_589_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_589_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_589_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_589_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_589_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_589_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_589_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_589_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_589_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_589_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_589_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_589_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_589_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_589_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_589_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_589_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_589_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_589_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_589_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_589_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_589_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_589_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_589_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_589_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_589_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_589_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_589_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_589_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_589_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_589_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_58_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_590_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_590_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_590_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_590_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_590_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_590_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_590_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_590_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_590_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_590_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_590_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_590_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_590_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_590_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_590_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_590_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_590_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_590_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_590_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_590_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_590_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_590_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_590_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_590_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_590_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_590_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_590_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_590_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_591_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_591_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_591_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_591_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_591_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_591_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_591_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_591_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_591_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_591_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_591_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_591_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_591_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_591_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_591_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_591_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_591_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_591_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_591_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_591_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_591_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_591_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_591_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_591_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_591_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_591_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_591_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_591_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_591_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_591_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_591_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_591_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_592_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_592_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_592_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_592_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_592_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_592_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_592_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_592_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_592_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_592_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_592_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_592_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_592_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_592_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_592_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_592_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_592_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_592_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_592_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_592_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_592_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_592_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_592_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_592_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_592_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_592_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_592_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_592_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_592_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_592_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_592_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_592_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_593_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_593_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_593_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_593_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_593_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_593_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_593_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_593_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_593_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_593_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_593_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_593_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_593_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_593_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_593_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_593_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_593_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_593_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_593_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_593_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_593_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_593_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_593_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_593_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_593_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_594_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_594_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_594_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_594_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_594_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_594_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_594_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_594_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_594_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_594_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_594_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_594_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_594_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_594_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_594_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_594_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_594_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_594_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_594_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_594_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_595_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_595_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_595_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_595_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_595_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_595_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_595_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_595_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_595_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_595_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_595_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_595_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_595_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_595_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_595_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_595_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_595_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_595_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_595_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_595_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_595_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_595_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_595_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_595_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_595_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_595_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_596_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_596_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_596_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_596_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_596_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_596_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_596_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_596_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_596_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_596_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_596_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_596_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_596_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_596_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_596_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_596_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_596_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_596_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_596_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_596_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_596_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_596_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_596_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_597_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_597_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_597_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_597_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_597_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_597_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_597_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_597_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_597_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_597_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_597_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_597_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_597_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_597_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_597_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_597_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_597_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_597_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_597_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_597_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_597_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_597_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_597_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_597_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_597_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_597_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_597_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_597_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_597_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_598_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_598_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_598_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_598_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_598_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_598_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_598_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_598_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_598_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_598_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_598_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_598_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_598_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_598_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_598_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_598_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_598_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_598_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_598_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_598_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_598_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_598_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_598_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_598_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_598_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_598_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_598_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_598_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_599_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_599_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_599_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_599_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_599_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_599_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_599_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_599_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_599_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_599_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_599_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_599_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_599_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_599_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_599_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_599_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_599_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_599_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_599_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_599_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_599_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_599_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_599_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_599_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_599_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_599_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_599_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_599_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_599_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_599_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_599_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_599_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_599_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_599_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_599_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_599_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_599_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_599_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_599_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_599_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_599_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_599_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_599_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_599_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_599_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_599_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_59_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_59_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_5_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_600_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_600_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_600_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_600_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_600_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_600_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_600_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_600_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_600_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_600_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_600_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_600_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_600_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_600_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_600_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_600_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_600_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_600_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_600_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_600_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_600_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_600_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_600_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_600_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_600_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_600_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_600_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_600_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_600_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_600_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_600_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_601_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_601_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_601_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_601_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_601_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_601_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_601_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_601_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_601_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_601_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_601_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_601_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_601_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_601_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_601_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_601_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_601_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_601_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_601_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_601_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_601_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_601_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_601_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_601_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_601_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_601_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_601_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_601_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_601_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_601_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_601_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_601_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_601_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_601_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_601_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_601_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_601_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_601_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_601_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_601_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_601_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_601_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_602_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_602_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_602_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_602_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_602_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_602_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_602_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_602_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_602_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_602_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_602_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_602_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_602_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_602_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_602_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_602_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_602_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_602_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_602_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_602_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_602_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_602_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_602_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_602_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_602_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_602_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_602_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_602_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_603_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_603_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_603_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_603_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_603_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_603_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_603_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_603_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_603_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_603_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_603_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_603_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_603_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_603_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_603_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_603_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_603_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_603_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_603_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_603_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_603_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_603_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_603_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_603_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_603_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_603_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_603_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_604_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_604_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_604_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_604_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_604_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_604_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_604_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_604_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_604_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_604_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_604_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_604_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_604_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_604_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_604_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_604_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_604_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_604_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_604_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_604_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_605_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_605_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_605_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_605_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_605_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_605_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_605_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_605_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_605_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_605_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_605_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_605_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_605_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_605_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_605_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_605_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_605_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_605_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_605_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_605_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_605_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_605_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_605_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_605_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_605_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_605_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_605_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_605_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_605_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_605_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_605_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_605_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_606_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_606_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_606_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_606_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_606_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_606_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_606_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_606_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_606_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_606_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_606_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_606_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_606_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_606_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_606_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_606_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_606_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_606_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_606_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_606_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_606_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_606_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_606_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_606_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_606_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_606_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_606_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_606_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_606_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_606_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_607_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_607_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_607_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_607_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_607_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_607_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_607_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_607_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_607_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_607_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_607_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_607_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_607_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_607_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_607_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_607_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_607_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_607_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_607_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_607_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_607_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_607_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_607_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_607_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_607_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_607_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_607_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_607_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_607_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_607_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_607_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_607_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_608_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_608_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_608_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_608_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_608_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_608_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_608_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_608_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_608_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_608_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_608_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_608_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_608_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_608_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_608_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_608_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_608_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_608_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_608_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_608_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_608_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_608_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_608_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_608_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_608_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_608_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_608_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_608_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_608_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_608_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_608_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_608_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_608_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_608_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_608_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_608_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_608_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_608_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_608_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_608_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_608_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_609_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_609_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_609_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_609_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_609_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_609_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_609_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_609_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_609_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_609_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_609_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_609_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_609_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_609_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_609_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_609_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_609_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_609_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_609_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_609_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_609_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_609_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_609_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_609_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_609_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_609_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_609_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_609_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_609_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_609_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_609_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_609_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_609_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_609_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_610_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_610_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_610_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_610_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_610_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_610_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_610_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_610_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_610_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_610_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_610_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_610_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_610_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_610_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_610_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_610_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_610_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_610_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_610_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_610_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_610_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_610_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_610_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_610_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_610_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_610_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_610_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_610_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_610_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_610_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_610_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_610_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_610_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_610_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_610_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_610_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_610_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_610_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_611_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_611_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_611_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_611_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_611_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_611_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_611_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_611_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_611_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_611_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_611_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_611_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_611_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_611_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_611_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_611_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_611_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_611_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_611_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_611_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_611_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_611_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_611_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_611_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_611_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_611_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_611_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_611_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_611_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_611_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_611_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_611_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_611_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_612_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_612_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_612_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_612_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_612_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_612_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_612_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_612_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_612_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_612_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_612_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_612_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_612_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_612_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_612_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_612_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_612_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_612_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_612_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_612_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_612_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_612_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_612_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_612_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_612_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_612_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_612_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_612_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_612_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_612_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_612_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_612_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_612_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_612_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_612_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_613_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_613_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_613_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_613_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_613_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_613_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_613_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_613_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_613_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_613_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_613_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_613_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_613_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_613_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_613_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_613_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_613_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_613_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_613_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_613_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_613_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_613_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_614_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_614_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_614_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_614_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_614_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_614_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_614_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_614_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_614_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_614_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_614_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_614_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_614_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_614_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_614_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_614_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_614_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_614_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_614_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_614_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_614_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_614_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_614_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_614_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_614_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_614_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_614_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_614_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_614_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_615_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_615_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_615_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_615_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_615_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_615_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_615_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_615_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_615_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_615_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_615_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_615_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_615_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_615_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_615_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_615_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_615_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_615_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_615_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_615_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_615_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_615_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_615_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_615_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_615_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_615_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_615_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_615_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_615_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_615_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_615_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_615_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_615_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_615_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_616_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_616_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_616_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_616_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_616_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_616_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_616_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_616_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_616_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_616_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_616_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_616_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_616_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_616_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_616_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_616_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_616_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_616_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_616_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_616_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_616_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_616_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_616_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_616_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_616_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_616_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_616_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_616_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_616_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_616_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_616_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_616_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_617_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_617_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_617_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_617_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_617_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_617_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_617_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_617_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_617_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_617_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_617_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_617_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_617_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_617_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_617_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_617_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_617_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_617_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_617_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_617_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_617_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_617_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_617_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_617_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_617_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_617_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_617_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_617_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_617_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_617_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_617_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_617_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_617_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_618_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_618_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_618_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_618_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_618_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_618_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_618_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_618_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_618_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_618_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_618_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_618_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_618_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_618_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_618_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_618_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_618_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_618_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_618_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_618_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_618_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_619_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_619_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_619_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_619_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_619_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_619_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_619_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_619_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_619_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_619_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_619_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_619_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_619_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_619_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_619_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_619_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_619_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_619_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_619_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_619_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_619_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_619_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_619_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_619_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_619_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_620_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_620_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_620_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_620_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_620_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_620_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_620_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_620_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_620_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_620_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_620_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_620_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_620_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_620_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_620_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_620_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_620_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_620_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_620_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_620_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_620_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_620_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_620_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_621_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_621_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_621_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_621_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_621_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_621_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_621_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_621_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_621_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_621_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_621_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_621_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_621_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_621_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_621_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_621_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_621_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_621_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_621_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_621_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_621_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_621_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_621_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_621_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_621_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_621_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_621_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_621_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_622_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_622_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_622_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_622_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_622_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_622_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_622_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_622_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_622_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_622_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_622_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_622_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_622_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_622_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_622_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_622_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_622_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_622_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_622_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_622_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_622_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_622_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_622_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_622_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_622_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_622_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_622_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_622_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_623_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_623_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_623_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_623_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_623_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_623_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_623_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_623_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_623_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_623_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_623_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_623_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_623_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_623_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_623_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_623_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_623_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_623_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_623_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_623_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_624_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_624_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_624_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_624_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_624_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_624_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_624_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_624_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_624_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_624_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_624_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_624_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_624_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_624_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_624_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_624_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_624_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_624_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_624_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_624_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_624_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_624_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_624_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_624_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_624_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_624_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_624_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_624_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_624_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_624_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_624_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_625_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_625_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_625_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_625_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_625_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_625_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_625_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_625_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_625_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_625_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_625_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_625_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_625_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_625_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_625_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_625_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_625_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_625_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_625_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_625_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_625_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_625_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_625_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_625_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_625_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_625_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_626_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_626_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_626_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_626_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_626_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_626_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_626_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_626_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_626_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_626_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_626_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_626_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_626_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_626_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_626_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_626_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_626_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_626_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_626_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_626_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_626_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_626_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_626_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_626_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_626_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_627_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_627_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_627_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_627_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_627_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_627_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_627_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_627_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_627_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_627_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_627_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_627_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_627_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_627_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_627_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_627_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_627_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_627_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_627_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_627_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_627_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_628_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_628_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_628_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_628_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_628_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_628_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_628_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_628_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_628_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_628_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_628_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_628_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_628_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_628_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_628_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_628_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_628_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_628_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_628_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_628_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_628_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_628_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_628_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_628_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_629_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_629_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_629_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_629_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_629_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_629_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_629_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_629_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_629_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_629_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_629_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_629_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_629_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_629_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_629_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_629_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_629_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_629_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_629_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_629_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_629_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_629_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_629_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_629_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_630_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_630_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_630_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_630_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_630_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_630_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_630_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_630_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_630_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_630_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_630_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_630_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_630_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_630_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_630_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_630_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_630_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_630_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_630_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_630_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_630_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_630_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_631_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_631_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_631_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_631_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_631_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_631_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_631_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_631_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_631_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_631_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_631_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_631_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_631_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_631_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_631_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_631_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_631_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_631_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_631_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_631_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_631_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_631_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_631_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_632_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_632_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_632_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_632_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_632_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_632_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_632_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_632_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_632_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_632_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_632_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_632_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_632_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_632_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_632_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_632_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_632_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_632_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_632_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_632_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_632_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_632_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_632_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_632_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_632_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_632_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_633_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_633_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_633_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_633_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_633_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_633_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_633_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_633_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_633_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_633_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_633_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_633_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_633_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_633_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_633_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_633_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_633_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_633_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_633_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_634_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_634_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_634_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_634_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_634_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_634_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_634_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_634_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_634_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_634_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_634_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_634_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_634_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_634_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_634_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_634_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_634_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_634_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_634_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_634_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_634_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_634_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_634_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_634_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_634_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_635_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_635_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_635_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_635_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_635_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_635_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_635_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_635_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_635_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_635_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_635_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_635_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_635_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_635_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_635_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_635_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_635_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_635_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_635_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_635_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_636_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_636_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_636_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_636_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_636_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_636_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_636_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_636_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_636_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_636_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_636_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_636_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_636_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_636_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_636_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_636_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_636_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_636_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_636_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_636_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_636_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_637_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_637_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_637_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_637_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_637_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_637_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_637_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_637_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_637_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_637_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_637_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_637_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_637_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_637_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_637_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_637_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_637_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_637_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_637_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_637_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_638_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_638_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_638_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_638_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_638_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_638_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_638_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_638_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_638_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_638_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_638_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_638_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_638_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_638_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_638_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_638_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_638_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_638_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_638_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_639_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_639_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_639_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_639_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_639_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_639_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_639_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_639_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_639_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_639_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_639_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_639_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_639_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_639_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_639_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_639_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_639_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_639_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_63_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_63_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_640_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_640_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_640_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_640_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_640_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_640_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_640_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_640_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_640_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_640_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_640_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_640_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_640_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_640_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_640_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_640_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_640_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_640_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_641_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_641_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_641_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_641_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_641_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_641_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_641_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_641_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_641_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_641_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_641_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_641_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_641_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_641_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_641_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_641_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_641_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_641_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_642_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_642_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_642_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_642_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_642_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_642_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_642_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_642_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_642_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_642_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_642_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_642_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_642_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_642_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_642_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_642_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_642_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_642_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_643_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_643_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_643_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_643_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_643_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_643_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_643_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_643_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_643_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_643_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_643_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_643_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_643_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_643_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_643_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_643_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_643_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_643_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_644_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_644_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_644_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_644_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_644_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_644_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_644_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_644_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_644_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_644_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_644_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_644_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_644_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_644_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_644_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_644_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_644_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_644_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_645_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_645_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_645_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_645_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_645_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_645_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_645_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_645_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_645_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_645_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_645_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_645_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_645_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_645_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_645_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_645_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_645_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_645_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_646_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_646_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_646_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_646_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_646_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_646_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_646_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_646_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_646_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_646_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_646_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_646_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_646_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_646_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_646_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_646_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_646_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_646_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_647_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_647_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_647_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_647_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_647_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_647_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_647_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_647_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_647_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_647_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_647_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_647_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_647_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_647_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_647_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_647_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_647_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_647_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_648_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_648_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_648_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_648_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_648_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_648_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_648_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_648_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_648_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_648_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_648_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_648_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_648_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_648_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_648_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_648_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_648_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_648_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_649_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_649_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_649_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_649_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_649_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_649_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_649_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_649_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_649_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_649_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_649_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_649_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_649_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_649_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_649_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_649_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_649_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_649_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_64_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_64_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_650_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_650_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_650_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_650_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_650_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_650_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_650_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_650_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_650_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_650_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_650_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_650_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_650_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_650_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_650_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_650_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_650_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_650_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_651_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_651_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_651_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_651_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_651_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_651_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_651_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_651_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_651_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_651_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_651_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_651_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_651_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_651_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_651_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_651_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_651_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_651_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_652_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_652_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_652_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_652_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_652_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_652_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_652_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_652_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_652_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_652_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_652_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_652_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_652_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_652_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_652_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_652_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_652_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_652_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_653_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_653_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_653_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_653_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_653_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_653_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_653_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_653_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_653_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_653_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_653_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_653_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_653_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_653_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_653_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_653_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_653_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_653_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_654_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_654_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_654_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_654_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_654_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_654_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_654_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_654_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_654_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_654_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_654_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_654_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_654_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_654_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_654_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_654_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_654_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_654_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_655_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_655_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_655_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_655_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_655_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_655_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_655_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_655_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_655_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_655_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_655_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_655_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_655_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_655_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_655_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_655_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_655_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_655_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_656_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_656_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_656_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_656_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_656_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_656_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_656_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_656_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_656_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_656_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_656_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_656_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_656_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_656_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_656_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_656_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_656_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_656_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_657_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_657_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_657_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_657_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_657_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_657_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_657_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_657_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_657_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_657_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_657_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_657_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_657_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_657_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_657_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_657_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_657_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_657_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_658_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_658_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_658_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_658_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_658_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_658_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_658_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_658_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_658_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_658_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_658_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_658_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_658_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_658_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_658_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_658_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_658_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_658_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_659_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_659_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_659_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_659_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_659_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_659_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_659_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_659_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_659_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_659_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_659_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_659_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_659_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_659_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_659_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_659_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_659_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_659_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_65_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_65_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_660_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_660_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_660_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_660_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_660_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_660_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_660_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_660_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_660_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_660_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_660_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_660_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_660_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_660_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_660_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_660_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_660_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_660_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_661_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_661_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_661_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_661_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_661_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_661_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_661_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_661_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_661_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_661_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_661_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_661_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_661_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_661_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_661_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_661_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_661_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_661_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_662_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_662_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_662_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_662_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_662_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_662_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_662_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_662_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_662_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_662_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_662_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_662_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_662_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_662_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_662_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_662_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_662_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_662_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_663_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_663_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_663_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_663_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_663_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_663_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_663_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_663_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_663_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_663_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_663_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_663_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_663_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_663_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_663_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_663_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_663_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_663_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_664_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_664_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_664_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_664_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_664_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_664_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_664_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_664_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_664_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_664_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_664_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_664_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_664_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_664_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_664_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_664_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_664_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_664_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_665_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_665_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_665_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_665_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_665_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_665_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_665_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_665_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_665_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_665_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_665_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_665_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_665_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_665_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_665_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_665_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_665_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_665_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_666_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_666_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_666_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_666_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_666_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_666_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_666_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_666_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_666_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_666_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_666_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_666_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_666_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_666_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_666_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_666_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_666_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_666_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_667_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_667_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_667_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_667_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_667_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_667_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_667_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_667_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_667_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_667_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_667_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_667_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_667_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_667_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_667_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_667_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_667_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_667_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_668_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_668_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_668_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_668_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_668_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_668_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_668_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_668_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_668_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_668_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_668_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_668_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_668_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_668_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_668_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_668_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_668_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_668_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_669_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_669_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_669_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_669_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_669_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_669_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_669_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_669_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_669_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_669_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_669_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_669_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_669_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_669_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_669_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_669_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_669_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_669_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_66_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_66_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_670_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_670_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_670_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_670_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_670_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_670_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_670_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_670_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_670_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_670_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_670_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_670_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_670_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_670_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_670_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_670_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_670_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_670_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_671_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_671_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_671_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_671_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_671_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_671_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_671_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_671_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_671_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_671_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_671_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_671_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_671_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_671_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_671_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_671_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_671_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_671_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_672_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_672_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_672_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_672_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_672_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_672_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_672_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_672_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_672_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_672_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_672_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_672_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_672_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_672_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_672_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_672_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_672_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_672_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_673_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_673_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_673_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_673_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_673_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_673_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_673_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_673_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_673_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_673_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_673_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_673_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_673_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_673_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_673_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_673_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_673_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_673_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_674_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_674_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_674_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_674_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_674_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_674_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_674_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_674_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_674_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_674_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_674_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_674_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_674_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_674_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_674_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_674_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_674_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_674_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_675_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_675_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_675_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_675_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_675_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_675_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_675_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_675_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_675_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_675_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_675_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_675_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_675_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_675_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_675_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_675_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_675_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_675_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_676_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_676_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_676_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_676_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_676_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_676_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_676_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_676_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_676_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_676_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_676_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_676_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_676_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_676_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_676_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_676_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_676_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_676_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_676_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_676_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_676_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_676_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_677_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_677_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_677_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_677_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_677_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_677_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_677_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_677_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_677_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_677_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_677_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_677_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_677_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_677_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_677_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_677_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_677_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_677_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_677_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_677_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_677_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_677_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_677_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_677_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_678_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_678_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_678_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_678_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_678_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_678_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_678_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_678_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_678_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_678_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_678_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_678_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_678_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_678_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_678_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_678_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_678_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_678_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_678_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_678_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_678_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_678_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_678_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_678_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_678_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_678_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_678_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_678_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_678_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_679_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_679_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_679_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_679_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_679_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_679_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_679_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_679_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_679_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_679_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_679_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_679_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_679_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_679_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_679_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_679_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_679_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_679_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_679_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_679_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_679_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_679_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_679_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_679_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_679_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_67_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_67_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_67_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_67_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_67_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_67_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_680_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_680_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_680_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_680_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_680_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_680_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_680_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_680_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_680_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_680_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_680_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_680_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_680_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_680_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_680_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_680_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_680_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_680_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_680_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_680_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_680_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_680_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_680_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_680_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_680_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_680_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_680_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_680_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_680_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_680_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_680_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_680_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_680_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_680_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_680_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_680_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_680_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_680_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_680_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_680_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_680_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_680_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_680_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_680_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_680_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_680_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_680_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_680_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_680_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_680_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_680_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_680_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_680_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_680_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_680_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_680_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_680_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_680_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_680_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_680_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_680_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_680_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_680_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_680_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_680_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_680_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_680_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_680_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_680_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_680_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_680_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_680_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_680_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_680_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_680_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_680_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_680_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_680_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_680_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_680_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_680_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_680_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_680_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_680_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_680_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_680_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_680_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_68_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_68_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_68_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_68_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_68_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_69_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_69_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_69_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_69_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_69_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_69_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_70_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_70_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_70_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_70_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_70_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_71_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_71_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_71_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_71_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_71_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_71_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_71_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_72_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_72_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_72_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_72_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_72_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_73_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_73_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_73_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_73_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_73_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_73_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_73_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_74_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_74_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_74_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_74_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_74_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_74_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_74_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_75_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_75_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_75_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_75_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_75_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_75_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_75_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_75_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_76_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_76_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_76_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_76_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_76_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_76_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_76_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_77_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_77_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_78_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_78_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_78_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_78_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_78_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_78_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_79_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_79_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_79_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_79_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_79_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_79_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_7_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_80_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_80_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_80_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_81_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_81_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_81_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_81_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_81_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_82_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_82_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_82_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_82_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_82_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_82_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_83_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_83_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_83_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_83_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_83_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_83_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_83_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_83_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_84_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_84_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_84_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_84_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_84_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_84_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_84_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_85_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_85_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_85_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_85_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_85_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_85_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_85_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_86_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_86_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_86_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_86_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_86_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_86_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_87_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_87_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_87_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_87_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_87_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_87_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_87_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_87_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_88_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_88_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_88_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_88_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_88_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_89_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_89_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_89_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_89_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_89_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_90_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_90_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_90_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_90_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_90_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_91_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_91_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_91_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_91_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_92_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_92_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_92_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_92_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_92_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_92_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_93_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_93_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_93_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_93_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_93_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_93_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_94_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_94_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_94_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_94_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_94_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_95_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_95_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_95_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_95_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_95_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_95_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_96_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_96_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_96_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_96_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_96_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_96_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_97_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_97_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_97_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_97_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_97_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_98_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_98_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_98_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_98_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_98_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_98_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_98_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_99_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_99_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_99_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_99_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_99_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_99_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_9_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Left_681 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_100_Left_781 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_100_Right_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_101_Left_782 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_101_Right_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_102_Left_783 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_102_Right_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_103_Left_784 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_103_Right_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_104_Left_785 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_104_Right_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_105_Left_786 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_105_Right_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_106_Left_787 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_106_Right_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_107_Left_788 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_107_Right_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_108_Left_789 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_108_Right_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_109_Left_790 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_109_Right_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Left_691 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_110_Left_791 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_110_Right_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_111_Left_792 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_111_Right_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_112_Left_793 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_112_Right_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_113_Left_794 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_113_Right_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_114_Left_795 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_114_Right_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_115_Left_796 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_115_Right_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_116_Left_797 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_116_Right_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_117_Left_798 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_117_Right_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_118_Left_799 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_118_Right_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_119_Left_800 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_119_Right_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Left_692 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_120_Left_801 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_120_Right_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_121_Left_802 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_121_Right_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_122_Left_803 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_122_Right_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_123_Left_804 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_123_Right_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_124_Left_805 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_124_Right_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_125_Left_806 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_125_Right_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_126_Left_807 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_126_Right_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_127_Left_808 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_127_Right_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_128_Left_809 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_128_Right_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_129_Left_810 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_129_Right_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Left_693 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_130_Left_811 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_130_Right_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_131_Left_812 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_131_Right_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_132_Left_813 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_132_Right_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_133_Left_814 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_133_Right_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_134_Left_815 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_134_Right_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_135_Left_816 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_135_Right_135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_136_Left_817 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_136_Right_136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_137_Left_818 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_137_Right_137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_138_Left_819 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_138_Right_138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_139_Left_820 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_139_Right_139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Left_694 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_140_Left_821 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_140_Right_140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_141_Left_822 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_141_Right_141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_142_Left_823 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_142_Right_142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_143_Left_824 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_143_Right_143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_144_Left_825 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_144_Right_144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_145_Left_826 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_145_Right_145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_146_Left_827 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_146_Right_146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_147_Left_828 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_147_Right_147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_148_Left_829 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_148_Right_148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_149_Left_830 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_149_Right_149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Left_695 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_150_Left_831 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_150_Right_150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_151_Left_832 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_151_Right_151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_152_Left_833 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_152_Right_152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_153_Left_834 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_153_Right_153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_154_Left_835 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_154_Right_154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_155_Left_836 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_155_Right_155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_156_Left_837 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_156_Right_156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_157_Left_838 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_157_Right_157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_158_Left_839 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_158_Right_158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_159_Left_840 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_159_Right_159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Left_696 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_160_Left_841 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_160_Right_160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_161_Left_842 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_161_Right_161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_162_Left_843 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_162_Right_162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_163_Left_844 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_163_Right_163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_164_Left_845 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_164_Right_164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_165_Left_846 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_165_Right_165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_166_Left_847 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_166_Right_166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_167_Left_848 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_167_Right_167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_168_Left_849 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_168_Right_168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_169_Left_850 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_169_Right_169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Left_697 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_170_Left_851 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_170_Right_170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_171_Left_852 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_171_Right_171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_172_Left_853 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_172_Right_172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_173_Left_854 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_173_Right_173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_174_Left_855 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_174_Right_174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_175_Left_856 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_175_Right_175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_176_Left_857 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_176_Right_176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_177_Left_858 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_177_Right_177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_178_Left_859 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_178_Right_178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_179_Left_860 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_179_Right_179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Left_698 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_180_Left_861 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_180_Right_180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_181_Left_862 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_181_Right_181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_182_Left_863 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_182_Right_182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_183_Left_864 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_183_Right_183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_184_Left_865 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_184_Right_184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_185_Left_866 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_185_Right_185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_186_Left_867 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_186_Right_186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_187_Left_868 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_187_Right_187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_188_Left_869 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_188_Right_188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_189_Left_870 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_189_Right_189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Left_699 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_190_Left_871 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_190_Right_190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_191_Left_872 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_191_Right_191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_192_Left_873 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_192_Right_192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_193_Left_874 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_193_Right_193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_194_Left_875 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_194_Right_194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_195_Left_876 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_195_Right_195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_196_Left_877 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_196_Right_196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_197_Left_878 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_197_Right_197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_198_Left_879 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_198_Right_198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_199_Left_880 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_199_Right_199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Left_700 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Left_682 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_200_Left_881 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_200_Right_200 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_201_Left_882 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_201_Right_201 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_202_Left_883 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_202_Right_202 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_203_Left_884 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_203_Right_203 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_204_Left_885 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_204_Right_204 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_205_Left_886 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_205_Right_205 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_206_Left_887 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_206_Right_206 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_207_Left_888 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_207_Right_207 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_208_Left_889 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_208_Right_208 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_209_Left_890 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_209_Right_209 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Left_701 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_210_Left_891 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_210_Right_210 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_211_Left_892 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_211_Right_211 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_212_Left_893 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_212_Right_212 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_213_Left_894 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_213_Right_213 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_214_Left_895 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_214_Right_214 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_215_Left_896 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_215_Right_215 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_216_Left_897 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_216_Right_216 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_217_Left_898 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_217_Right_217 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_218_Left_899 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_218_Right_218 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_219_Left_900 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_219_Right_219 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Left_702 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_220_Left_901 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_220_Right_220 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_221_Left_902 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_221_Right_221 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_222_Left_903 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_222_Right_222 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_223_Left_904 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_223_Right_223 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_224_Left_905 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_224_Right_224 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_225_Left_906 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_225_Right_225 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_226_Left_907 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_226_Right_226 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_227_Left_908 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_227_Right_227 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_228_Left_909 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_228_Right_228 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_229_Left_910 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_229_Right_229 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Left_703 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_230_Left_911 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_230_Right_230 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_231_Left_912 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_231_Right_231 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_232_Left_913 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_232_Right_232 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_233_Left_914 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_233_Right_233 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_234_Left_915 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_234_Right_234 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_235_Left_916 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_235_Right_235 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_236_Left_917 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_236_Right_236 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_237_Left_918 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_237_Right_237 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_238_Left_919 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_238_Right_238 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_239_Left_920 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_239_Right_239 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Left_704 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_240_Left_921 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_240_Right_240 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_241_Left_922 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_241_Right_241 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_242_Left_923 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_242_Right_242 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_243_Left_924 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_243_Right_243 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_244_Left_925 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_244_Right_244 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_245_Left_926 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_245_Right_245 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_246_Left_927 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_246_Right_246 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_247_Left_928 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_247_Right_247 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_248_Left_929 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_248_Right_248 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_249_Left_930 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_249_Right_249 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Left_705 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_250_Left_931 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_250_Right_250 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_251_Left_932 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_251_Right_251 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_252_Left_933 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_252_Right_252 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_253_Left_934 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_253_Right_253 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_254_Left_935 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_254_Right_254 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_255_Left_936 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_255_Right_255 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_256_Left_937 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_256_Right_256 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_257_Left_938 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_257_Right_257 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_258_Left_939 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_258_Right_258 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_259_Left_940 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_259_Right_259 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Left_706 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_260_Left_941 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_260_Right_260 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_261_Left_942 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_261_Right_261 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_262_Left_943 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_262_Right_262 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_263_Left_944 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_263_Right_263 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_264_Left_945 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_264_Right_264 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_265_Left_946 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_265_Right_265 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_266_Left_947 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_266_Right_266 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_267_Left_948 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_267_Right_267 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_268_Left_949 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_268_Right_268 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_269_Left_950 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_269_Right_269 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Left_707 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Right_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_270_Left_951 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_270_Right_270 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_271_Left_952 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_271_Right_271 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_272_Left_953 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_272_Right_272 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_273_Left_954 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_273_Right_273 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_274_Left_955 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_274_Right_274 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_275_Left_956 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_275_Right_275 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_276_Left_957 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_276_Right_276 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_277_Left_958 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_277_Right_277 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_278_Left_959 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_278_Right_278 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_279_Left_960 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_279_Right_279 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Left_708 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Right_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_280_Left_961 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_280_Right_280 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_281_Left_962 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_281_Right_281 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_282_Left_963 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_282_Right_282 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_283_Left_964 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_283_Right_283 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_284_Left_965 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_284_Right_284 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_285_Left_966 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_285_Right_285 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_286_Left_967 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_286_Right_286 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_287_Left_968 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_287_Right_287 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_288_Left_969 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_288_Right_288 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_289_Left_970 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_289_Right_289 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Left_709 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Right_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_290_Left_971 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_290_Right_290 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_291_Left_972 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_291_Right_291 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_292_Left_973 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_292_Right_292 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_293_Left_974 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_293_Right_293 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_294_Left_975 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_294_Right_294 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_295_Left_976 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_295_Right_295 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_296_Left_977 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_296_Right_296 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_297_Left_978 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_297_Right_297 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_298_Left_979 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_298_Right_298 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_299_Left_980 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_299_Right_299 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Left_710 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Right_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Left_683 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_300_Left_981 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_300_Right_300 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_301_Left_982 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_301_Right_301 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_302_Left_983 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_302_Right_302 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_303_Left_984 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_303_Right_303 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_304_Left_985 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_304_Right_304 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_305_Left_986 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_305_Right_305 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_306_Left_987 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_306_Right_306 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_307_Left_988 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_307_Right_307 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_308_Left_989 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_308_Right_308 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_309_Left_990 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_309_Right_309 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Left_711 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Right_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_310_Left_991 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_310_Right_310 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_311_Left_992 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_311_Right_311 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_312_Left_993 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_312_Right_312 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_313_Left_994 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_313_Right_313 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_314_Left_995 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_314_Right_314 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_315_Left_996 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_315_Right_315 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_316_Left_997 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_316_Right_316 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_317_Left_998 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_317_Right_317 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_318_Left_999 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_318_Right_318 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_319_Left_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_319_Right_319 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Left_712 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Right_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_320_Left_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_320_Right_320 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_321_Left_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_321_Right_321 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_322_Left_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_322_Right_322 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_323_Left_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_323_Right_323 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_324_Left_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_324_Right_324 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_325_Left_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_325_Right_325 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_326_Left_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_326_Right_326 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_327_Left_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_327_Right_327 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_328_Left_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_328_Right_328 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_329_Left_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_329_Right_329 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Left_713 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Right_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_330_Left_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_330_Right_330 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_331_Left_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_331_Right_331 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_332_Left_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_332_Right_332 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_333_Left_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_333_Right_333 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_334_Left_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_334_Right_334 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_335_Left_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_335_Right_335 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_336_Left_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_336_Right_336 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_337_Left_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_337_Right_337 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_338_Left_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_338_Right_338 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_339_Left_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_339_Right_339 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Left_714 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Right_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_340_Left_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_340_Right_340 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_341_Left_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_341_Right_341 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_342_Left_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_342_Right_342 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_343_Left_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_343_Right_343 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_344_Left_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_344_Right_344 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_345_Left_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_345_Right_345 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_346_Left_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_346_Right_346 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_347_Left_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_347_Right_347 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_348_Left_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_348_Right_348 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_349_Left_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_349_Right_349 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Left_715 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Right_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_350_Left_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_350_Right_350 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_351_Left_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_351_Right_351 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_352_Left_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_352_Right_352 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_353_Left_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_353_Right_353 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_354_Left_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_354_Right_354 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_355_Left_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_355_Right_355 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_356_Left_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_356_Right_356 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_357_Left_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_357_Right_357 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_358_Left_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_358_Right_358 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_359_Left_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_359_Right_359 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Left_716 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Right_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_360_Left_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_360_Right_360 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_361_Left_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_361_Right_361 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_362_Left_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_362_Right_362 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_363_Left_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_363_Right_363 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_364_Left_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_364_Right_364 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_365_Left_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_365_Right_365 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_366_Left_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_366_Right_366 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_367_Left_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_367_Right_367 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_368_Left_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_368_Right_368 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_369_Left_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_369_Right_369 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Left_717 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Right_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_370_Left_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_370_Right_370 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_371_Left_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_371_Right_371 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_372_Left_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_372_Right_372 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_373_Left_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_373_Right_373 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_374_Left_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_374_Right_374 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_375_Left_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_375_Right_375 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_376_Left_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_376_Right_376 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_377_Left_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_377_Right_377 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_378_Left_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_378_Right_378 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_379_Left_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_379_Right_379 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Left_718 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Right_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_380_Left_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_380_Right_380 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_381_Left_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_381_Right_381 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_382_Left_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_382_Right_382 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_383_Left_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_383_Right_383 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_384_Left_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_384_Right_384 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_385_Left_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_385_Right_385 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_386_Left_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_386_Right_386 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_387_Left_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_387_Right_387 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_388_Left_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_388_Right_388 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_389_Left_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_389_Right_389 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Left_719 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Right_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_390_Left_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_390_Right_390 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_391_Left_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_391_Right_391 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_392_Left_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_392_Right_392 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_393_Left_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_393_Right_393 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_394_Left_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_394_Right_394 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_395_Left_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_395_Right_395 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_396_Left_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_396_Right_396 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_397_Left_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_397_Right_397 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_398_Left_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_398_Right_398 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_399_Left_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_399_Right_399 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Left_720 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Right_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Left_684 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_400_Left_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_400_Right_400 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_401_Left_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_401_Right_401 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_402_Left_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_402_Right_402 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_403_Left_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_403_Right_403 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_404_Left_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_404_Right_404 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_405_Left_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_405_Right_405 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_406_Left_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_406_Right_406 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_407_Left_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_407_Right_407 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_408_Left_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_408_Right_408 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_409_Left_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_409_Right_409 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Left_721 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Right_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_410_Left_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_410_Right_410 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_411_Left_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_411_Right_411 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_412_Left_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_412_Right_412 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_413_Left_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_413_Right_413 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_414_Left_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_414_Right_414 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_415_Left_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_415_Right_415 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_416_Left_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_416_Right_416 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_417_Left_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_417_Right_417 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_418_Left_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_418_Right_418 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_419_Left_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_419_Right_419 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Left_722 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Right_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_420_Left_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_420_Right_420 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_421_Left_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_421_Right_421 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_422_Left_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_422_Right_422 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_423_Left_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_423_Right_423 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_424_Left_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_424_Right_424 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_425_Left_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_425_Right_425 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_426_Left_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_426_Right_426 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_427_Left_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_427_Right_427 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_428_Left_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_428_Right_428 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_429_Left_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_429_Right_429 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Left_723 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Right_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_430_Left_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_430_Right_430 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_431_Left_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_431_Right_431 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_432_Left_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_432_Right_432 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_433_Left_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_433_Right_433 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_434_Left_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_434_Right_434 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_435_Left_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_435_Right_435 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_436_Left_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_436_Right_436 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_437_Left_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_437_Right_437 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_438_Left_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_438_Right_438 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_439_Left_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_439_Right_439 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Left_724 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Right_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_440_Left_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_440_Right_440 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_441_Left_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_441_Right_441 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_442_Left_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_442_Right_442 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_443_Left_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_443_Right_443 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_444_Left_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_444_Right_444 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_445_Left_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_445_Right_445 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_446_Left_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_446_Right_446 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_447_Left_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_447_Right_447 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_448_Left_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_448_Right_448 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_449_Left_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_449_Right_449 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Left_725 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Right_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_450_Left_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_450_Right_450 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_451_Left_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_451_Right_451 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_452_Left_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_452_Right_452 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_453_Left_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_453_Right_453 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_454_Left_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_454_Right_454 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_455_Left_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_455_Right_455 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_456_Left_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_456_Right_456 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_457_Left_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_457_Right_457 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_458_Left_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_458_Right_458 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_459_Left_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_459_Right_459 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Left_726 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Right_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_460_Left_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_460_Right_460 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_461_Left_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_461_Right_461 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_462_Left_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_462_Right_462 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_463_Left_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_463_Right_463 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_464_Left_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_464_Right_464 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_465_Left_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_465_Right_465 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_466_Left_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_466_Right_466 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_467_Left_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_467_Right_467 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_468_Left_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_468_Right_468 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_469_Left_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_469_Right_469 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Left_727 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Right_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_470_Left_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_470_Right_470 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_471_Left_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_471_Right_471 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_472_Left_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_472_Right_472 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_473_Left_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_473_Right_473 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_474_Left_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_474_Right_474 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_475_Left_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_475_Right_475 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_476_Left_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_476_Right_476 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_477_Left_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_477_Right_477 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_478_Left_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_478_Right_478 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_479_Left_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_479_Right_479 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_Left_728 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_Right_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_480_Left_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_480_Right_480 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_481_Left_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_481_Right_481 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_482_Left_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_482_Right_482 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_483_Left_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_483_Right_483 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_484_Left_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_484_Right_484 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_485_Left_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_485_Right_485 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_486_Left_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_486_Right_486 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_487_Left_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_487_Right_487 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_488_Left_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_488_Right_488 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_489_Left_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_489_Right_489 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_Left_729 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_Right_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_490_Left_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_490_Right_490 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_491_Left_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_491_Right_491 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_492_Left_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_492_Right_492 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_493_Left_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_493_Right_493 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_494_Left_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_494_Right_494 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_495_Left_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_495_Right_495 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_496_Left_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_496_Right_496 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_497_Left_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_497_Right_497 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_498_Left_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_498_Right_498 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_499_Left_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_499_Right_499 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_Left_730 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_Right_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Left_685 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_500_Left_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_500_Right_500 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_501_Left_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_501_Right_501 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_502_Left_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_502_Right_502 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_503_Left_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_503_Right_503 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_504_Left_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_504_Right_504 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_505_Left_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_505_Right_505 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_506_Left_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_506_Right_506 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_507_Left_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_507_Right_507 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_508_Left_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_508_Right_508 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_509_Left_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_509_Right_509 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_Left_731 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_Right_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_510_Left_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_510_Right_510 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_511_Left_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_511_Right_511 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_512_Left_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_512_Right_512 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_513_Left_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_513_Right_513 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_514_Left_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_514_Right_514 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_515_Left_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_515_Right_515 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_516_Left_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_516_Right_516 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_517_Left_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_517_Right_517 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_518_Left_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_518_Right_518 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_519_Left_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_519_Right_519 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_Left_732 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_Right_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_520_Left_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_520_Right_520 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_521_Left_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_521_Right_521 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_522_Left_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_522_Right_522 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_523_Left_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_523_Right_523 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_524_Left_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_524_Right_524 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_525_Left_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_525_Right_525 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_526_Left_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_526_Right_526 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_527_Left_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_527_Right_527 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_528_Left_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_528_Right_528 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_529_Left_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_529_Right_529 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_Left_733 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_Right_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_530_Left_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_530_Right_530 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_531_Left_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_531_Right_531 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_532_Left_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_532_Right_532 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_533_Left_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_533_Right_533 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_534_Left_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_534_Right_534 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_535_Left_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_535_Right_535 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_536_Left_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_536_Right_536 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_537_Left_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_537_Right_537 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_538_Left_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_538_Right_538 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_539_Left_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_539_Right_539 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_Left_734 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_Right_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_540_Left_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_540_Right_540 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_541_Left_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_541_Right_541 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_542_Left_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_542_Right_542 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_543_Left_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_543_Right_543 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_544_Left_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_544_Right_544 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_545_Left_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_545_Right_545 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_546_Left_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_546_Right_546 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_547_Left_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_547_Right_547 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_548_Left_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_548_Right_548 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_549_Left_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_549_Right_549 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_Left_735 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_Right_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_550_Left_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_550_Right_550 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_551_Left_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_551_Right_551 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_552_Left_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_552_Right_552 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_553_Left_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_553_Right_553 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_554_Left_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_554_Right_554 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_555_Left_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_555_Right_555 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_556_Left_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_556_Right_556 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_557_Left_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_557_Right_557 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_558_Left_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_558_Right_558 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_559_Left_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_559_Right_559 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_Left_736 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_Right_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_560_Left_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_560_Right_560 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_561_Left_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_561_Right_561 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_562_Left_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_562_Right_562 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_563_Left_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_563_Right_563 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_564_Left_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_564_Right_564 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_565_Left_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_565_Right_565 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_566_Left_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_566_Right_566 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_567_Left_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_567_Right_567 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_568_Left_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_568_Right_568 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_569_Left_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_569_Right_569 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_Left_737 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_Right_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_570_Left_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_570_Right_570 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_571_Left_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_571_Right_571 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_572_Left_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_572_Right_572 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_573_Left_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_573_Right_573 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_574_Left_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_574_Right_574 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_575_Left_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_575_Right_575 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_576_Left_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_576_Right_576 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_577_Left_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_577_Right_577 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_578_Left_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_578_Right_578 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_579_Left_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_579_Right_579 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_Left_738 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_Right_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_580_Left_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_580_Right_580 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_581_Left_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_581_Right_581 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_582_Left_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_582_Right_582 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_583_Left_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_583_Right_583 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_584_Left_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_584_Right_584 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_585_Left_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_585_Right_585 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_586_Left_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_586_Right_586 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_587_Left_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_587_Right_587 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_588_Left_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_588_Right_588 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_589_Left_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_589_Right_589 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_Left_739 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_Right_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_590_Left_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_590_Right_590 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_591_Left_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_591_Right_591 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_592_Left_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_592_Right_592 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_593_Left_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_593_Right_593 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_594_Left_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_594_Right_594 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_595_Left_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_595_Right_595 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_596_Left_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_596_Right_596 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_597_Left_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_597_Right_597 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_598_Left_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_598_Right_598 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_599_Left_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_599_Right_599 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_Left_740 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_Right_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Left_686 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_600_Left_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_600_Right_600 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_601_Left_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_601_Right_601 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_602_Left_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_602_Right_602 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_603_Left_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_603_Right_603 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_604_Left_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_604_Right_604 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_605_Left_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_605_Right_605 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_606_Left_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_606_Right_606 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_607_Left_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_607_Right_607 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_608_Left_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_608_Right_608 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_609_Left_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_609_Right_609 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_Left_741 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_Right_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_610_Left_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_610_Right_610 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_611_Left_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_611_Right_611 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_612_Left_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_612_Right_612 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_613_Left_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_613_Right_613 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_614_Left_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_614_Right_614 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_615_Left_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_615_Right_615 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_616_Left_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_616_Right_616 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_617_Left_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_617_Right_617 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_618_Left_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_618_Right_618 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_619_Left_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_619_Right_619 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_Left_742 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_Right_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_620_Left_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_620_Right_620 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_621_Left_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_621_Right_621 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_622_Left_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_622_Right_622 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_623_Left_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_623_Right_623 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_624_Left_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_624_Right_624 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_625_Left_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_625_Right_625 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_626_Left_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_626_Right_626 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_627_Left_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_627_Right_627 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_628_Left_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_628_Right_628 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_629_Left_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_629_Right_629 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_Left_743 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_Right_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_630_Left_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_630_Right_630 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_631_Left_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_631_Right_631 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_632_Left_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_632_Right_632 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_633_Left_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_633_Right_633 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_634_Left_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_634_Right_634 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_635_Left_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_635_Right_635 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_636_Left_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_636_Right_636 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_637_Left_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_637_Right_637 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_638_Left_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_638_Right_638 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_639_Left_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_639_Right_639 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_Left_744 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_Right_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_640_Left_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_640_Right_640 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_641_Left_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_641_Right_641 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_642_Left_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_642_Right_642 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_643_Left_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_643_Right_643 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_644_Left_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_644_Right_644 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_645_Left_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_645_Right_645 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_646_Left_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_646_Right_646 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_647_Left_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_647_Right_647 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_648_Left_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_648_Right_648 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_649_Left_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_649_Right_649 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_Left_745 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_Right_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_650_Left_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_650_Right_650 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_651_Left_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_651_Right_651 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_652_Left_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_652_Right_652 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_653_Left_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_653_Right_653 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_654_Left_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_654_Right_654 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_655_Left_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_655_Right_655 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_656_Left_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_656_Right_656 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_657_Left_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_657_Right_657 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_658_Left_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_658_Right_658 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_659_Left_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_659_Right_659 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_Left_746 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_Right_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_660_Left_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_660_Right_660 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_661_Left_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_661_Right_661 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_662_Left_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_662_Right_662 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_663_Left_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_663_Right_663 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_664_Left_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_664_Right_664 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_665_Left_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_665_Right_665 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_666_Left_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_666_Right_666 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_667_Left_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_667_Right_667 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_668_Left_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_668_Right_668 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_669_Left_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_669_Right_669 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_Left_747 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_Right_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_670_Left_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_670_Right_670 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_671_Left_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_671_Right_671 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_672_Left_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_672_Right_672 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_673_Left_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_673_Right_673 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_674_Left_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_674_Right_674 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_675_Left_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_675_Right_675 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_676_Left_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_676_Right_676 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_677_Left_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_677_Right_677 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_678_Left_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_678_Right_678 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_679_Left_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_679_Right_679 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_Left_748 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_Right_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_680_Left_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_680_Right_680 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_Left_749 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_Right_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_Left_750 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_Right_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Left_687 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_Left_751 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_Right_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_Left_752 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_Right_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_Left_753 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_Right_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_Left_754 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_Right_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_Left_755 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_Right_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_Left_756 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_Right_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_Left_757 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_Right_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_Left_758 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_Right_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_Left_759 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_Right_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_Left_760 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_Right_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Left_688 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_Left_761 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_Right_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_Left_762 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_Right_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_Left_763 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_Right_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_83_Left_764 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_83_Right_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_84_Left_765 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_84_Right_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_85_Left_766 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_85_Right_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_86_Left_767 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_86_Right_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_87_Left_768 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_87_Right_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_88_Left_769 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_88_Right_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_89_Left_770 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_89_Right_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Left_689 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_90_Left_771 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_90_Right_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_91_Left_772 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_91_Right_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_92_Left_773 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_92_Right_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_93_Left_774 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_93_Right_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_94_Left_775 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_94_Right_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_95_Left_776 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_95_Right_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_96_Left_777 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_96_Right_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_97_Left_778 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_97_Right_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_98_Left_779 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_98_Right_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_99_Left_780 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_99_Right_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Left_690 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_2157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_2158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_2159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_2161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_2162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_2165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_2168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_2169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_2170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_2171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_2173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_2174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_2175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_2176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_2178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_2180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_2181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_2182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_2183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_2184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_2185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_2186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_2187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_2188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_2189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_2190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_2191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_2192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_2193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_2194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_2197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_2204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_2205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_2206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_2208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_2210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_2211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_2213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_2214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_2215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_2218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_2220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_2221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_2222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_2223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_2224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_2225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_2226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_2227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_2228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_2229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_2232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_2233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_2239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_2240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_2241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_2243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_2244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_2245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_2246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_2247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_2248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_2249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_2250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_2251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_2252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_2253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_2254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_2255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_2256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_2257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_2258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_2259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_2260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_2261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_2262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_2263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_2264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_2265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_2268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_2269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_2272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_2275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_2276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_2278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_2279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_2280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_2281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_2282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_2283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_2284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_2285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_2286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_2287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_2288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_2289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_2290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_2291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_2292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_2293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_2294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_2295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_2296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_2297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_2298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_2299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_2300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_2303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_2304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_2307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_2310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_2311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_2313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_2374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_2375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_2378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_2381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_2383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_2384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_2385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_2386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_2387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_2388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_2389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_2390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_2391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_2392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_2393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_2394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_2395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_2396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_2397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_2398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_2399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_2400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_2401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_2402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_2403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_2404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_2405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_2406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_2407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_2410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_2414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_2418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_2419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_2420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_2421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_2422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_2423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_2424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_2425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_2426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_2427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_2428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_2429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_2430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_2431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_2432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_2433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_2434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_2435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_2436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_2437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_2438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_2439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_2440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_2441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_2442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_2445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_2457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_2458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_2459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_2460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_2461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_2462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_2463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_2464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_2465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_2466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_2467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_2468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_2469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_2470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_2471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_2472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_2473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_2474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_2475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_2476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_2477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_2478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_2482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_2485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_2488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_2489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_2490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_2491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_2492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_2493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_2494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_2495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_2497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_2499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_2501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_2503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_2505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_2506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_2507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_2508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_2509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_2510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_2511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_2513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_2517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_2520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_2523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_2524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_2525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_2526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_2529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_2530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_2532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_2533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_2534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_2537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_2539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_2540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_2541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_2542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_2543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_2544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_2545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_2546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_2547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_2548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_2549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_2552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_2553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_2556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_2560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_2561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_2563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_2564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_2565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_2566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_2567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_2568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_2569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_2570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_2571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_2572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_2573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_2574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_2575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_2576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_2577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_2578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_2579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_2580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_2581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_2582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_2583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_2584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_2587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_2588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_2594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_2596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_2597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_2599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_2600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_2601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_2602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_2603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_2604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_2605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_2606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_2607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_2608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_2609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_2610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_2611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_2612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_2613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_2614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_2615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_2616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_2617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_2618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_2619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_2620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_2623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_2631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_2632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_2634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_2635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_2636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_2637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_2638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_2639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_2644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_2646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_2647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_2650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_2652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_2653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_2654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_2655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_2658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_2659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_2665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_2667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_2668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_2670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_2671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_2672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_2673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_2675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_2676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_2678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_2679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_2680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_2681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_2682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_2683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_2684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_2686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_2687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_2688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_2689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_2690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_2691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_2694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_2695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_2698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_2701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_2702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_2703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_2704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_2705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_2707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_2708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_2709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_2711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_2712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_2714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_2715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_2716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_2717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_2718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_2719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_2720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_2721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_2722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_2723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_2724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_2725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_2726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_2729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_2730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_2733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_2736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_2737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_2738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_2739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_2740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_183_2742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_183_2743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_183_2744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_183_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_183_2746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_183_2747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_183_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_2749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_2750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_2751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_2752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_2753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_2754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_2755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_2756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_185_2757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_185_2758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_185_2759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_185_2760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_185_2761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_185_2762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_185_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_2765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_2766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_2769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_187_2772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_187_2773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_187_2774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_187_2775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_187_2776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_187_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_187_2778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_2779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_2780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_2782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_2783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_2785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_2786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_189_2787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_189_2788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_189_2789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_189_2790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_189_2791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_189_2792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_189_2793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_2794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_2795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_2796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_2797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_2800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_2801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_191_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_191_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_191_2804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_191_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_191_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_191_2807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_191_2808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_2809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_2810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_2811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_2813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_2814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_193_2817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_193_2818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_193_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_193_2820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_193_2821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_193_2822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_193_2823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_2824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_2825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_2826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_2827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_2828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_2829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_2830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_2831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_2832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_2833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_2836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_2837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_196_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_196_2840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_196_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_196_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_196_2843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_196_2844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_196_2845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_196_2846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_197_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_197_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_197_2849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_197_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_197_2851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_197_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_197_2853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_198_2854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_198_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_198_2856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_198_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_198_2858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_198_2859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_198_2860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_198_2861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_199_2862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_199_2863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_199_2864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_199_2865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_199_2866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_199_2867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_199_2868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_200_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_200_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_200_2871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_200_2872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_200_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_200_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_200_2875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_200_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_201_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_201_2878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_201_2879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_201_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_201_2881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_201_2882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_201_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_202_2884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_202_2885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_202_2886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_202_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_202_2888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_202_2889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_202_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_202_2891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_203_2892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_203_2893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_203_2894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_203_2895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_203_2896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_203_2897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_203_2898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_204_2899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_204_2900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_204_2901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_204_2902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_204_2903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_204_2904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_204_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_204_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_205_2907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_205_2908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_205_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_205_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_205_2911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_205_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_205_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_206_2914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_206_2915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_206_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_206_2917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_206_2918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_206_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_206_2920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_206_2921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_207_2922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_207_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_207_2924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_207_2925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_207_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_207_2927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_207_2928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_208_2929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_208_2930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_208_2931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_208_2932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_208_2933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_208_2934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_208_2935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_208_2936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_209_2937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_209_2938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_209_2939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_209_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_209_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_209_2942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_209_2943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_210_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_210_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_210_2946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_210_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_210_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_210_2949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_210_2950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_210_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_211_2952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_211_2953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_211_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_211_2955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_211_2956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_211_2957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_211_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_212_2959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_212_2960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_212_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_212_2962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_212_2963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_212_2964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_212_2965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_212_2966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_213_2967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_213_2968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_213_2969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_213_2970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_213_2971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_213_2972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_213_2973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_214_2974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_214_2975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_214_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_214_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_214_2978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_214_2979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_214_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_214_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_215_2982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_215_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_215_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_215_2985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_215_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_215_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_215_2988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_216_2989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_216_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_216_2991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_216_2992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_216_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_216_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_216_2995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_216_2996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_217_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_217_2998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_217_2999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_217_3000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_217_3001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_217_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_217_3003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_218_3004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_218_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_218_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_218_3007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_218_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_218_3009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_218_3010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_218_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_219_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_219_3013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_219_3014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_219_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_219_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_219_3017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_219_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_220_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_220_3020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_220_3021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_220_3022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_220_3023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_220_3024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_220_3025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_220_3026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_221_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_221_3028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_221_3029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_221_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_221_3031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_221_3032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_221_3033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_222_3034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_222_3035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_222_3036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_222_3037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_222_3038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_222_3039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_222_3040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_222_3041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_223_3042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_223_3043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_223_3044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_223_3045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_223_3046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_223_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_223_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_224_3049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_224_3050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_224_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_224_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_224_3053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_224_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_224_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_224_3056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_225_3057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_225_3058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_225_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_225_3060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_225_3061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_225_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_225_3063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_226_3064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_226_3065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_226_3066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_226_3067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_226_3068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_226_3069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_226_3070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_226_3071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_227_3072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_227_3073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_227_3074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_227_3075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_227_3076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_227_3077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_227_3078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_228_3079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_228_3080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_228_3081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_228_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_228_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_228_3084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_228_3085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_228_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_229_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_229_3088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_229_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_229_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_229_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_229_3092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_229_3093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_230_3094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_230_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_230_3096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_230_3097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_230_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_230_3099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_230_3100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_230_3101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_231_3102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_231_3103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_231_3104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_231_3105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_231_3106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_231_3107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_231_3108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_232_3109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_232_3110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_232_3111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_232_3112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_232_3113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_232_3114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_232_3115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_232_3116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_233_3117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_233_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_233_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_233_3120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_233_3121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_233_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_233_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_234_3124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_234_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_234_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_234_3127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_234_3128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_234_3129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_234_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_234_3131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_235_3132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_235_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_235_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_235_3135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_235_3136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_235_3137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_235_3138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_236_3139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_236_3140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_236_3141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_236_3142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_236_3143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_236_3144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_236_3145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_236_3146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_237_3147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_237_3148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_237_3149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_237_3150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_237_3151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_237_3152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_237_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_238_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_238_3155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_238_3156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_238_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_238_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_238_3159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_238_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_238_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_239_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_239_3163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_239_3164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_239_3165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_239_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_239_3167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_239_3168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_240_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_240_3170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_240_3171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_240_3172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_240_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_240_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_240_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_240_3176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_241_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_241_3178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_241_3179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_241_3180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_241_3181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_241_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_241_3183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_242_3184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_242_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_242_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_242_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_242_3188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_242_3189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_242_3190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_242_3191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_243_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_243_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_243_3194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_243_3195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_243_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_243_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_243_3198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_244_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_244_3200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_244_3201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_244_3202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_244_3203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_244_3204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_244_3205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_244_3206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_245_3207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_245_3208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_245_3209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_245_3210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_245_3211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_245_3212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_245_3213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_246_3214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_246_3215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_246_3216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_246_3217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_246_3218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_246_3219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_246_3220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_246_3221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_247_3222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_247_3223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_247_3224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_247_3225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_247_3226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_247_3227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_247_3228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_248_3229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_248_3230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_248_3231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_248_3232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_248_3233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_248_3234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_248_3235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_248_3236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_249_3237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_249_3238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_249_3239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_249_3240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_249_3241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_249_3242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_249_3243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_250_3244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_250_3245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_250_3246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_250_3247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_250_3248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_250_3249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_250_3250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_250_3251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_251_3252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_251_3253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_251_3254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_251_3255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_251_3256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_251_3257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_251_3258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_252_3259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_252_3260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_252_3261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_252_3262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_252_3263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_252_3264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_252_3265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_252_3266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_253_3267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_253_3268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_253_3269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_253_3270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_253_3271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_253_3272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_253_3273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_254_3274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_254_3275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_254_3276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_254_3277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_254_3278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_254_3279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_254_3280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_254_3281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_255_3282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_255_3283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_255_3284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_255_3285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_255_3286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_255_3287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_255_3288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_256_3289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_256_3290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_256_3291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_256_3292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_256_3293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_256_3294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_256_3295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_256_3296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_257_3297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_257_3298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_257_3299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_257_3300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_257_3301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_257_3302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_257_3303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_258_3304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_258_3305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_258_3306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_258_3307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_258_3308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_258_3309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_258_3310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_258_3311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_259_3312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_259_3313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_259_3314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_259_3315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_259_3316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_259_3317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_259_3318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_260_3319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_260_3320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_260_3321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_260_3322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_260_3323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_260_3324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_260_3325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_260_3326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_261_3327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_261_3328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_261_3329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_261_3330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_261_3331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_261_3332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_261_3333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_262_3334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_262_3335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_262_3336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_262_3337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_262_3338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_262_3339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_262_3340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_262_3341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_263_3342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_263_3343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_263_3344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_263_3345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_263_3346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_263_3347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_263_3348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_264_3349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_264_3350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_264_3351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_264_3352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_264_3353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_264_3354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_264_3355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_264_3356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_265_3357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_265_3358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_265_3359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_265_3360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_265_3361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_265_3362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_265_3363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_266_3364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_266_3365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_266_3366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_266_3367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_266_3368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_266_3369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_266_3370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_266_3371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_267_3372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_267_3373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_267_3374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_267_3375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_267_3376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_267_3377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_267_3378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_268_3379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_268_3380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_268_3381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_268_3382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_268_3383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_268_3384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_268_3385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_268_3386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_269_3387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_269_3388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_269_3389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_269_3390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_269_3391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_269_3392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_269_3393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_270_3394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_270_3395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_270_3396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_270_3397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_270_3398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_270_3399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_270_3400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_270_3401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_271_3402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_271_3403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_271_3404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_271_3405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_271_3406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_271_3407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_271_3408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_272_3409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_272_3410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_272_3411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_272_3412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_272_3413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_272_3414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_272_3415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_272_3416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_273_3417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_273_3418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_273_3419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_273_3420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_273_3421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_273_3422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_273_3423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_274_3424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_274_3425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_274_3426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_274_3427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_274_3428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_274_3429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_274_3430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_274_3431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_275_3432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_275_3433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_275_3434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_275_3435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_275_3436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_275_3437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_275_3438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_276_3439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_276_3440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_276_3441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_276_3442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_276_3443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_276_3444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_276_3445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_276_3446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_277_3447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_277_3448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_277_3449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_277_3450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_277_3451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_277_3452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_277_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_278_3454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_278_3455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_278_3456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_278_3457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_278_3458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_278_3459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_278_3460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_278_3461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_279_3462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_279_3463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_279_3464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_279_3465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_279_3466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_279_3467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_279_3468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_280_3469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_280_3470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_280_3471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_280_3472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_280_3473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_280_3474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_280_3475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_280_3476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_281_3477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_281_3478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_281_3479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_281_3480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_281_3481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_281_3482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_281_3483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_282_3484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_282_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_282_3486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_282_3487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_282_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_282_3489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_282_3490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_282_3491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_283_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_283_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_283_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_283_3495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_283_3496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_283_3497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_283_3498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_284_3499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_284_3500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_284_3501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_284_3502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_284_3503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_284_3504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_284_3505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_284_3506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_285_3507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_285_3508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_285_3509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_285_3510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_285_3511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_285_3512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_285_3513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_286_3514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_286_3515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_286_3516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_286_3517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_286_3518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_286_3519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_286_3520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_286_3521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_287_3522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_287_3523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_287_3524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_287_3525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_287_3526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_287_3527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_287_3528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_288_3529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_288_3530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_288_3531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_288_3532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_288_3533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_288_3534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_288_3535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_288_3536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_289_3537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_289_3538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_289_3539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_289_3540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_289_3541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_289_3542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_289_3543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_290_3544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_290_3545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_290_3546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_290_3547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_290_3548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_290_3549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_290_3550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_290_3551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_291_3552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_291_3553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_291_3554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_291_3555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_291_3556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_291_3557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_291_3558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_292_3559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_292_3560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_292_3561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_292_3562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_292_3563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_292_3564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_292_3565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_292_3566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_293_3567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_293_3568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_293_3569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_293_3570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_293_3571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_293_3572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_293_3573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_294_3574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_294_3575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_294_3576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_294_3577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_294_3578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_294_3579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_294_3580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_294_3581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_295_3582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_295_3583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_295_3584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_295_3585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_295_3586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_295_3587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_295_3588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_296_3589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_296_3590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_296_3591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_296_3592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_296_3593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_296_3594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_296_3595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_296_3596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_297_3597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_297_3598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_297_3599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_297_3600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_297_3601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_297_3602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_297_3603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_298_3604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_298_3605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_298_3606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_298_3607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_298_3608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_298_3609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_298_3610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_298_3611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_299_3612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_299_3613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_299_3614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_299_3615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_299_3616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_299_3617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_299_3618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_300_3619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_300_3620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_300_3621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_300_3622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_300_3623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_300_3624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_300_3625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_300_3626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_301_3627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_301_3628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_301_3629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_301_3630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_301_3631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_301_3632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_301_3633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_302_3634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_302_3635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_302_3636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_302_3637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_302_3638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_302_3639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_302_3640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_302_3641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_303_3642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_303_3643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_303_3644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_303_3645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_303_3646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_303_3647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_303_3648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_304_3649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_304_3650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_304_3651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_304_3652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_304_3653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_304_3654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_304_3655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_304_3656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_305_3657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_305_3658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_305_3659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_305_3660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_305_3661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_305_3662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_305_3663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_306_3664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_306_3665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_306_3666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_306_3667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_306_3668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_306_3669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_306_3670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_306_3671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_307_3672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_307_3673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_307_3674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_307_3675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_307_3676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_307_3677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_307_3678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_308_3679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_308_3680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_308_3681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_308_3682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_308_3683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_308_3684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_308_3685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_308_3686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_309_3687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_309_3688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_309_3689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_309_3690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_309_3691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_309_3692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_309_3693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_310_3694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_310_3695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_310_3696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_310_3697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_310_3698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_310_3699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_310_3700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_310_3701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_311_3702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_311_3703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_311_3704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_311_3705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_311_3706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_311_3707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_311_3708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_312_3709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_312_3710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_312_3711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_312_3712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_312_3713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_312_3714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_312_3715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_312_3716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_313_3717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_313_3718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_313_3719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_313_3720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_313_3721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_313_3722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_313_3723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_314_3724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_314_3725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_314_3726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_314_3727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_314_3728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_314_3729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_314_3730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_314_3731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_315_3732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_315_3733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_315_3734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_315_3735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_315_3736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_315_3737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_315_3738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_316_3739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_316_3740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_316_3741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_316_3742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_316_3743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_316_3744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_316_3745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_316_3746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_317_3747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_317_3748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_317_3749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_317_3750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_317_3751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_317_3752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_317_3753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_318_3754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_318_3755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_318_3756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_318_3757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_318_3758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_318_3759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_318_3760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_318_3761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_319_3762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_319_3763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_319_3764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_319_3765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_319_3766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_319_3767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_319_3768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_320_3769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_320_3770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_320_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_320_3772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_320_3773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_320_3774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_320_3775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_320_3776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_321_3777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_321_3778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_321_3779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_321_3780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_321_3781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_321_3782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_321_3783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_322_3784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_322_3785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_322_3786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_322_3787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_322_3788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_322_3789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_322_3790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_322_3791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_323_3792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_323_3793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_323_3794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_323_3795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_323_3796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_323_3797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_323_3798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_3799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_3800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_3801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_3802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_3804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_3805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_324_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_325_3807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_325_3808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_325_3809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_325_3810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_325_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_325_3812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_325_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_326_3814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_326_3815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_326_3816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_326_3817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_326_3818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_326_3819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_326_3820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_326_3821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_3822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_3823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_3824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_3825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_3826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_3827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_327_3828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_328_3829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_328_3830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_328_3831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_328_3832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_328_3833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_328_3834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_328_3835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_328_3836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_329_3837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_329_3838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_329_3839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_329_3840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_329_3841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_329_3842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_329_3843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_330_3844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_330_3845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_330_3846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_330_3847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_330_3848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_330_3849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_330_3850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_330_3851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_331_3852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_331_3853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_331_3854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_331_3855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_331_3856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_331_3857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_331_3858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_332_3859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_332_3860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_332_3861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_332_3862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_332_3863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_332_3864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_332_3865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_332_3866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_333_3867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_333_3868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_333_3869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_333_3870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_333_3871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_333_3872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_333_3873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_334_3874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_334_3875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_334_3876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_334_3877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_334_3878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_334_3879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_334_3880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_334_3881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_335_3882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_335_3883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_335_3884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_335_3885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_335_3886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_335_3887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_335_3888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_336_3889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_336_3890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_336_3891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_336_3892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_336_3893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_336_3894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_336_3895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_336_3896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_337_3897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_337_3898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_337_3899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_337_3900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_337_3901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_337_3902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_337_3903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_338_3904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_338_3905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_338_3906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_338_3907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_338_3908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_338_3909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_338_3910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_338_3911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_339_3912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_339_3913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_339_3914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_339_3915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_339_3916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_339_3917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_339_3918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_340_3919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_340_3920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_340_3921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_340_3922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_340_3923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_340_3924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_340_3925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_340_3926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_341_3927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_341_3928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_341_3929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_341_3930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_341_3931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_341_3932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_341_3933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_342_3934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_342_3935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_342_3936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_342_3937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_342_3938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_342_3939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_342_3940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_342_3941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_343_3942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_343_3943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_343_3944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_343_3945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_343_3946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_343_3947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_343_3948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_344_3949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_344_3950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_344_3951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_344_3952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_344_3953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_344_3954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_344_3955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_344_3956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_345_3957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_345_3958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_345_3959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_345_3960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_345_3961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_345_3962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_345_3963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_346_3964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_346_3965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_346_3966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_346_3967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_346_3968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_346_3969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_346_3970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_346_3971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_347_3972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_347_3973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_347_3974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_347_3975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_347_3976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_347_3977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_347_3978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_348_3979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_348_3980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_348_3981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_348_3982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_348_3983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_348_3984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_348_3985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_348_3986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_349_3987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_349_3988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_349_3989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_349_3990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_349_3991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_349_3992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_349_3993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_350_3994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_350_3995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_350_3996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_350_3997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_350_3998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_350_3999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_350_4000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_350_4001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_351_4002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_351_4003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_351_4004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_351_4005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_351_4006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_351_4007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_351_4008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_352_4009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_352_4010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_352_4011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_352_4012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_352_4013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_352_4014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_352_4015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_352_4016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_353_4017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_353_4018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_353_4019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_353_4020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_353_4021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_353_4022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_353_4023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_354_4024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_354_4025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_354_4026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_354_4027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_354_4028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_354_4029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_354_4030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_354_4031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_355_4032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_355_4033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_355_4034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_355_4035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_355_4036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_355_4037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_355_4038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_356_4039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_356_4040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_356_4041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_356_4042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_356_4043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_356_4044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_356_4045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_356_4046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_357_4047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_357_4048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_357_4049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_357_4050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_357_4051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_357_4052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_357_4053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_358_4054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_358_4055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_358_4056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_358_4057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_358_4058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_358_4059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_358_4060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_358_4061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_359_4062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_359_4063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_359_4064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_359_4065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_359_4066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_359_4067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_359_4068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_360_4069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_360_4070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_360_4071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_360_4072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_360_4073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_360_4074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_360_4075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_360_4076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_361_4077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_361_4078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_361_4079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_361_4080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_361_4081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_361_4082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_361_4083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_362_4084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_362_4085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_362_4086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_362_4087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_362_4088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_362_4089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_362_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_362_4091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_363_4092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_363_4093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_363_4094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_363_4095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_363_4096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_363_4097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_363_4098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_364_4099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_364_4100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_364_4101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_364_4102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_364_4103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_364_4104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_364_4105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_364_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_365_4107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_365_4108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_365_4109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_365_4110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_365_4111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_365_4112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_365_4113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_366_4114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_366_4115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_366_4116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_366_4117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_366_4118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_366_4119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_366_4120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_366_4121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_367_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_367_4123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_367_4124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_367_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_367_4126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_367_4127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_367_4128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_368_4129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_368_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_368_4131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_368_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_368_4133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_368_4134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_368_4135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_368_4136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_369_4137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_369_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_369_4139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_369_4140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_369_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_369_4142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_369_4143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_370_4144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_370_4145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_370_4146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_370_4147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_370_4148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_370_4149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_370_4150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_370_4151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_371_4152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_371_4153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_371_4154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_371_4155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_371_4156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_371_4157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_371_4158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_372_4159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_372_4160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_372_4161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_372_4162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_372_4163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_372_4164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_372_4165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_372_4166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_373_4167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_373_4168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_373_4169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_373_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_373_4171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_373_4172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_373_4173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_374_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_374_4175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_374_4176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_374_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_374_4178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_374_4179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_374_4180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_374_4181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_375_4182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_375_4183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_375_4184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_375_4185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_375_4186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_375_4187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_375_4188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_376_4189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_376_4190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_376_4191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_376_4192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_376_4193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_376_4194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_376_4195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_376_4196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_377_4197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_377_4198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_377_4199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_377_4200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_377_4201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_377_4202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_377_4203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_378_4204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_378_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_378_4206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_378_4207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_378_4208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_378_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_378_4210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_378_4211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_379_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_379_4213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_379_4214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_379_4215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_379_4216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_379_4217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_379_4218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_380_4219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_380_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_380_4221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_380_4222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_380_4223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_380_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_380_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_380_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_381_4227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_381_4228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_381_4229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_381_4230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_381_4231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_381_4232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_381_4233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_382_4234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_382_4235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_382_4236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_382_4237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_382_4238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_382_4239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_382_4240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_382_4241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_383_4242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_383_4243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_383_4244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_383_4245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_383_4246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_383_4247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_383_4248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_384_4249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_384_4250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_384_4251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_384_4252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_384_4253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_384_4254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_384_4255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_384_4256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_385_4257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_385_4258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_385_4259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_385_4260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_385_4261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_385_4262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_385_4263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_386_4264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_386_4265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_386_4266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_386_4267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_386_4268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_386_4269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_386_4270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_386_4271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_387_4272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_387_4273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_387_4274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_387_4275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_387_4276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_387_4277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_387_4278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_388_4279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_388_4280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_388_4281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_388_4282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_388_4283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_388_4284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_388_4285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_388_4286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_389_4287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_389_4288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_389_4289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_389_4290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_389_4291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_389_4292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_389_4293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_390_4294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_390_4295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_390_4296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_390_4297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_390_4298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_390_4299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_390_4300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_390_4301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_391_4302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_391_4303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_391_4304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_391_4305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_391_4306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_391_4307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_391_4308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_392_4309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_392_4310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_392_4311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_392_4312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_392_4313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_392_4314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_392_4315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_392_4316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_393_4317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_393_4318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_393_4319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_393_4320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_393_4321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_393_4322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_393_4323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_394_4324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_394_4325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_394_4326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_394_4327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_394_4328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_394_4329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_394_4330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_394_4331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_395_4332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_395_4333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_395_4334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_395_4335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_395_4336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_395_4337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_395_4338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_396_4339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_396_4340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_396_4341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_396_4342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_396_4343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_396_4344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_396_4345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_396_4346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_397_4347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_397_4348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_397_4349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_397_4350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_397_4351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_397_4352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_397_4353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_398_4354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_398_4355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_398_4356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_398_4357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_398_4358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_398_4359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_398_4360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_398_4361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_399_4362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_399_4363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_399_4364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_399_4365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_399_4366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_399_4367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_399_4368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_400_4369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_400_4370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_400_4371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_400_4372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_400_4373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_400_4374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_400_4375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_400_4376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_401_4377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_401_4378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_401_4379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_401_4380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_401_4381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_401_4382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_401_4383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_402_4384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_402_4385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_402_4386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_402_4387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_402_4388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_402_4389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_402_4390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_402_4391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_403_4392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_403_4393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_403_4394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_403_4395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_403_4396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_403_4397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_403_4398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_404_4399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_404_4400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_404_4401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_404_4402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_404_4403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_404_4404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_404_4405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_404_4406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_405_4407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_405_4408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_405_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_405_4410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_405_4411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_405_4412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_405_4413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_406_4414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_406_4415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_406_4416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_406_4417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_406_4418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_406_4419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_406_4420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_406_4421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_407_4422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_407_4423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_407_4424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_407_4425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_407_4426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_407_4427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_407_4428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_408_4429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_408_4430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_408_4431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_408_4432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_408_4433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_408_4434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_408_4435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_408_4436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_409_4437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_409_4438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_409_4439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_409_4440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_409_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_409_4442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_409_4443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_410_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_410_4445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_410_4446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_410_4447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_410_4448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_410_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_410_4450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_410_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_411_4452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_411_4453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_411_4454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_411_4455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_411_4456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_411_4457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_411_4458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_412_4459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_412_4460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_412_4461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_412_4462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_412_4463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_412_4464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_412_4465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_412_4466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_413_4467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_413_4468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_413_4469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_413_4470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_413_4471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_413_4472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_413_4473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_414_4474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_414_4475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_414_4476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_414_4477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_414_4478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_414_4479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_414_4480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_414_4481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_415_4482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_415_4483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_415_4484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_415_4485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_415_4486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_415_4487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_415_4488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_416_4489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_416_4490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_416_4491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_416_4492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_416_4493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_416_4494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_416_4495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_416_4496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_417_4497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_417_4498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_417_4499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_417_4500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_417_4501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_417_4502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_417_4503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_418_4504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_418_4505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_418_4506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_418_4507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_418_4508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_418_4509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_418_4510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_418_4511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_419_4512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_419_4513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_419_4514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_419_4515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_419_4516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_419_4517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_419_4518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_420_4519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_420_4520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_420_4521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_420_4522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_420_4523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_420_4524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_420_4525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_420_4526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_421_4527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_421_4528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_421_4529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_421_4530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_421_4531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_421_4532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_421_4533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_422_4534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_422_4535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_422_4536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_422_4537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_422_4538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_422_4539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_422_4540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_422_4541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_423_4542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_423_4543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_423_4544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_423_4545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_423_4546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_423_4547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_423_4548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_424_4549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_424_4550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_424_4551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_424_4552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_424_4553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_424_4554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_424_4555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_424_4556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_425_4557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_425_4558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_425_4559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_425_4560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_425_4561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_425_4562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_425_4563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_426_4564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_426_4565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_426_4566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_426_4567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_426_4568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_426_4569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_426_4570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_426_4571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_427_4572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_427_4573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_427_4574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_427_4575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_427_4576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_427_4577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_427_4578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_428_4579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_428_4580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_428_4581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_428_4582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_428_4583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_428_4584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_428_4585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_428_4586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_429_4587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_429_4588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_429_4589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_429_4590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_429_4591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_429_4592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_429_4593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_430_4594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_430_4595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_430_4596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_430_4597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_430_4598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_430_4599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_430_4600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_430_4601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_431_4602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_431_4603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_431_4604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_431_4605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_431_4606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_431_4607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_431_4608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_432_4609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_432_4610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_432_4611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_432_4612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_432_4613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_432_4614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_432_4615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_432_4616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_433_4617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_433_4618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_433_4619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_433_4620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_433_4621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_433_4622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_433_4623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_434_4624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_434_4625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_434_4626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_434_4627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_434_4628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_434_4629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_434_4630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_434_4631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_435_4632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_435_4633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_435_4634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_435_4635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_435_4636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_435_4637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_435_4638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_436_4639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_436_4640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_436_4641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_436_4642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_436_4643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_436_4644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_436_4645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_436_4646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_437_4647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_437_4648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_437_4649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_437_4650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_437_4651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_437_4652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_437_4653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_438_4654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_438_4655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_438_4656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_438_4657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_438_4658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_438_4659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_438_4660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_438_4661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_439_4662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_439_4663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_439_4664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_439_4665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_439_4666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_439_4667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_439_4668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_440_4669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_440_4670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_440_4671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_440_4672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_440_4673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_440_4674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_440_4675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_440_4676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_441_4677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_441_4678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_441_4679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_441_4680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_441_4681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_441_4682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_441_4683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_442_4684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_442_4685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_442_4686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_442_4687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_442_4688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_442_4689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_442_4690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_442_4691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_443_4692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_443_4693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_443_4694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_443_4695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_443_4696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_443_4697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_443_4698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_444_4699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_444_4700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_444_4701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_444_4702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_444_4703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_444_4704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_444_4705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_444_4706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_445_4707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_445_4708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_445_4709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_445_4710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_445_4711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_445_4712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_445_4713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_446_4714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_446_4715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_446_4716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_446_4717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_446_4718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_446_4719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_446_4720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_446_4721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_447_4722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_447_4723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_447_4724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_447_4725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_447_4726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_447_4727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_447_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_448_4729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_448_4730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_448_4731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_448_4732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_448_4733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_448_4734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_448_4735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_448_4736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_449_4737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_449_4738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_449_4739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_449_4740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_449_4741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_449_4742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_449_4743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_450_4744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_450_4745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_450_4746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_450_4747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_450_4748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_450_4749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_450_4750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_450_4751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_451_4752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_451_4753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_451_4754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_451_4755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_451_4756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_451_4757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_451_4758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_452_4759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_452_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_452_4761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_452_4762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_452_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_452_4764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_452_4765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_452_4766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_453_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_453_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_453_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_453_4770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_453_4771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_453_4772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_453_4773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_454_4774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_454_4775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_454_4776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_454_4777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_454_4778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_454_4779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_454_4780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_454_4781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_455_4782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_455_4783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_455_4784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_455_4785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_455_4786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_455_4787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_455_4788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_456_4789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_456_4790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_456_4791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_456_4792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_456_4793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_456_4794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_456_4795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_456_4796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_457_4797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_457_4798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_457_4799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_457_4800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_457_4801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_457_4802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_457_4803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_458_4804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_458_4805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_458_4806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_458_4807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_458_4808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_458_4809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_458_4810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_458_4811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_459_4812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_459_4813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_459_4814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_459_4815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_459_4816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_459_4817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_459_4818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_460_4819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_460_4820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_460_4821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_460_4822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_460_4823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_460_4824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_460_4825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_460_4826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_461_4827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_461_4828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_461_4829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_461_4830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_461_4831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_461_4832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_461_4833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_462_4834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_462_4835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_462_4836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_462_4837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_462_4838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_462_4839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_462_4840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_462_4841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_463_4842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_463_4843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_463_4844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_463_4845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_463_4846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_463_4847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_463_4848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_464_4849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_464_4850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_464_4851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_464_4852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_464_4853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_464_4854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_464_4855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_464_4856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_465_4857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_465_4858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_465_4859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_465_4860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_465_4861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_465_4862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_465_4863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_466_4864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_466_4865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_466_4866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_466_4867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_466_4868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_466_4869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_466_4870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_466_4871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_467_4872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_467_4873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_467_4874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_467_4875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_467_4876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_467_4877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_467_4878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_468_4879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_468_4880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_468_4881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_468_4882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_468_4883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_468_4884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_468_4885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_468_4886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_469_4887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_469_4888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_469_4889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_469_4890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_469_4891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_469_4892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_469_4893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_470_4894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_470_4895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_470_4896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_470_4897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_470_4898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_470_4899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_470_4900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_470_4901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_471_4902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_471_4903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_471_4904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_471_4905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_471_4906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_471_4907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_471_4908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_472_4909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_472_4910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_472_4911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_472_4912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_472_4913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_472_4914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_472_4915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_472_4916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_473_4917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_473_4918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_473_4919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_473_4920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_473_4921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_473_4922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_473_4923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_474_4924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_474_4925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_474_4926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_474_4927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_474_4928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_474_4929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_474_4930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_474_4931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_475_4932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_475_4933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_475_4934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_475_4935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_475_4936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_475_4937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_475_4938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_476_4939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_476_4940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_476_4941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_476_4942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_476_4943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_476_4944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_476_4945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_476_4946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_477_4947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_477_4948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_477_4949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_477_4950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_477_4951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_477_4952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_477_4953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_478_4954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_478_4955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_478_4956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_478_4957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_478_4958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_478_4959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_478_4960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_478_4961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_479_4962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_479_4963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_479_4964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_479_4965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_479_4966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_479_4967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_479_4968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_480_4969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_480_4970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_480_4971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_480_4972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_480_4973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_480_4974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_480_4975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_480_4976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_481_4977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_481_4978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_481_4979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_481_4980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_481_4981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_481_4982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_481_4983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_482_4984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_482_4985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_482_4986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_482_4987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_482_4988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_482_4989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_482_4990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_482_4991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_483_4992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_483_4993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_483_4994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_483_4995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_483_4996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_483_4997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_483_4998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_484_4999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_484_5000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_484_5001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_484_5002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_484_5003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_484_5004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_484_5005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_484_5006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_485_5007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_485_5008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_485_5009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_485_5010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_485_5011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_485_5012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_485_5013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_486_5014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_486_5015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_486_5016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_486_5017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_486_5018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_486_5019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_486_5020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_486_5021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_487_5022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_487_5023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_487_5024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_487_5025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_487_5026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_487_5027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_487_5028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_488_5029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_488_5030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_488_5031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_488_5032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_488_5033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_488_5034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_488_5035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_488_5036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_489_5037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_489_5038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_489_5039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_489_5040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_489_5041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_489_5042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_489_5043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_490_5044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_490_5045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_490_5046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_490_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_490_5048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_490_5049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_490_5050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_490_5051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_491_5052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_491_5053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_491_5054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_491_5055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_491_5056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_491_5057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_491_5058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_492_5059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_492_5060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_492_5061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_492_5062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_492_5063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_492_5064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_492_5065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_492_5066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_493_5067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_493_5068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_493_5069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_493_5070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_493_5071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_493_5072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_493_5073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_494_5074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_494_5075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_494_5076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_494_5077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_494_5078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_494_5079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_494_5080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_494_5081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_495_5082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_495_5083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_495_5084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_495_5085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_495_5086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_495_5087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_495_5088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_496_5089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_496_5090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_496_5091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_496_5092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_496_5093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_496_5094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_496_5095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_496_5096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_497_5097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_497_5098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_497_5099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_497_5100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_497_5101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_497_5102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_497_5103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_498_5104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_498_5105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_498_5106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_498_5107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_498_5108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_498_5109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_498_5110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_498_5111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_499_5112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_499_5113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_499_5114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_499_5115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_499_5116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_499_5117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_499_5118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_500_5119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_500_5120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_500_5121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_500_5122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_500_5123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_500_5124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_500_5125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_500_5126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_501_5127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_501_5128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_501_5129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_501_5130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_501_5131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_501_5132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_501_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_502_5134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_502_5135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_502_5136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_502_5137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_502_5138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_502_5139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_502_5140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_502_5141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_503_5142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_503_5143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_503_5144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_503_5145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_503_5146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_503_5147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_503_5148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_504_5149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_504_5150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_504_5151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_504_5152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_504_5153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_504_5154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_504_5155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_504_5156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_505_5157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_505_5158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_505_5159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_505_5160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_505_5161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_505_5162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_505_5163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_506_5164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_506_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_506_5166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_506_5167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_506_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_506_5169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_506_5170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_506_5171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_507_5172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_507_5173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_507_5174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_507_5175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_507_5176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_507_5177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_507_5178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_508_5179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_508_5180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_508_5181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_508_5182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_508_5183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_508_5184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_508_5185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_508_5186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_509_5187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_509_5188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_509_5189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_509_5190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_509_5191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_509_5192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_509_5193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_510_5194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_510_5195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_510_5196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_510_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_510_5198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_510_5199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_510_5200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_510_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_511_5202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_511_5203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_511_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_511_5205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_511_5206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_511_5207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_511_5208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_512_5209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_512_5210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_512_5211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_512_5212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_512_5213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_512_5214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_512_5215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_512_5216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_513_5217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_513_5218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_513_5219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_513_5220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_513_5221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_513_5222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_513_5223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_514_5224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_514_5225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_514_5226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_514_5227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_514_5228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_514_5229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_514_5230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_514_5231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_515_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_515_5233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_515_5234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_515_5235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_515_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_515_5237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_515_5238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_516_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_516_5240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_516_5241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_516_5242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_516_5243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_516_5244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_516_5245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_516_5246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_517_5247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_517_5248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_517_5249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_517_5250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_517_5251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_517_5252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_517_5253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_518_5254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_518_5255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_518_5256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_518_5257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_518_5258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_518_5259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_518_5260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_518_5261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_519_5262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_519_5263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_519_5264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_519_5265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_519_5266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_519_5267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_519_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_520_5269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_520_5270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_520_5271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_520_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_520_5273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_520_5274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_520_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_520_5276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_521_5277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_521_5278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_521_5279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_521_5280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_521_5281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_521_5282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_521_5283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_522_5284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_522_5285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_522_5286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_522_5287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_522_5288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_522_5289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_522_5290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_522_5291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_523_5292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_523_5293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_523_5294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_523_5295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_523_5296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_523_5297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_523_5298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_524_5299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_524_5300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_524_5301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_524_5302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_524_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_524_5304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_524_5305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_524_5306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_525_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_525_5308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_525_5309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_525_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_525_5311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_525_5312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_525_5313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_526_5314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_526_5315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_526_5316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_526_5317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_526_5318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_526_5319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_526_5320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_526_5321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_527_5322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_527_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_527_5324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_527_5325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_527_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_527_5327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_527_5328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_528_5329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_528_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_528_5331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_528_5332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_528_5333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_528_5334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_528_5335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_528_5336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_529_5337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_529_5338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_529_5339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_529_5340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_529_5341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_529_5342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_529_5343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_530_5344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_530_5345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_530_5346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_530_5347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_530_5348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_530_5349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_530_5350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_530_5351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_531_5352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_531_5353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_531_5354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_531_5355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_531_5356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_531_5357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_531_5358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_532_5359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_532_5360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_532_5361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_532_5362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_532_5363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_532_5364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_532_5365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_532_5366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_533_5367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_533_5368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_533_5369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_533_5370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_533_5371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_533_5372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_533_5373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_534_5374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_534_5375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_534_5376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_534_5377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_534_5378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_534_5379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_534_5380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_534_5381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_535_5382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_535_5383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_535_5384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_535_5385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_535_5386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_535_5387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_535_5388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_536_5389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_536_5390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_536_5391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_536_5392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_536_5393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_536_5394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_536_5395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_536_5396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_537_5397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_537_5398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_537_5399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_537_5400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_537_5401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_537_5402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_537_5403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_538_5404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_538_5405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_538_5406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_538_5407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_538_5408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_538_5409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_538_5410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_538_5411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_539_5412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_539_5413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_539_5414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_539_5415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_539_5416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_539_5417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_539_5418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_540_5419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_540_5420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_540_5421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_540_5422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_540_5423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_540_5424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_540_5425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_540_5426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_541_5427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_541_5428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_541_5429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_541_5430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_541_5431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_541_5432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_541_5433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_542_5434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_542_5435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_542_5436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_542_5437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_542_5438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_542_5439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_542_5440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_542_5441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_543_5442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_543_5443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_543_5444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_543_5445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_543_5446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_543_5447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_543_5448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_544_5449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_544_5450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_544_5451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_544_5452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_544_5453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_544_5454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_544_5455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_544_5456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_545_5457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_545_5458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_545_5459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_545_5460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_545_5461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_545_5462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_545_5463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_546_5464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_546_5465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_546_5466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_546_5467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_546_5468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_546_5469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_546_5470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_546_5471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_547_5472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_547_5473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_547_5474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_547_5475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_547_5476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_547_5477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_547_5478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_548_5479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_548_5480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_548_5481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_548_5482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_548_5483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_548_5484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_548_5485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_548_5486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_549_5487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_549_5488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_549_5489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_549_5490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_549_5491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_549_5492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_549_5493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_550_5494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_550_5495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_550_5496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_550_5497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_550_5498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_550_5499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_550_5500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_550_5501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_551_5502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_551_5503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_551_5504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_551_5505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_551_5506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_551_5507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_551_5508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_552_5509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_552_5510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_552_5511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_552_5512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_552_5513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_552_5514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_552_5515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_552_5516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_553_5517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_553_5518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_553_5519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_553_5520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_553_5521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_553_5522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_553_5523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_554_5524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_554_5525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_554_5526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_554_5527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_554_5528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_554_5529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_554_5530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_554_5531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_555_5532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_555_5533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_555_5534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_555_5535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_555_5536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_555_5537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_555_5538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_556_5539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_556_5540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_556_5541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_556_5542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_556_5543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_556_5544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_556_5545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_556_5546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_557_5547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_557_5548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_557_5549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_557_5550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_557_5551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_557_5552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_557_5553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_558_5554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_558_5555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_558_5556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_558_5557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_558_5558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_558_5559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_558_5560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_558_5561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_559_5562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_559_5563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_559_5564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_559_5565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_559_5566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_559_5567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_559_5568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_560_5569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_560_5570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_560_5571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_560_5572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_560_5573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_560_5574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_560_5575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_560_5576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_561_5577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_561_5578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_561_5579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_561_5580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_561_5581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_561_5582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_561_5583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_562_5584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_562_5585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_562_5586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_562_5587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_562_5588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_562_5589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_562_5590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_562_5591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_563_5592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_563_5593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_563_5594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_563_5595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_563_5596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_563_5597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_563_5598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_564_5599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_564_5600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_564_5601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_564_5602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_564_5603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_564_5604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_564_5605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_564_5606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_565_5607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_565_5608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_565_5609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_565_5610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_565_5611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_565_5612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_565_5613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_566_5614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_566_5615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_566_5616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_566_5617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_566_5618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_566_5619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_566_5620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_566_5621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_567_5622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_567_5623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_567_5624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_567_5625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_567_5626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_567_5627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_567_5628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_568_5629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_568_5630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_568_5631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_568_5632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_568_5633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_568_5634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_568_5635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_568_5636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_569_5637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_569_5638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_569_5639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_569_5640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_569_5641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_569_5642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_569_5643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_570_5644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_570_5645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_570_5646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_570_5647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_570_5648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_570_5649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_570_5650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_570_5651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_571_5652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_571_5653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_571_5654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_571_5655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_571_5656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_571_5657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_571_5658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_572_5659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_572_5660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_572_5661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_572_5662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_572_5663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_572_5664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_572_5665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_572_5666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_573_5667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_573_5668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_573_5669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_573_5670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_573_5671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_573_5672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_573_5673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_574_5674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_574_5675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_574_5676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_574_5677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_574_5678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_574_5679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_574_5680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_574_5681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_575_5682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_575_5683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_575_5684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_575_5685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_575_5686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_575_5687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_575_5688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_576_5689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_576_5690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_576_5691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_576_5692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_576_5693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_576_5694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_576_5695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_576_5696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_577_5697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_577_5698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_577_5699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_577_5700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_577_5701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_577_5702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_577_5703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_578_5704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_578_5705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_578_5706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_578_5707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_578_5708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_578_5709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_578_5710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_578_5711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_579_5712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_579_5713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_579_5714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_579_5715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_579_5716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_579_5717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_579_5718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_580_5719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_580_5720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_580_5721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_580_5722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_580_5723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_580_5724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_580_5725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_580_5726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_581_5727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_581_5728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_581_5729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_581_5730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_581_5731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_581_5732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_581_5733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_582_5734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_582_5735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_582_5736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_582_5737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_582_5738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_582_5739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_582_5740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_582_5741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_583_5742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_583_5743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_583_5744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_583_5745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_583_5746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_583_5747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_583_5748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_584_5749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_584_5750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_584_5751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_584_5752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_584_5753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_584_5754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_584_5755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_584_5756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_585_5757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_585_5758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_585_5759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_585_5760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_585_5761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_585_5762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_585_5763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_586_5764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_586_5765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_586_5766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_586_5767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_586_5768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_586_5769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_586_5770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_586_5771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_587_5772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_587_5773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_587_5774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_587_5775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_587_5776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_587_5777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_587_5778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_588_5779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_588_5780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_588_5781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_588_5782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_588_5783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_588_5784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_588_5785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_588_5786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_589_5787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_589_5788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_589_5789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_589_5790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_589_5791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_589_5792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_589_5793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_590_5794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_590_5795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_590_5796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_590_5797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_590_5798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_590_5799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_590_5800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_590_5801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_591_5802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_591_5803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_591_5804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_591_5805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_591_5806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_591_5807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_591_5808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_592_5809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_592_5810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_592_5811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_592_5812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_592_5813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_592_5814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_592_5815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_592_5816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_593_5817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_593_5818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_593_5819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_593_5820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_593_5821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_593_5822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_593_5823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_594_5824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_594_5825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_594_5826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_594_5827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_594_5828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_594_5829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_594_5830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_594_5831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_595_5832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_595_5833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_595_5834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_595_5835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_595_5836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_595_5837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_595_5838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_596_5839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_596_5840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_596_5841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_596_5842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_596_5843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_596_5844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_596_5845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_596_5846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_597_5847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_597_5848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_597_5849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_597_5850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_597_5851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_597_5852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_597_5853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_598_5854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_598_5855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_598_5856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_598_5857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_598_5858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_598_5859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_598_5860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_598_5861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_599_5862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_599_5863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_599_5864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_599_5865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_599_5866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_599_5867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_599_5868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_600_5869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_600_5870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_600_5871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_600_5872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_600_5873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_600_5874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_600_5875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_600_5876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_601_5877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_601_5878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_601_5879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_601_5880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_601_5881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_601_5882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_601_5883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_602_5884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_602_5885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_602_5886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_602_5887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_602_5888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_602_5889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_602_5890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_602_5891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_603_5892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_603_5893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_603_5894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_603_5895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_603_5896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_603_5897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_603_5898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_604_5899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_604_5900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_604_5901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_604_5902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_604_5903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_604_5904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_604_5905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_604_5906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_605_5907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_605_5908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_605_5909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_605_5910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_605_5911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_605_5912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_605_5913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_606_5914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_606_5915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_606_5916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_606_5917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_606_5918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_606_5919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_606_5920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_606_5921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_607_5922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_607_5923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_607_5924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_607_5925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_607_5926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_607_5927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_607_5928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_608_5929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_608_5930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_608_5931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_608_5932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_608_5933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_608_5934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_608_5935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_608_5936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_609_5937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_609_5938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_609_5939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_609_5940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_609_5941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_609_5942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_609_5943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_610_5944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_610_5945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_610_5946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_610_5947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_610_5948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_610_5949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_610_5950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_610_5951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_611_5952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_611_5953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_611_5954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_611_5955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_611_5956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_611_5957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_611_5958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_612_5959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_612_5960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_612_5961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_612_5962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_612_5963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_612_5964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_612_5965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_612_5966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_613_5967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_613_5968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_613_5969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_613_5970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_613_5971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_613_5972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_613_5973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_614_5974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_614_5975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_614_5976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_614_5977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_614_5978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_614_5979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_614_5980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_614_5981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_615_5982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_615_5983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_615_5984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_615_5985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_615_5986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_615_5987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_615_5988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_616_5989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_616_5990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_616_5991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_616_5992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_616_5993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_616_5994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_616_5995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_616_5996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_617_5997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_617_5998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_617_5999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_617_6000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_617_6001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_617_6002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_617_6003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_618_6004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_618_6005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_618_6006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_618_6007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_618_6008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_618_6009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_618_6010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_618_6011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_619_6012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_619_6013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_619_6014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_619_6015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_619_6016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_619_6017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_619_6018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_620_6019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_620_6020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_620_6021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_620_6022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_620_6023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_620_6024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_620_6025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_620_6026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_621_6027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_621_6028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_621_6029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_621_6030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_621_6031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_621_6032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_621_6033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_622_6034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_622_6035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_622_6036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_622_6037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_622_6038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_622_6039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_622_6040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_622_6041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_623_6042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_623_6043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_623_6044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_623_6045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_623_6046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_623_6047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_623_6048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_624_6049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_624_6050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_624_6051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_624_6052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_624_6053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_624_6054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_624_6055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_624_6056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_625_6057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_625_6058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_625_6059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_625_6060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_625_6061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_625_6062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_625_6063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_626_6064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_626_6065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_626_6066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_626_6067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_626_6068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_626_6069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_626_6070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_626_6071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_627_6072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_627_6073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_627_6074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_627_6075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_627_6076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_627_6077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_627_6078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_628_6079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_628_6080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_628_6081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_628_6082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_628_6083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_628_6084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_628_6085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_628_6086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_629_6087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_629_6088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_629_6089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_629_6090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_629_6091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_629_6092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_629_6093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_630_6094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_630_6095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_630_6096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_630_6097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_630_6098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_630_6099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_630_6100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_630_6101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_631_6102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_631_6103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_631_6104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_631_6105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_631_6106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_631_6107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_631_6108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_632_6109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_632_6110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_632_6111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_632_6112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_632_6113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_632_6114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_632_6115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_632_6116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_633_6117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_633_6118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_633_6119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_633_6120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_633_6121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_633_6122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_633_6123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_634_6124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_634_6125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_634_6126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_634_6127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_634_6128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_634_6129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_634_6130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_634_6131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_635_6132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_635_6133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_635_6134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_635_6135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_635_6136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_635_6137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_635_6138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_636_6139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_636_6140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_636_6141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_636_6142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_636_6143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_636_6144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_636_6145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_636_6146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_637_6147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_637_6148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_637_6149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_637_6150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_637_6151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_637_6152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_637_6153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_638_6154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_638_6155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_638_6156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_638_6157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_638_6158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_638_6159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_638_6160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_638_6161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_639_6162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_639_6163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_639_6164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_639_6165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_639_6166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_639_6167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_639_6168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_640_6169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_640_6170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_640_6171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_640_6172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_640_6173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_640_6174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_640_6175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_640_6176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_641_6177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_641_6178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_641_6179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_641_6180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_641_6181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_641_6182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_641_6183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_642_6184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_642_6185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_642_6186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_642_6187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_642_6188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_642_6189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_642_6190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_642_6191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_643_6192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_643_6193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_643_6194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_643_6195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_643_6196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_643_6197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_643_6198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_644_6199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_644_6200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_644_6201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_644_6202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_644_6203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_644_6204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_644_6205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_644_6206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_645_6207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_645_6208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_645_6209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_645_6210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_645_6211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_645_6212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_645_6213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_646_6214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_646_6215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_646_6216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_646_6217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_646_6218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_646_6219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_646_6220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_646_6221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_647_6222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_647_6223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_647_6224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_647_6225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_647_6226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_647_6227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_647_6228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_648_6229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_648_6230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_648_6231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_648_6232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_648_6233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_648_6234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_648_6235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_648_6236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_649_6237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_649_6238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_649_6239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_649_6240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_649_6241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_649_6242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_649_6243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_650_6244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_650_6245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_650_6246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_650_6247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_650_6248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_650_6249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_650_6250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_650_6251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_651_6252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_651_6253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_651_6254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_651_6255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_651_6256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_651_6257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_651_6258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_652_6259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_652_6260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_652_6261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_652_6262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_652_6263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_652_6264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_652_6265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_652_6266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_653_6267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_653_6268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_653_6269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_653_6270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_653_6271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_653_6272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_653_6273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_654_6274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_654_6275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_654_6276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_654_6277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_654_6278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_654_6279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_654_6280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_654_6281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_655_6282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_655_6283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_655_6284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_655_6285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_655_6286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_655_6287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_655_6288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_656_6289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_656_6290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_656_6291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_656_6292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_656_6293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_656_6294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_656_6295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_656_6296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_657_6297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_657_6298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_657_6299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_657_6300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_657_6301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_657_6302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_657_6303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_658_6304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_658_6305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_658_6306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_658_6307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_658_6308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_658_6309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_658_6310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_658_6311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_659_6312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_659_6313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_659_6314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_659_6315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_659_6316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_659_6317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_659_6318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_660_6319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_660_6320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_660_6321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_660_6322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_660_6323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_660_6324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_660_6325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_660_6326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_661_6327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_661_6328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_661_6329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_661_6330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_661_6331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_661_6332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_661_6333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_662_6334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_662_6335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_662_6336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_662_6337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_662_6338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_662_6339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_662_6340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_662_6341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_663_6342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_663_6343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_663_6344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_663_6345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_663_6346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_663_6347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_663_6348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_664_6349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_664_6350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_664_6351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_664_6352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_664_6353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_664_6354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_664_6355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_664_6356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_665_6357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_665_6358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_665_6359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_665_6360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_665_6361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_665_6362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_665_6363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_666_6364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_666_6365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_666_6366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_666_6367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_666_6368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_666_6369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_666_6370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_666_6371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_667_6372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_667_6373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_667_6374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_667_6375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_667_6376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_667_6377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_667_6378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_668_6379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_668_6380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_668_6381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_668_6382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_668_6383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_668_6384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_668_6385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_668_6386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_669_6387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_669_6388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_669_6389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_669_6390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_669_6391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_669_6392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_669_6393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_670_6394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_670_6395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_670_6396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_670_6397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_670_6398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_670_6399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_670_6400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_670_6401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_671_6402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_671_6403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_671_6404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_671_6405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_671_6406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_671_6407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_671_6408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_672_6409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_672_6410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_672_6411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_672_6412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_672_6413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_672_6414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_672_6415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_672_6416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_673_6417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_673_6418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_673_6419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_673_6420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_673_6421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_673_6422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_673_6423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_674_6424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_674_6425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_674_6426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_674_6427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_674_6428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_674_6429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_674_6430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_674_6431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_675_6432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_675_6433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_675_6434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_675_6435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_675_6436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_675_6437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_675_6438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_676_6439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_676_6440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_676_6441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_676_6442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_676_6443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_676_6444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_676_6445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_676_6446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_677_6447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_677_6448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_677_6449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_677_6450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_677_6451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_677_6452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_677_6453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_678_6454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_678_6455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_678_6456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_678_6457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_678_6458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_678_6459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_678_6460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_678_6461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_679_6462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_679_6463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_679_6464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_679_6465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_679_6466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_679_6467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_679_6468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_680_6469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_680_6470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_680_6471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_680_6472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_680_6473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_680_6474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_680_6475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_680_6476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_680_6477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_680_6478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_680_6479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_680_6480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_680_6481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_680_6482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_680_6483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2335_ (.I(_0216_),
    .Z(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2336_ (.I(_0956_),
    .Z(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2337_ (.I(_0207_),
    .Z(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2338_ (.I(_0958_),
    .Z(_0959_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2339_ (.I(_0151_),
    .Z(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2340_ (.I(_0960_),
    .Z(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2341_ (.A1(net878),
    .A2(_0959_),
    .A3(_0961_),
    .ZN(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2342_ (.A1(_0955_),
    .A2(_0957_),
    .B(_0962_),
    .ZN(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2343_ (.A1(net862),
    .A2(_0952_),
    .B1(_0954_),
    .B2(net785),
    .C(_0963_),
    .ZN(_0964_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2344_ (.I(_0227_),
    .Z(_0965_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2345_ (.I(_0965_),
    .Z(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2346_ (.I(_0231_),
    .Z(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2347_ (.I(_0967_),
    .Z(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _2348_ (.I(net474),
    .ZN(_0969_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2349_ (.I(_0095_),
    .Z(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2350_ (.I(_0970_),
    .Z(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2351_ (.I(_0239_),
    .Z(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2352_ (.I(_0972_),
    .Z(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _2353_ (.I(net831),
    .ZN(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _2354_ (.A1(_0969_),
    .A2(_0971_),
    .A3(_0762_),
    .B1(_0973_),
    .B2(_0974_),
    .ZN(_0975_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2355_ (.A1(net801),
    .A2(_0966_),
    .B1(_0968_),
    .B2(net816),
    .C(_0975_),
    .ZN(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2356_ (.I(_0245_),
    .Z(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _2357_ (.I(_0977_),
    .Z(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2358_ (.I(_0248_),
    .Z(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _2359_ (.I(_0979_),
    .Z(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2360_ (.I(net194),
    .ZN(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2361_ (.I(_0252_),
    .Z(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2362_ (.I(_0982_),
    .Z(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2363_ (.I(_0255_),
    .Z(_0984_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2364_ (.I(_0984_),
    .Z(_0985_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_8 _2365_ (.I(net769),
    .ZN(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _2366_ (.A1(_0981_),
    .A2(_0983_),
    .B1(_0985_),
    .B2(_0986_),
    .ZN(_0987_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _2367_ (.A1(net179),
    .A2(_0978_),
    .B1(_0980_),
    .B2(net888),
    .C(_0987_),
    .ZN(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2368_ (.I(_0261_),
    .Z(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2369_ (.I(_0989_),
    .Z(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2370_ (.I(_0264_),
    .Z(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2371_ (.I(_0991_),
    .Z(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _2372_ (.I(net145),
    .ZN(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2373_ (.I(_0268_),
    .Z(_0994_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _2374_ (.I(_0994_),
    .Z(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2375_ (.I(_0271_),
    .Z(_0996_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _2376_ (.I(_0996_),
    .Z(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2377_ (.I(net611),
    .ZN(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _2378_ (.A1(_0993_),
    .A2(_0995_),
    .B1(_0997_),
    .B2(_0998_),
    .ZN(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2379_ (.A1(net766),
    .A2(_0990_),
    .B1(_0992_),
    .B2(net753),
    .C(_0999_),
    .ZN(_1000_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _2380_ (.A1(net1813),
    .A2(net1811),
    .A3(_0988_),
    .A4(_1000_),
    .ZN(_1001_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2381_ (.I(_0278_),
    .Z(_1002_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2382_ (.I(_1002_),
    .Z(_1003_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2383_ (.I(_0281_),
    .Z(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2384_ (.I(_1004_),
    .Z(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2385_ (.A1(net614),
    .A2(_1003_),
    .B1(_1005_),
    .B2(net629),
    .ZN(_1006_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2386_ (.I(_0285_),
    .Z(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2387_ (.I(_1007_),
    .Z(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2388_ (.I(_0289_),
    .Z(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2389_ (.I(_1009_),
    .Z(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2390_ (.A1(net645),
    .A2(_1008_),
    .B1(_1010_),
    .B2(net536),
    .ZN(_1011_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2391_ (.I(_0294_),
    .Z(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2392_ (.I(_1012_),
    .Z(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2393_ (.I(_0297_),
    .Z(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2394_ (.I(_1014_),
    .Z(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2395_ (.A1(net551),
    .A2(_1013_),
    .B1(_1015_),
    .B2(net568),
    .ZN(_1016_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2396_ (.I(_0301_),
    .Z(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2397_ (.I(_1017_),
    .Z(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2398_ (.I(_0304_),
    .Z(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2399_ (.I(_1019_),
    .Z(_1020_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2400_ (.A1(net412),
    .A2(_1018_),
    .B1(_1020_),
    .B2(net583),
    .ZN(_1021_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _2401_ (.A1(_1006_),
    .A2(_1011_),
    .A3(_1016_),
    .A4(_1021_),
    .ZN(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2402_ (.I(_0309_),
    .Z(_1023_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2403_ (.I(_1023_),
    .Z(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2404_ (.I(_0313_),
    .Z(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2405_ (.I(_1025_),
    .Z(_1026_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2406_ (.A1(net303),
    .A2(_1024_),
    .B1(_1026_),
    .B2(net54),
    .ZN(_1027_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2407_ (.I(_0317_),
    .Z(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _2408_ (.I(_1028_),
    .Z(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2409_ (.I(_0320_),
    .Z(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2410_ (.I(_1030_),
    .Z(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2411_ (.A1(net318),
    .A2(_1029_),
    .B1(_1031_),
    .B2(net70),
    .ZN(_1032_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2412_ (.I(_0324_),
    .Z(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _2413_ (.I(_1033_),
    .Z(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2414_ (.I(_0327_),
    .Z(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _2415_ (.I(_1035_),
    .Z(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2416_ (.A1(net24),
    .A2(_1034_),
    .B1(_1036_),
    .B2(net39),
    .ZN(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2417_ (.I(_0331_),
    .Z(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2418_ (.I(_1038_),
    .Z(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2419_ (.I(_0334_),
    .Z(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _2420_ (.I(_1040_),
    .Z(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2421_ (.A1(net85),
    .A2(_1039_),
    .B1(_1041_),
    .B2(net117),
    .ZN(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _2422_ (.A1(_1027_),
    .A2(_1032_),
    .A3(_1037_),
    .A4(_1042_),
    .ZN(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _2423_ (.A1(_1001_),
    .A2(_1022_),
    .A3(_1043_),
    .ZN(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2424_ (.A1(_0847_),
    .A2(_0849_),
    .B1(_0950_),
    .B2(_1044_),
    .ZN(_2321_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2425_ (.I(net896),
    .ZN(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2426_ (.I(net506),
    .ZN(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2427_ (.A1(_1046_),
    .A2(_0852_),
    .A3(_0853_),
    .ZN(_1047_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2428_ (.A1(net521),
    .A2(_0856_),
    .A3(_0858_),
    .Z(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2429_ (.I(net599),
    .ZN(_1049_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _2430_ (.A1(_1049_),
    .A2(_0862_),
    .A3(_0725_),
    .ZN(_1050_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2431_ (.I(net491),
    .ZN(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _2432_ (.A1(_1051_),
    .A2(_0866_),
    .A3(_0868_),
    .ZN(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _2433_ (.A1(_1047_),
    .A2(_1048_),
    .A3(_1050_),
    .A4(_1052_),
    .ZN(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2434_ (.I(net460),
    .ZN(_1054_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2435_ (.I(net443),
    .ZN(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _2436_ (.A1(_1054_),
    .A2(_0877_),
    .A3(_0878_),
    .B1(_0880_),
    .B2(_1055_),
    .ZN(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2437_ (.A1(net397),
    .A2(_0872_),
    .B1(_0874_),
    .B2(net428),
    .C(_1056_),
    .ZN(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _2438_ (.I(net288),
    .ZN(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2439_ (.I(net382),
    .ZN(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _2440_ (.A1(_1058_),
    .A2(_0736_),
    .A3(_0890_),
    .B1(_0892_),
    .B2(_1059_),
    .ZN(_1060_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2441_ (.A1(net210),
    .A2(_0885_),
    .B1(_0887_),
    .B2(net227),
    .C(_1060_),
    .ZN(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2442_ (.I(net164),
    .ZN(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2443_ (.I(net149),
    .ZN(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _2444_ (.A1(_1062_),
    .A2(_0902_),
    .A3(_0903_),
    .B1(_0905_),
    .B2(_1063_),
    .ZN(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2445_ (.A1(net258),
    .A2(_0897_),
    .B1(_0899_),
    .B2(net242),
    .C(_1064_),
    .ZN(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _2446_ (.A1(_1053_),
    .A2(_1057_),
    .A3(_1061_),
    .A4(_1065_),
    .ZN(_1066_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2447_ (.A1(net467),
    .A2(_0911_),
    .B1(_0913_),
    .B2(net102),
    .ZN(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2448_ (.A1(net661),
    .A2(_0916_),
    .B1(_0918_),
    .B2(net133),
    .ZN(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2449_ (.A1(net724),
    .A2(_0921_),
    .B1(_0923_),
    .B2(net708),
    .ZN(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2450_ (.A1(net677),
    .A2(_0926_),
    .B1(_0928_),
    .B2(net693),
    .ZN(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _2451_ (.A1(_1067_),
    .A2(_1068_),
    .A3(_1069_),
    .A4(_1070_),
    .ZN(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2452_ (.A1(net351),
    .A2(_0932_),
    .B1(_0934_),
    .B2(net739),
    .ZN(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2453_ (.A1(net9),
    .A2(_0937_),
    .B1(_0939_),
    .B2(net311),
    .ZN(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2454_ (.A1(net366),
    .A2(_0942_),
    .B1(_0944_),
    .B2(net273),
    .ZN(_1074_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2455_ (.A1(net336),
    .A2(_0947_),
    .B(_0753_),
    .ZN(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _2456_ (.A1(_1072_),
    .A2(_1073_),
    .A3(_1074_),
    .A4(_1075_),
    .ZN(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _2457_ (.A1(_1066_),
    .A2(_1071_),
    .A3(_1076_),
    .ZN(_1077_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2458_ (.I(net848),
    .ZN(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2459_ (.A1(net879),
    .A2(_0959_),
    .A3(_0961_),
    .ZN(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2460_ (.A1(_1078_),
    .A2(_0957_),
    .B(_1079_),
    .ZN(_1080_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2461_ (.A1(net863),
    .A2(_0952_),
    .B1(_0954_),
    .B2(net786),
    .C(_1080_),
    .ZN(_1081_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _2462_ (.I(net475),
    .ZN(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _2463_ (.I(net832),
    .ZN(_1083_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _2464_ (.A1(_1082_),
    .A2(_0971_),
    .A3(_0762_),
    .B1(_0973_),
    .B2(_1083_),
    .ZN(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2465_ (.A1(net802),
    .A2(_0966_),
    .B1(_0968_),
    .B2(net817),
    .C(_1084_),
    .ZN(_1085_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2466_ (.I(net195),
    .ZN(_1086_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_8 _2467_ (.I(net770),
    .ZN(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _2468_ (.A1(_1086_),
    .A2(_0983_),
    .B1(_0985_),
    .B2(_1087_),
    .ZN(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2469_ (.A1(net180),
    .A2(_0978_),
    .B1(_0980_),
    .B2(net889),
    .C(_1088_),
    .ZN(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _2470_ (.I(net156),
    .ZN(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2471_ (.I(net622),
    .ZN(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _2472_ (.A1(_1090_),
    .A2(_0995_),
    .B1(_0997_),
    .B2(_1091_),
    .ZN(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2473_ (.A1(net777),
    .A2(_0990_),
    .B1(_0992_),
    .B2(net754),
    .C(_1092_),
    .ZN(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _2474_ (.A1(net1809),
    .A2(net1807),
    .A3(_1089_),
    .A4(_1093_),
    .ZN(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2475_ (.A1(net615),
    .A2(_1003_),
    .B1(_1005_),
    .B2(net630),
    .ZN(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2476_ (.A1(net646),
    .A2(_1008_),
    .B1(_1010_),
    .B2(net537),
    .ZN(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2477_ (.A1(net552),
    .A2(_1013_),
    .B1(_1015_),
    .B2(net569),
    .ZN(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2478_ (.A1(net413),
    .A2(_1018_),
    .B1(_1020_),
    .B2(net584),
    .ZN(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _2479_ (.A1(_1095_),
    .A2(_1096_),
    .A3(_1097_),
    .A4(_1098_),
    .ZN(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2480_ (.A1(net304),
    .A2(_1024_),
    .B1(_1026_),
    .B2(net55),
    .ZN(_1100_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2481_ (.A1(net319),
    .A2(_1029_),
    .B1(_1031_),
    .B2(net71),
    .ZN(_1101_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2482_ (.A1(net25),
    .A2(_1034_),
    .B1(_1036_),
    .B2(net40),
    .ZN(_1102_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2483_ (.A1(net86),
    .A2(_1039_),
    .B1(_1041_),
    .B2(net118),
    .ZN(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _2484_ (.A1(_1100_),
    .A2(_1101_),
    .A3(_1102_),
    .A4(_1103_),
    .ZN(_1104_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _2485_ (.A1(_1094_),
    .A2(_1099_),
    .A3(_1104_),
    .ZN(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2486_ (.A1(_1045_),
    .A2(_0849_),
    .B1(_1077_),
    .B2(_1105_),
    .ZN(_2322_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _2487_ (.I(net12),
    .ZN(_1106_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2488_ (.I(net507),
    .ZN(_1107_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2489_ (.A1(_1107_),
    .A2(_0852_),
    .A3(_0853_),
    .ZN(_1108_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2490_ (.A1(net523),
    .A2(_0856_),
    .A3(_0858_),
    .Z(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2491_ (.I(net601),
    .ZN(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2492_ (.I(_0053_),
    .Z(_1111_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _2493_ (.A1(_1110_),
    .A2(_0862_),
    .A3(_1111_),
    .ZN(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2494_ (.I(net492),
    .ZN(_1113_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _2495_ (.A1(_1113_),
    .A2(_0866_),
    .A3(_0868_),
    .ZN(_1114_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _2496_ (.A1(_1108_),
    .A2(_1109_),
    .A3(_1112_),
    .A4(_1114_),
    .ZN(_1115_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2497_ (.I(net461),
    .ZN(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2498_ (.I(net446),
    .ZN(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _2499_ (.A1(_1116_),
    .A2(_0877_),
    .A3(_0878_),
    .B1(_0880_),
    .B2(_1117_),
    .ZN(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2500_ (.A1(net398),
    .A2(_0872_),
    .B1(_0874_),
    .B2(net429),
    .C(_1118_),
    .ZN(_1119_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _2501_ (.I(net290),
    .ZN(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2502_ (.I(_0735_),
    .Z(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2503_ (.I(net383),
    .ZN(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _2504_ (.A1(_1120_),
    .A2(_1121_),
    .A3(_0890_),
    .B1(_0892_),
    .B2(_1122_),
    .ZN(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2505_ (.A1(net212),
    .A2(_0885_),
    .B1(_0887_),
    .B2(net228),
    .C(_1123_),
    .ZN(_1124_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2506_ (.I(net165),
    .ZN(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2507_ (.I(net150),
    .ZN(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _2508_ (.A1(_1125_),
    .A2(_0902_),
    .A3(_0903_),
    .B1(_0905_),
    .B2(_1126_),
    .ZN(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2509_ (.A1(net259),
    .A2(_0897_),
    .B1(_0899_),
    .B2(net243),
    .C(_1127_),
    .ZN(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _2510_ (.A1(_1115_),
    .A2(_1119_),
    .A3(_1124_),
    .A4(_1128_),
    .ZN(_1129_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2511_ (.A1(net478),
    .A2(_0911_),
    .B1(_0913_),
    .B2(net103),
    .ZN(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2512_ (.A1(net662),
    .A2(_0916_),
    .B1(_0918_),
    .B2(net135),
    .ZN(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2513_ (.A1(net725),
    .A2(_0921_),
    .B1(_0923_),
    .B2(net709),
    .ZN(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2514_ (.A1(net679),
    .A2(_0926_),
    .B1(_0928_),
    .B2(net694),
    .ZN(_1133_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _2515_ (.A1(_1130_),
    .A2(_1131_),
    .A3(_1132_),
    .A4(_1133_),
    .ZN(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2516_ (.A1(net352),
    .A2(_0932_),
    .B1(_0934_),
    .B2(net740),
    .ZN(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2517_ (.A1(net10),
    .A2(_0937_),
    .B1(_0939_),
    .B2(net322),
    .ZN(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2518_ (.A1(net368),
    .A2(_0942_),
    .B1(_0944_),
    .B2(net274),
    .ZN(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2519_ (.I(_0012_),
    .Z(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2520_ (.A1(net337),
    .A2(_0947_),
    .B(_1138_),
    .ZN(_1139_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _2521_ (.A1(_1135_),
    .A2(_1136_),
    .A3(_1137_),
    .A4(_1139_),
    .ZN(_1140_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _2522_ (.A1(_1129_),
    .A2(_1134_),
    .A3(_1140_),
    .ZN(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2523_ (.I(net849),
    .ZN(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2524_ (.A1(net880),
    .A2(_0959_),
    .A3(_0961_),
    .ZN(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2525_ (.A1(_1142_),
    .A2(_0957_),
    .B(_1143_),
    .ZN(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2526_ (.A1(net864),
    .A2(_0952_),
    .B1(_0954_),
    .B2(net787),
    .C(_1144_),
    .ZN(_1145_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _2527_ (.I(net476),
    .ZN(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2528_ (.I(_0066_),
    .Z(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2529_ (.I(_1147_),
    .Z(_1148_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _2530_ (.I(net834),
    .ZN(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _2531_ (.A1(_1146_),
    .A2(_0971_),
    .A3(_1148_),
    .B1(_0973_),
    .B2(_1149_),
    .ZN(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2532_ (.A1(net803),
    .A2(_0966_),
    .B1(_0968_),
    .B2(net818),
    .C(_1150_),
    .ZN(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2533_ (.I(net196),
    .ZN(_1152_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_8 _2534_ (.I(net771),
    .ZN(_1153_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _2535_ (.A1(_1152_),
    .A2(_0983_),
    .B1(_0985_),
    .B2(_1153_),
    .ZN(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _2536_ (.A1(net181),
    .A2(_0978_),
    .B1(_0980_),
    .B2(net890),
    .C(_1154_),
    .ZN(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _2537_ (.I(net167),
    .ZN(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2538_ (.I(net633),
    .ZN(_1157_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _2539_ (.A1(_1156_),
    .A2(_0995_),
    .B1(_0997_),
    .B2(_1157_),
    .ZN(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2540_ (.A1(net789),
    .A2(_0990_),
    .B1(_0992_),
    .B2(net756),
    .C(_1158_),
    .ZN(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _2541_ (.A1(net1805),
    .A2(net1803),
    .A3(_1155_),
    .A4(_1159_),
    .ZN(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2542_ (.A1(net616),
    .A2(_1003_),
    .B1(_1005_),
    .B2(net631),
    .ZN(_1161_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2543_ (.A1(net647),
    .A2(_1008_),
    .B1(_1010_),
    .B2(net538),
    .ZN(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2544_ (.A1(net553),
    .A2(_1013_),
    .B1(_1015_),
    .B2(net570),
    .ZN(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2545_ (.A1(net414),
    .A2(_1018_),
    .B1(_1020_),
    .B2(net585),
    .ZN(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _2546_ (.A1(_1161_),
    .A2(_1162_),
    .A3(_1163_),
    .A4(_1164_),
    .ZN(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2547_ (.A1(net305),
    .A2(_1024_),
    .B1(_1026_),
    .B2(net57),
    .ZN(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2548_ (.A1(net320),
    .A2(_1029_),
    .B1(_1031_),
    .B2(net72),
    .ZN(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2549_ (.A1(net26),
    .A2(_1034_),
    .B1(_1036_),
    .B2(net41),
    .ZN(_1168_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2550_ (.A1(net87),
    .A2(_1039_),
    .B1(_1041_),
    .B2(net119),
    .ZN(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _2551_ (.A1(_1166_),
    .A2(_1167_),
    .A3(_1168_),
    .A4(_1169_),
    .ZN(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _2552_ (.A1(_1160_),
    .A2(_1165_),
    .A3(_1170_),
    .ZN(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2553_ (.A1(_1106_),
    .A2(_0849_),
    .B1(_1141_),
    .B2(_1171_),
    .ZN(_2310_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2554_ (.I(net23),
    .ZN(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2555_ (.I(net508),
    .ZN(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2556_ (.A1(_1173_),
    .A2(_0852_),
    .A3(_0853_),
    .ZN(_1174_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2557_ (.A1(net524),
    .A2(_0856_),
    .A3(_0858_),
    .Z(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2558_ (.I(net602),
    .ZN(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _2559_ (.A1(_1176_),
    .A2(_0862_),
    .A3(_1111_),
    .ZN(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2560_ (.I(net493),
    .ZN(_1178_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _2561_ (.A1(_1178_),
    .A2(_0866_),
    .A3(_0868_),
    .ZN(_1179_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _2562_ (.A1(_1174_),
    .A2(_1175_),
    .A3(_1177_),
    .A4(_1179_),
    .ZN(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2563_ (.I(net462),
    .ZN(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2564_ (.I(net447),
    .ZN(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _2565_ (.A1(_1181_),
    .A2(_0877_),
    .A3(_0878_),
    .B1(_0880_),
    .B2(_1182_),
    .ZN(_1183_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2566_ (.A1(net399),
    .A2(_0872_),
    .B1(_0874_),
    .B2(net430),
    .C(_1183_),
    .ZN(_1184_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _2567_ (.I(net291),
    .ZN(_1185_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2568_ (.I(net384),
    .ZN(_1186_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _2569_ (.A1(_1185_),
    .A2(_1121_),
    .A3(_0890_),
    .B1(_0892_),
    .B2(_1186_),
    .ZN(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2570_ (.A1(net213),
    .A2(_0885_),
    .B1(_0887_),
    .B2(net229),
    .C(_1187_),
    .ZN(_1188_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2571_ (.I(net166),
    .ZN(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2572_ (.I(net151),
    .ZN(_1190_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _2573_ (.A1(_1189_),
    .A2(_0902_),
    .A3(_0903_),
    .B1(_0905_),
    .B2(_1190_),
    .ZN(_1191_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2574_ (.A1(net260),
    .A2(_0897_),
    .B1(_0899_),
    .B2(net244),
    .C(_1191_),
    .ZN(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _2575_ (.A1(_1180_),
    .A2(_1184_),
    .A3(_1188_),
    .A4(_1192_),
    .ZN(_1193_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2576_ (.A1(net489),
    .A2(_0911_),
    .B1(_0913_),
    .B2(net104),
    .ZN(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2577_ (.A1(net663),
    .A2(_0916_),
    .B1(_0918_),
    .B2(net136),
    .ZN(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2578_ (.A1(net726),
    .A2(_0921_),
    .B1(_0923_),
    .B2(net710),
    .ZN(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2579_ (.A1(net680),
    .A2(_0926_),
    .B1(_0928_),
    .B2(net695),
    .ZN(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _2580_ (.A1(_1194_),
    .A2(_1195_),
    .A3(_1196_),
    .A4(_1197_),
    .ZN(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2581_ (.A1(net353),
    .A2(_0932_),
    .B1(_0934_),
    .B2(net741),
    .ZN(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2582_ (.A1(net11),
    .A2(_0937_),
    .B1(_0939_),
    .B2(net333),
    .ZN(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2583_ (.A1(net369),
    .A2(_0942_),
    .B1(_0944_),
    .B2(net275),
    .ZN(_1201_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2584_ (.A1(net338),
    .A2(_0947_),
    .B(_1138_),
    .ZN(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _2585_ (.A1(_1199_),
    .A2(_1200_),
    .A3(_1201_),
    .A4(_1202_),
    .ZN(_1203_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _2586_ (.A1(_1193_),
    .A2(_1198_),
    .A3(_1203_),
    .ZN(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2587_ (.I(net850),
    .ZN(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2588_ (.A1(net881),
    .A2(_0959_),
    .A3(_0961_),
    .ZN(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2589_ (.A1(_1205_),
    .A2(_0957_),
    .B(_1206_),
    .ZN(_1207_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2590_ (.A1(net865),
    .A2(_0952_),
    .B1(_0954_),
    .B2(net788),
    .C(_1207_),
    .ZN(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _2591_ (.I(net477),
    .ZN(_1209_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _2592_ (.I(net835),
    .ZN(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _2593_ (.A1(_1209_),
    .A2(_0971_),
    .A3(_1148_),
    .B1(_0973_),
    .B2(_1210_),
    .ZN(_1211_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2594_ (.A1(net804),
    .A2(_0966_),
    .B1(_0968_),
    .B2(net819),
    .C(_1211_),
    .ZN(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2595_ (.I(net197),
    .ZN(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_8 _2596_ (.I(net772),
    .ZN(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _2597_ (.A1(_1213_),
    .A2(_0983_),
    .B1(_0985_),
    .B2(_1214_),
    .ZN(_1215_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2598_ (.A1(net182),
    .A2(_0978_),
    .B1(_0980_),
    .B2(net891),
    .C(_1215_),
    .ZN(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _2599_ (.I(net178),
    .ZN(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2600_ (.I(net644),
    .ZN(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _2601_ (.A1(_1217_),
    .A2(_0995_),
    .B1(_0997_),
    .B2(_1218_),
    .ZN(_1219_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2602_ (.A1(net800),
    .A2(_0990_),
    .B1(_0992_),
    .B2(net757),
    .C(_1219_),
    .ZN(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _2603_ (.A1(net1801),
    .A2(net1799),
    .A3(_1216_),
    .A4(_1220_),
    .ZN(_1221_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2604_ (.A1(net617),
    .A2(_1003_),
    .B1(_1005_),
    .B2(net632),
    .ZN(_1222_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2605_ (.A1(net648),
    .A2(_1008_),
    .B1(_1010_),
    .B2(net539),
    .ZN(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2606_ (.A1(net554),
    .A2(_1013_),
    .B1(_1015_),
    .B2(net571),
    .ZN(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2607_ (.A1(net415),
    .A2(_1018_),
    .B1(_1020_),
    .B2(net586),
    .ZN(_1225_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _2608_ (.A1(_1222_),
    .A2(_1223_),
    .A3(_1224_),
    .A4(_1225_),
    .ZN(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2609_ (.A1(net306),
    .A2(_1024_),
    .B1(_1026_),
    .B2(net58),
    .ZN(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2610_ (.A1(net321),
    .A2(_1029_),
    .B1(_1031_),
    .B2(net73),
    .ZN(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2611_ (.A1(net27),
    .A2(_1034_),
    .B1(_1036_),
    .B2(net42),
    .ZN(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2612_ (.A1(net88),
    .A2(_1039_),
    .B1(_1041_),
    .B2(net120),
    .ZN(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _2613_ (.A1(_1227_),
    .A2(_1228_),
    .A3(_1229_),
    .A4(_1230_),
    .ZN(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _2614_ (.A1(_1221_),
    .A2(_1226_),
    .A3(_1231_),
    .ZN(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2615_ (.A1(_1172_),
    .A2(_0849_),
    .B1(_1204_),
    .B2(_1232_),
    .ZN(_2311_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2616_ (.I(net34),
    .ZN(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2617_ (.I(_0848_),
    .Z(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2618_ (.I(net509),
    .ZN(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2619_ (.I(_0851_),
    .Z(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2620_ (.I(_0531_),
    .Z(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2621_ (.A1(_1235_),
    .A2(_1236_),
    .A3(_1237_),
    .ZN(_1238_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2622_ (.I(_0855_),
    .Z(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2623_ (.I(_0857_),
    .Z(_1240_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2624_ (.A1(net525),
    .A2(_1239_),
    .A3(_1240_),
    .Z(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2625_ (.I(net603),
    .ZN(_1242_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2626_ (.I(_0861_),
    .Z(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _2627_ (.A1(_1242_),
    .A2(_1243_),
    .A3(_1111_),
    .ZN(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2628_ (.I(net494),
    .ZN(_1245_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2629_ (.I(_0865_),
    .Z(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2630_ (.I(_0867_),
    .Z(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2631_ (.A1(_1245_),
    .A2(_1246_),
    .A3(_1247_),
    .ZN(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _2632_ (.A1(_1238_),
    .A2(_1241_),
    .A3(_1244_),
    .A4(_1248_),
    .ZN(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2633_ (.I(_0871_),
    .Z(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2634_ (.I(_0873_),
    .Z(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2635_ (.I(net463),
    .ZN(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2636_ (.I(_0876_),
    .Z(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2637_ (.I(_0079_),
    .Z(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2638_ (.I(_0879_),
    .Z(_1255_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2639_ (.I(net448),
    .ZN(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _2640_ (.A1(_1252_),
    .A2(_1253_),
    .A3(_1254_),
    .B1(_1255_),
    .B2(_1256_),
    .ZN(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2641_ (.A1(net401),
    .A2(_1250_),
    .B1(_1251_),
    .B2(net431),
    .C(_1257_),
    .ZN(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _2642_ (.I(_0884_),
    .Z(_1259_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _2643_ (.I(_0886_),
    .Z(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _2644_ (.I(net292),
    .ZN(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2645_ (.I(_0889_),
    .Z(_1262_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2646_ (.I(_0891_),
    .Z(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2647_ (.I(net385),
    .ZN(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _2648_ (.A1(_1261_),
    .A2(_1121_),
    .A3(_1262_),
    .B1(_1263_),
    .B2(_1264_),
    .ZN(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2649_ (.A1(net214),
    .A2(_1259_),
    .B1(_1260_),
    .B2(net230),
    .C(_1265_),
    .ZN(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _2650_ (.I(_0896_),
    .Z(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _2651_ (.I(_0898_),
    .Z(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2652_ (.I(net168),
    .ZN(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _2653_ (.I(_0901_),
    .Z(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2654_ (.I(_0127_),
    .Z(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2655_ (.I(_0904_),
    .Z(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2656_ (.I(net152),
    .ZN(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _2657_ (.A1(_1269_),
    .A2(_1270_),
    .A3(_1271_),
    .B1(_1272_),
    .B2(_1273_),
    .ZN(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2658_ (.A1(net261),
    .A2(_1267_),
    .B1(_1268_),
    .B2(net246),
    .C(_1274_),
    .ZN(_1275_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _2659_ (.A1(_1249_),
    .A2(_1258_),
    .A3(_1266_),
    .A4(_1275_),
    .ZN(_1276_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2660_ (.I(_0910_),
    .Z(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2661_ (.I(_0912_),
    .Z(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2662_ (.A1(net500),
    .A2(_1277_),
    .B1(_1278_),
    .B2(net105),
    .ZN(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2663_ (.I(_0915_),
    .Z(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2664_ (.I(_0917_),
    .Z(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2665_ (.A1(net664),
    .A2(_1280_),
    .B1(_1281_),
    .B2(net137),
    .ZN(_1282_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2666_ (.I(_0920_),
    .Z(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2667_ (.I(_0922_),
    .Z(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2668_ (.A1(net727),
    .A2(_1283_),
    .B1(_1284_),
    .B2(net712),
    .ZN(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _2669_ (.I(_0925_),
    .Z(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _2670_ (.I(_0927_),
    .Z(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2671_ (.A1(net681),
    .A2(_1286_),
    .B1(_1287_),
    .B2(net696),
    .ZN(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _2672_ (.A1(_1279_),
    .A2(_1282_),
    .A3(_1285_),
    .A4(_1288_),
    .ZN(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _2673_ (.I(_0931_),
    .Z(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _2674_ (.I(_0933_),
    .Z(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2675_ (.A1(net354),
    .A2(_1290_),
    .B1(_1291_),
    .B2(net742),
    .ZN(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _2676_ (.I(_0936_),
    .Z(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _2677_ (.I(_0938_),
    .Z(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2678_ (.A1(net13),
    .A2(_1293_),
    .B1(_1294_),
    .B2(net345),
    .ZN(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2679_ (.I(_0941_),
    .Z(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2680_ (.I(_0943_),
    .Z(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2681_ (.A1(net370),
    .A2(_1296_),
    .B1(_1297_),
    .B2(net276),
    .ZN(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _2682_ (.I(_0946_),
    .Z(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2683_ (.A1(net339),
    .A2(_1299_),
    .B(_1138_),
    .ZN(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _2684_ (.A1(_1292_),
    .A2(_1295_),
    .A3(_1298_),
    .A4(_1300_),
    .ZN(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2685_ (.A1(_1276_),
    .A2(_1289_),
    .A3(_1301_),
    .ZN(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _2686_ (.I(_0951_),
    .Z(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2687_ (.I(_0953_),
    .Z(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2688_ (.I(net851),
    .ZN(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2689_ (.I(_0956_),
    .Z(_1306_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2690_ (.I(_0958_),
    .Z(_1307_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2691_ (.I(_0960_),
    .Z(_1308_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2692_ (.A1(net882),
    .A2(_1307_),
    .A3(_1308_),
    .ZN(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2693_ (.A1(_1305_),
    .A2(_1306_),
    .B(_1309_),
    .ZN(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2694_ (.A1(net867),
    .A2(_1303_),
    .B1(_1304_),
    .B2(net790),
    .C(_1310_),
    .ZN(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2695_ (.I(_0965_),
    .Z(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2696_ (.I(_0967_),
    .Z(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _2697_ (.I(net479),
    .ZN(_1314_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2698_ (.I(_0970_),
    .Z(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2699_ (.I(_0972_),
    .Z(_1316_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2700_ (.I(net836),
    .ZN(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _2701_ (.A1(_1314_),
    .A2(_1315_),
    .A3(_1148_),
    .B1(_1316_),
    .B2(_1317_),
    .ZN(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2702_ (.A1(net805),
    .A2(_1312_),
    .B1(_1313_),
    .B2(net820),
    .C(_1318_),
    .ZN(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _2703_ (.I(_0977_),
    .Z(_1320_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2704_ (.I(_0979_),
    .Z(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _2705_ (.I(net198),
    .ZN(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2706_ (.I(_0982_),
    .Z(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2707_ (.I(_0984_),
    .Z(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_8 _2708_ (.I(net773),
    .ZN(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _2709_ (.A1(_1322_),
    .A2(_1323_),
    .B1(_1324_),
    .B2(_1325_),
    .ZN(_1326_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2710_ (.A1(net183),
    .A2(_1320_),
    .B1(_1321_),
    .B2(net892),
    .C(_1326_),
    .ZN(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2711_ (.I(_0989_),
    .Z(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2712_ (.I(_0991_),
    .Z(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _2713_ (.I(net189),
    .ZN(_1330_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _2714_ (.I(_0994_),
    .Z(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _2715_ (.I(_0996_),
    .Z(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2716_ (.I(net655),
    .ZN(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _2717_ (.A1(_1330_),
    .A2(_1331_),
    .B1(_1332_),
    .B2(_1333_),
    .ZN(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2718_ (.A1(net811),
    .A2(_1328_),
    .B1(_1329_),
    .B2(net758),
    .C(_1334_),
    .ZN(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _2719_ (.A1(net1797),
    .A2(net1795),
    .A3(_1327_),
    .A4(_1335_),
    .ZN(_1336_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _2720_ (.I(_1002_),
    .Z(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _2721_ (.I(_1004_),
    .Z(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2722_ (.A1(net618),
    .A2(_1337_),
    .B1(_1338_),
    .B2(net634),
    .ZN(_1339_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2723_ (.I(_1007_),
    .Z(_1340_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2724_ (.I(_1009_),
    .Z(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2725_ (.A1(net649),
    .A2(_1340_),
    .B1(_1341_),
    .B2(net540),
    .ZN(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _2726_ (.I(_1012_),
    .Z(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2727_ (.I(_1014_),
    .Z(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2728_ (.A1(net557),
    .A2(_1343_),
    .B1(_1344_),
    .B2(net572),
    .ZN(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2729_ (.I(_1017_),
    .Z(_1346_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2730_ (.I(_1019_),
    .Z(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2731_ (.A1(net416),
    .A2(_1346_),
    .B1(_1347_),
    .B2(net587),
    .ZN(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _2732_ (.A1(_1339_),
    .A2(_1342_),
    .A3(_1345_),
    .A4(_1348_),
    .ZN(_1349_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2733_ (.I(_1023_),
    .Z(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2734_ (.I(_1025_),
    .Z(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2735_ (.A1(net307),
    .A2(_1350_),
    .B1(_1351_),
    .B2(net59),
    .ZN(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2736_ (.I(_1028_),
    .Z(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2737_ (.I(_1030_),
    .Z(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2738_ (.A1(net323),
    .A2(_1353_),
    .B1(_1354_),
    .B2(net74),
    .ZN(_1355_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2739_ (.I(_1033_),
    .Z(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2740_ (.I(_1035_),
    .Z(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2741_ (.A1(net28),
    .A2(_1356_),
    .B1(_1357_),
    .B2(net43),
    .ZN(_1358_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2742_ (.I(_1038_),
    .Z(_1359_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2743_ (.I(_1040_),
    .Z(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2744_ (.A1(net90),
    .A2(_1359_),
    .B1(_1360_),
    .B2(net121),
    .ZN(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _2745_ (.A1(_1352_),
    .A2(_1355_),
    .A3(_1358_),
    .A4(_1361_),
    .ZN(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _2746_ (.A1(_1336_),
    .A2(_1349_),
    .A3(_1362_),
    .ZN(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2747_ (.A1(_1233_),
    .A2(_1234_),
    .B1(net1704),
    .B2(_1363_),
    .ZN(_2312_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2748_ (.I(net45),
    .ZN(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2749_ (.I(net510),
    .ZN(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2750_ (.A1(_1365_),
    .A2(_1236_),
    .A3(_1237_),
    .ZN(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2751_ (.A1(net526),
    .A2(_1239_),
    .A3(_1240_),
    .Z(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2752_ (.I(net604),
    .ZN(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _2753_ (.A1(_1368_),
    .A2(_1243_),
    .A3(_1111_),
    .ZN(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2754_ (.I(net495),
    .ZN(_1370_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2755_ (.A1(_1370_),
    .A2(_1246_),
    .A3(_1247_),
    .ZN(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _2756_ (.A1(_1366_),
    .A2(_1367_),
    .A3(_1369_),
    .A4(_1371_),
    .ZN(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2757_ (.I(net464),
    .ZN(_1373_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2758_ (.I(net449),
    .ZN(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _2759_ (.A1(_1373_),
    .A2(_1253_),
    .A3(_1254_),
    .B1(_1255_),
    .B2(_1374_),
    .ZN(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2760_ (.A1(net402),
    .A2(_1250_),
    .B1(_1251_),
    .B2(net432),
    .C(_1375_),
    .ZN(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _2761_ (.I(net293),
    .ZN(_1377_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _2762_ (.I(net386),
    .ZN(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _2763_ (.A1(_1377_),
    .A2(_1121_),
    .A3(_1262_),
    .B1(_1263_),
    .B2(_1378_),
    .ZN(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2764_ (.A1(net215),
    .A2(_1259_),
    .B1(_1260_),
    .B2(net231),
    .C(_1379_),
    .ZN(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2765_ (.I(net169),
    .ZN(_1381_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2766_ (.I(net153),
    .ZN(_1382_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _2767_ (.A1(_1381_),
    .A2(_1270_),
    .A3(_1271_),
    .B1(_1272_),
    .B2(_1382_),
    .ZN(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2768_ (.A1(net262),
    .A2(_1267_),
    .B1(_1268_),
    .B2(net247),
    .C(_1383_),
    .ZN(_1384_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _2769_ (.A1(_1372_),
    .A2(_1376_),
    .A3(_1380_),
    .A4(_1384_),
    .ZN(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2770_ (.A1(net511),
    .A2(_1277_),
    .B1(_1278_),
    .B2(net106),
    .ZN(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2771_ (.A1(net665),
    .A2(_1280_),
    .B1(_1281_),
    .B2(net138),
    .ZN(_1387_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2772_ (.A1(net728),
    .A2(_1283_),
    .B1(_1284_),
    .B2(net713),
    .ZN(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2773_ (.A1(net682),
    .A2(_1286_),
    .B1(_1287_),
    .B2(net697),
    .ZN(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _2774_ (.A1(_1386_),
    .A2(_1387_),
    .A3(_1388_),
    .A4(_1389_),
    .ZN(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2775_ (.A1(net355),
    .A2(_1290_),
    .B1(_1291_),
    .B2(net743),
    .ZN(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2776_ (.A1(net14),
    .A2(_1293_),
    .B1(_1294_),
    .B2(net356),
    .ZN(_1392_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2777_ (.A1(net371),
    .A2(_1296_),
    .B1(_1297_),
    .B2(net277),
    .ZN(_1393_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2778_ (.A1(net340),
    .A2(_1299_),
    .B(_1138_),
    .ZN(_1394_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _2779_ (.A1(_1391_),
    .A2(_1392_),
    .A3(_1393_),
    .A4(_1394_),
    .ZN(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _2780_ (.A1(_1385_),
    .A2(_1390_),
    .A3(_1395_),
    .ZN(_1396_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2781_ (.I(net852),
    .ZN(_1397_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2782_ (.A1(net883),
    .A2(_1307_),
    .A3(_1308_),
    .ZN(_1398_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2783_ (.A1(_1397_),
    .A2(_1306_),
    .B(_1398_),
    .ZN(_1399_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2784_ (.A1(net868),
    .A2(_1303_),
    .B1(_1304_),
    .B2(net791),
    .C(_1399_),
    .ZN(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _2785_ (.I(net480),
    .ZN(_1401_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _2786_ (.I(net837),
    .ZN(_1402_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _2787_ (.A1(_1401_),
    .A2(_1315_),
    .A3(_1148_),
    .B1(_1316_),
    .B2(_1402_),
    .ZN(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2788_ (.A1(net806),
    .A2(_1312_),
    .B1(_1313_),
    .B2(net821),
    .C(_1403_),
    .ZN(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _2789_ (.I(net199),
    .ZN(_1405_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_8 _2790_ (.I(net774),
    .ZN(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _2791_ (.A1(_1405_),
    .A2(_1323_),
    .B1(_1324_),
    .B2(_1406_),
    .ZN(_1407_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2792_ (.A1(net184),
    .A2(_1320_),
    .B1(_1321_),
    .B2(net893),
    .C(_1407_),
    .ZN(_1408_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _2793_ (.I(net200),
    .ZN(_1409_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2794_ (.I(net666),
    .ZN(_1410_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _2795_ (.A1(_1409_),
    .A2(_1331_),
    .B1(_1332_),
    .B2(_1410_),
    .ZN(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2796_ (.A1(net822),
    .A2(_1328_),
    .B1(_1329_),
    .B2(net759),
    .C(_1411_),
    .ZN(_1412_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _2797_ (.A1(net1793),
    .A2(net1791),
    .A3(_1408_),
    .A4(_1412_),
    .ZN(_1413_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2798_ (.A1(net619),
    .A2(_1337_),
    .B1(_1338_),
    .B2(net635),
    .ZN(_1414_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2799_ (.A1(net650),
    .A2(_1340_),
    .B1(_1341_),
    .B2(net541),
    .ZN(_1415_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2800_ (.A1(net558),
    .A2(_1343_),
    .B1(_1344_),
    .B2(net573),
    .ZN(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2801_ (.A1(net417),
    .A2(_1346_),
    .B1(_1347_),
    .B2(net588),
    .ZN(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _2802_ (.A1(_1414_),
    .A2(_1415_),
    .A3(_1416_),
    .A4(_1417_),
    .ZN(_1418_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2803_ (.A1(net308),
    .A2(_1350_),
    .B1(_1351_),
    .B2(net60),
    .ZN(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2804_ (.A1(net324),
    .A2(_1353_),
    .B1(_1354_),
    .B2(net75),
    .ZN(_1420_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2805_ (.A1(net29),
    .A2(_1356_),
    .B1(_1357_),
    .B2(net44),
    .ZN(_1421_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2806_ (.A1(net91),
    .A2(_1359_),
    .B1(_1360_),
    .B2(net122),
    .ZN(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _2807_ (.A1(_1419_),
    .A2(_1420_),
    .A3(_1421_),
    .A4(_1422_),
    .ZN(_1423_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _2808_ (.A1(_1413_),
    .A2(_1418_),
    .A3(_1423_),
    .ZN(_1424_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2809_ (.A1(_1364_),
    .A2(_1234_),
    .B1(_1396_),
    .B2(_1424_),
    .ZN(_2313_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2810_ (.I(net897),
    .ZN(_1425_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2811_ (.I(net1305),
    .ZN(_1426_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2812_ (.A1(_1426_),
    .A2(_1236_),
    .A3(_1237_),
    .ZN(_1427_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2813_ (.A1(net1319),
    .A2(_1239_),
    .A3(_1240_),
    .Z(_1428_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2814_ (.I(net1386),
    .ZN(_1429_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _2815_ (.I(_0028_),
    .Z(_1430_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _2816_ (.A1(_1429_),
    .A2(_1243_),
    .A3(_1430_),
    .ZN(_1431_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2817_ (.I(net1292),
    .ZN(_1432_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2818_ (.A1(_1432_),
    .A2(_1246_),
    .A3(_1247_),
    .ZN(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _2819_ (.A1(_1427_),
    .A2(_1428_),
    .A3(_1431_),
    .A4(_1433_),
    .ZN(_1434_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2820_ (.I(net1266),
    .ZN(_1435_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2821_ (.I(net1253),
    .ZN(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _2822_ (.A1(_1435_),
    .A2(_1253_),
    .A3(_1254_),
    .B1(_1255_),
    .B2(_1436_),
    .ZN(_1437_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2823_ (.A1(net1212),
    .A2(_1250_),
    .B1(_1251_),
    .B2(net1239),
    .C(_1437_),
    .ZN(_1438_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _2824_ (.I(net1120),
    .ZN(_1439_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2825_ (.I(_0735_),
    .Z(_1440_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2826_ (.I(net1199),
    .ZN(_1441_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _2827_ (.A1(_1439_),
    .A2(_1440_),
    .A3(_1262_),
    .B1(_1263_),
    .B2(_1441_),
    .ZN(_1442_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2828_ (.A1(net1053),
    .A2(_1259_),
    .B1(_1260_),
    .B2(net1066),
    .C(_1442_),
    .ZN(_1443_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2829_ (.I(net1013),
    .ZN(_1444_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2830_ (.I(net999),
    .ZN(_1445_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _2831_ (.A1(_1444_),
    .A2(_1270_),
    .A3(_1271_),
    .B1(_1272_),
    .B2(_1445_),
    .ZN(_1446_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2832_ (.A1(net1092),
    .A2(_1267_),
    .B1(_1268_),
    .B2(net1079),
    .C(_1446_),
    .ZN(_1447_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _2833_ (.A1(net1790),
    .A2(net1789),
    .A3(_1443_),
    .A4(_1447_),
    .ZN(_1448_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2834_ (.A1(net1196),
    .A2(_1277_),
    .B1(_1278_),
    .B2(net959),
    .ZN(_1449_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2835_ (.A1(net1438),
    .A2(_1280_),
    .B1(_1281_),
    .B2(net986),
    .ZN(_1450_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2836_ (.A1(net1492),
    .A2(_1283_),
    .B1(_1284_),
    .B2(net1479),
    .ZN(_1451_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2837_ (.A1(net1453),
    .A2(_1286_),
    .B1(_1287_),
    .B2(net1466),
    .ZN(_1452_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _2838_ (.A1(_1449_),
    .A2(_1450_),
    .A3(_1451_),
    .A4(_1452_),
    .ZN(_1453_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2839_ (.A1(net1172),
    .A2(_1290_),
    .B1(_1291_),
    .B2(net1505),
    .ZN(_1454_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2840_ (.A1(net1647),
    .A2(_1293_),
    .B1(_1294_),
    .B2(net1063),
    .ZN(_1455_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2841_ (.A1(net1186),
    .A2(_1296_),
    .B1(_1297_),
    .B2(net1105),
    .ZN(_1456_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2842_ (.I(_0011_),
    .Z(_1457_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2843_ (.A1(net1159),
    .A2(_1299_),
    .B(_1457_),
    .ZN(_1458_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _2844_ (.A1(_1454_),
    .A2(_1455_),
    .A3(_1456_),
    .A4(_1458_),
    .ZN(_1459_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _2845_ (.A1(_1448_),
    .A2(_1453_),
    .A3(_1459_),
    .ZN(_1460_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2846_ (.I(net1599),
    .ZN(_1461_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2847_ (.A1(net1625),
    .A2(_1307_),
    .A3(_1308_),
    .ZN(_1462_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2848_ (.A1(_1461_),
    .A2(_1306_),
    .B(_1462_),
    .ZN(_1463_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2849_ (.A1(net1612),
    .A2(_1303_),
    .B1(_1304_),
    .B2(net1545),
    .C(_1463_),
    .ZN(_1464_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _2850_ (.I(net1279),
    .ZN(_1465_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2851_ (.I(_1147_),
    .Z(_1466_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2852_ (.I(net1586),
    .ZN(_1467_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _2853_ (.A1(_1465_),
    .A2(_1315_),
    .A3(_1466_),
    .B1(_1316_),
    .B2(_1467_),
    .ZN(_1468_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2854_ (.A1(net1558),
    .A2(_1312_),
    .B1(_1313_),
    .B2(net1572),
    .C(_1468_),
    .ZN(_1469_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2855_ (.I(net1039),
    .ZN(_1470_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_8 _2856_ (.I(net1532),
    .ZN(_1471_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _2857_ (.A1(_1470_),
    .A2(_1323_),
    .B1(_1324_),
    .B2(_1471_),
    .ZN(_1472_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _2858_ (.A1(net1026),
    .A2(_1320_),
    .B1(_1321_),
    .B2(net1596),
    .C(_1472_),
    .ZN(_1473_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _2859_ (.I(net930),
    .ZN(_1474_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2860_ (.I(net1329),
    .ZN(_1475_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _2861_ (.A1(_1474_),
    .A2(_1331_),
    .B1(_1332_),
    .B2(_1475_),
    .ZN(_1476_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2862_ (.A1(net1463),
    .A2(_1328_),
    .B1(_1329_),
    .B2(net1519),
    .C(_1476_),
    .ZN(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _2863_ (.A1(net1787),
    .A2(net1785),
    .A3(_1473_),
    .A4(_1477_),
    .ZN(_1478_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2864_ (.A1(net1399),
    .A2(_1337_),
    .B1(_1338_),
    .B2(net1412),
    .ZN(_1479_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2865_ (.A1(net1425),
    .A2(_1340_),
    .B1(_1341_),
    .B2(net1332),
    .ZN(_1480_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2866_ (.A1(net1346),
    .A2(_1343_),
    .B1(_1344_),
    .B2(net1359),
    .ZN(_1481_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2867_ (.A1(net1225),
    .A2(_1346_),
    .B1(_1347_),
    .B2(net1372),
    .ZN(_1482_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _2868_ (.A1(_1479_),
    .A2(_1480_),
    .A3(_1481_),
    .A4(_1482_),
    .ZN(_1483_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2869_ (.A1(net1133),
    .A2(_1350_),
    .B1(_1351_),
    .B2(net920),
    .ZN(_1484_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2870_ (.A1(net1146),
    .A2(_1353_),
    .B1(_1354_),
    .B2(net933),
    .ZN(_1485_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2871_ (.A1(net1660),
    .A2(_1356_),
    .B1(_1357_),
    .B2(net906),
    .ZN(_1486_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2872_ (.A1(net946),
    .A2(_1359_),
    .B1(_1360_),
    .B2(net972),
    .ZN(_1487_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _2873_ (.A1(_1484_),
    .A2(_1485_),
    .A3(_1486_),
    .A4(_1487_),
    .ZN(_1488_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2874_ (.A1(_1478_),
    .A2(_1483_),
    .A3(_1488_),
    .ZN(_1489_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2875_ (.A1(_1425_),
    .A2(_1234_),
    .B1(_1460_),
    .B2(_1489_),
    .ZN(_2323_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2876_ (.I(net1008),
    .ZN(_1490_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2877_ (.I(net1306),
    .ZN(_1491_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2878_ (.A1(_1491_),
    .A2(_1236_),
    .A3(_1237_),
    .ZN(_1492_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _2879_ (.A1(net1320),
    .A2(_1239_),
    .A3(_1240_),
    .Z(_1493_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2880_ (.I(net1387),
    .ZN(_1494_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _2881_ (.A1(_1494_),
    .A2(_1243_),
    .A3(_1430_),
    .ZN(_1495_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2882_ (.I(net1293),
    .ZN(_1496_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2883_ (.A1(_1496_),
    .A2(_1246_),
    .A3(_1247_),
    .ZN(_1497_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _2884_ (.A1(_1492_),
    .A2(_1493_),
    .A3(_1495_),
    .A4(_1497_),
    .ZN(_1498_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2885_ (.I(net1267),
    .ZN(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2886_ (.I(net1254),
    .ZN(_1500_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _2887_ (.A1(_1499_),
    .A2(_1253_),
    .A3(_1254_),
    .B1(_1255_),
    .B2(_1500_),
    .ZN(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2888_ (.A1(net1213),
    .A2(_1250_),
    .B1(_1251_),
    .B2(net1240),
    .C(_1501_),
    .ZN(_1502_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _2889_ (.I(net1121),
    .ZN(_1503_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2890_ (.I(net1200),
    .ZN(_1504_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _2891_ (.A1(_1503_),
    .A2(_1440_),
    .A3(_1262_),
    .B1(_1263_),
    .B2(_1504_),
    .ZN(_1505_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2892_ (.A1(net1054),
    .A2(_1259_),
    .B1(_1260_),
    .B2(net1067),
    .C(_1505_),
    .ZN(_1506_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2893_ (.I(net1014),
    .ZN(_1507_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2894_ (.I(net1000),
    .ZN(_1508_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _2895_ (.A1(_1507_),
    .A2(_1270_),
    .A3(_1271_),
    .B1(_1272_),
    .B2(_1508_),
    .ZN(_1509_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2896_ (.A1(net1093),
    .A2(_1267_),
    .B1(_1268_),
    .B2(net1080),
    .C(_1509_),
    .ZN(_1510_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _2897_ (.A1(net1784),
    .A2(net1783),
    .A3(_1506_),
    .A4(_1510_),
    .ZN(_1511_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2898_ (.A1(net1207),
    .A2(_1277_),
    .B1(_1278_),
    .B2(net960),
    .ZN(_1512_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2899_ (.A1(net1439),
    .A2(_1280_),
    .B1(_1281_),
    .B2(net987),
    .ZN(_1513_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2900_ (.A1(net1493),
    .A2(_1283_),
    .B1(_1284_),
    .B2(net1480),
    .ZN(_1514_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2901_ (.A1(net1454),
    .A2(_1286_),
    .B1(_1287_),
    .B2(net1467),
    .ZN(_1515_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _2902_ (.A1(_1512_),
    .A2(_1513_),
    .A3(_1514_),
    .A4(_1515_),
    .ZN(_1516_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2903_ (.A1(net1173),
    .A2(_1290_),
    .B1(_1291_),
    .B2(net1506),
    .ZN(_1517_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2904_ (.A1(net1648),
    .A2(_1293_),
    .B1(_1294_),
    .B2(net1074),
    .ZN(_1518_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2905_ (.A1(net1187),
    .A2(_1296_),
    .B1(_1297_),
    .B2(net1106),
    .ZN(_1519_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2906_ (.A1(net1160),
    .A2(_1299_),
    .B(_1457_),
    .ZN(_1520_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _2907_ (.A1(_1517_),
    .A2(_1518_),
    .A3(_1519_),
    .A4(_1520_),
    .ZN(_1521_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _2908_ (.A1(_1511_),
    .A2(_1516_),
    .A3(_1521_),
    .ZN(_1522_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2909_ (.I(net1600),
    .ZN(_1523_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2910_ (.A1(net1626),
    .A2(_1307_),
    .A3(_1308_),
    .ZN(_1524_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2911_ (.A1(_1523_),
    .A2(_1306_),
    .B(_1524_),
    .ZN(_1525_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2912_ (.A1(net1613),
    .A2(_1303_),
    .B1(_1304_),
    .B2(net1546),
    .C(_1525_),
    .ZN(_1526_));
 gf180mcu_fd_sc_mcu7t5v0__inv_4 _2913_ (.I(net1280),
    .ZN(_1527_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2914_ (.I(net1587),
    .ZN(_1528_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _2915_ (.A1(_1527_),
    .A2(_1315_),
    .A3(_1466_),
    .B1(_1316_),
    .B2(_1528_),
    .ZN(_1529_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2916_ (.A1(net1559),
    .A2(_1312_),
    .B1(_1313_),
    .B2(net1573),
    .C(_1529_),
    .ZN(_1530_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2917_ (.I(net1040),
    .ZN(_1531_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_8 _2918_ (.I(net1533),
    .ZN(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _2919_ (.A1(_1531_),
    .A2(_1323_),
    .B1(_1324_),
    .B2(_1532_),
    .ZN(_1533_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _2920_ (.A1(net1027),
    .A2(_1320_),
    .B1(_1321_),
    .B2(net1607),
    .C(_1533_),
    .ZN(_1534_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _2921_ (.I(net941),
    .ZN(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2922_ (.I(net1340),
    .ZN(_1536_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _2923_ (.A1(_1535_),
    .A2(_1331_),
    .B1(_1332_),
    .B2(_1536_),
    .ZN(_1537_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2924_ (.A1(net1474),
    .A2(_1328_),
    .B1(_1329_),
    .B2(net1520),
    .C(_1537_),
    .ZN(_1538_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _2925_ (.A1(net1781),
    .A2(net1779),
    .A3(_1534_),
    .A4(_1538_),
    .ZN(_1539_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2926_ (.A1(net1400),
    .A2(_1337_),
    .B1(_1338_),
    .B2(net1413),
    .ZN(_1540_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2927_ (.A1(net1426),
    .A2(_1340_),
    .B1(_1341_),
    .B2(net1333),
    .ZN(_1541_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2928_ (.A1(net1347),
    .A2(_1343_),
    .B1(_1344_),
    .B2(net1360),
    .ZN(_1542_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2929_ (.A1(net1226),
    .A2(_1346_),
    .B1(_1347_),
    .B2(net1373),
    .ZN(_1543_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _2930_ (.A1(_1540_),
    .A2(_1541_),
    .A3(_1542_),
    .A4(_1543_),
    .ZN(_1544_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2931_ (.A1(net1134),
    .A2(_1350_),
    .B1(_1351_),
    .B2(net921),
    .ZN(_1545_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2932_ (.A1(net1147),
    .A2(_1353_),
    .B1(_1354_),
    .B2(net934),
    .ZN(_1546_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2933_ (.A1(net1661),
    .A2(_1356_),
    .B1(_1357_),
    .B2(net907),
    .ZN(_1547_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2934_ (.A1(net947),
    .A2(_1359_),
    .B1(_1360_),
    .B2(net973),
    .ZN(_1548_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _2935_ (.A1(_1545_),
    .A2(_1546_),
    .A3(_1547_),
    .A4(_1548_),
    .ZN(_1549_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2936_ (.A1(_1539_),
    .A2(_1544_),
    .A3(_1549_),
    .ZN(_1550_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2937_ (.A1(_1490_),
    .A2(_1234_),
    .B1(_1522_),
    .B2(_1550_),
    .ZN(_2326_));
 gf180mcu_fd_sc_mcu7t5v0__inv_3 _2938_ (.I(net1119),
    .ZN(_1551_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2939_ (.I(_0848_),
    .Z(_1552_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2940_ (.I(net1308),
    .ZN(_1553_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2941_ (.I(_0851_),
    .Z(_1554_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2942_ (.I(_0531_),
    .Z(_1555_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2943_ (.A1(_1553_),
    .A2(_1554_),
    .A3(_1555_),
    .ZN(_1556_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2944_ (.I(_0855_),
    .Z(_1557_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2945_ (.I(_0857_),
    .Z(_1558_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _2946_ (.A1(net1321),
    .A2(_1557_),
    .A3(_1558_),
    .Z(_1559_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2947_ (.I(net1388),
    .ZN(_1560_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _2948_ (.I(_0861_),
    .Z(_1561_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _2949_ (.A1(_1560_),
    .A2(_1561_),
    .A3(_1430_),
    .ZN(_1562_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2950_ (.I(net1294),
    .ZN(_1563_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2951_ (.I(_0865_),
    .Z(_1564_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2952_ (.I(_0867_),
    .Z(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2953_ (.A1(_1563_),
    .A2(_1564_),
    .A3(_1565_),
    .ZN(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _2954_ (.A1(_1556_),
    .A2(_1559_),
    .A3(_1562_),
    .A4(_1566_),
    .ZN(_1567_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _2955_ (.I(_0871_),
    .Z(_1568_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _2956_ (.I(_0873_),
    .Z(_1569_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2957_ (.I(net1268),
    .ZN(_1570_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2958_ (.I(_0876_),
    .Z(_1571_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2959_ (.I(_0288_),
    .Z(_1572_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2960_ (.I(_0879_),
    .Z(_1573_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2961_ (.I(net1255),
    .ZN(_1574_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _2962_ (.A1(_1570_),
    .A2(_1571_),
    .A3(_1572_),
    .B1(_1573_),
    .B2(_1574_),
    .ZN(_1575_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2963_ (.A1(net1214),
    .A2(_1568_),
    .B1(_1569_),
    .B2(net1242),
    .C(_1575_),
    .ZN(_1576_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2964_ (.I(_0884_),
    .Z(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2965_ (.I(_0886_),
    .Z(_1578_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _2966_ (.I(net1122),
    .ZN(_1579_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2967_ (.I(_0889_),
    .Z(_1580_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2968_ (.I(_0891_),
    .Z(_1581_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2969_ (.I(net1201),
    .ZN(_1582_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _2970_ (.A1(_1579_),
    .A2(_1440_),
    .A3(_1580_),
    .B1(_1581_),
    .B2(_1582_),
    .ZN(_1583_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2971_ (.A1(net1055),
    .A2(_1577_),
    .B1(_1578_),
    .B2(net1068),
    .C(_1583_),
    .ZN(_1584_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2972_ (.I(_0896_),
    .Z(_1585_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2973_ (.I(_0898_),
    .Z(_1586_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2974_ (.I(net1015),
    .ZN(_1587_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2975_ (.I(_0901_),
    .Z(_1588_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _2976_ (.I(_0102_),
    .Z(_1589_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2977_ (.I(_0904_),
    .Z(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2978_ (.I(net1001),
    .ZN(_1591_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _2979_ (.A1(_1587_),
    .A2(_1588_),
    .A3(_1589_),
    .B1(_1590_),
    .B2(_1591_),
    .ZN(_1592_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2980_ (.A1(net1094),
    .A2(_1585_),
    .B1(_1586_),
    .B2(net1081),
    .C(_1592_),
    .ZN(_1593_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _2981_ (.A1(_1567_),
    .A2(_1576_),
    .A3(_1584_),
    .A4(_1593_),
    .ZN(_1594_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2982_ (.I(_0910_),
    .Z(_1595_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2983_ (.I(_0912_),
    .Z(_1596_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2984_ (.A1(net1218),
    .A2(_1595_),
    .B1(_1596_),
    .B2(net961),
    .ZN(_1597_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2985_ (.I(_0915_),
    .Z(_1598_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2986_ (.I(_0917_),
    .Z(_1599_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2987_ (.A1(net1441),
    .A2(_1598_),
    .B1(_1599_),
    .B2(net988),
    .ZN(_1600_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2988_ (.I(_0920_),
    .Z(_1601_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2989_ (.I(_0922_),
    .Z(_1602_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2990_ (.A1(net1494),
    .A2(_1601_),
    .B1(_1602_),
    .B2(net1481),
    .ZN(_1603_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2991_ (.I(_0925_),
    .Z(_1604_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2992_ (.I(_0927_),
    .Z(_1605_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2993_ (.A1(net1455),
    .A2(_1604_),
    .B1(_1605_),
    .B2(net1468),
    .ZN(_1606_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _2994_ (.A1(_1597_),
    .A2(_1600_),
    .A3(_1603_),
    .A4(_1606_),
    .ZN(_1607_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2995_ (.I(_0931_),
    .Z(_1608_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2996_ (.I(_0933_),
    .Z(_1609_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2997_ (.A1(net1175),
    .A2(_1608_),
    .B1(_1609_),
    .B2(net1508),
    .ZN(_1610_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2998_ (.I(_0936_),
    .Z(_1611_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2999_ (.I(_0938_),
    .Z(_1612_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _3000_ (.A1(net1649),
    .A2(_1611_),
    .B1(_1612_),
    .B2(net1085),
    .ZN(_1613_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3001_ (.I(_0941_),
    .Z(_1614_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3002_ (.I(_0943_),
    .Z(_1615_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3003_ (.A1(net1188),
    .A2(_1614_),
    .B1(_1615_),
    .B2(net1108),
    .ZN(_1616_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3004_ (.I(_0946_),
    .Z(_1617_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3005_ (.A1(net1161),
    .A2(_1617_),
    .B(_1457_),
    .ZN(_1618_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3006_ (.A1(_1610_),
    .A2(_1613_),
    .A3(_1616_),
    .A4(_1618_),
    .ZN(_1619_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3007_ (.A1(_1594_),
    .A2(_1607_),
    .A3(_1619_),
    .ZN(_1620_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3008_ (.I(_0951_),
    .Z(_1621_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3009_ (.I(_0953_),
    .Z(_1622_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3010_ (.I(net1601),
    .ZN(_1623_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3011_ (.I(_0956_),
    .Z(_1624_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3012_ (.I(_0958_),
    .Z(_1625_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3013_ (.I(_0960_),
    .Z(_1626_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3014_ (.A1(net1627),
    .A2(_1625_),
    .A3(_1626_),
    .ZN(_1627_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3015_ (.A1(_1623_),
    .A2(_1624_),
    .B(_1627_),
    .ZN(_1628_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3016_ (.A1(net1614),
    .A2(_1621_),
    .B1(_1622_),
    .B2(net1547),
    .C(_1628_),
    .ZN(_1629_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3017_ (.I(_0965_),
    .Z(_1630_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3018_ (.I(_0967_),
    .Z(_1631_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _3019_ (.I(net1281),
    .ZN(_1632_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3020_ (.I(_0970_),
    .Z(_1633_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3021_ (.I(_0972_),
    .Z(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3022_ (.I(net1588),
    .ZN(_1635_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _3023_ (.A1(_1632_),
    .A2(_1633_),
    .A3(_1466_),
    .B1(_1634_),
    .B2(_1635_),
    .ZN(_1636_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3024_ (.A1(net1560),
    .A2(_1630_),
    .B1(_1631_),
    .B2(net1575),
    .C(_1636_),
    .ZN(_1637_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3025_ (.I(_0977_),
    .Z(_1638_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3026_ (.I(_0979_),
    .Z(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3027_ (.I(net1042),
    .ZN(_1640_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3028_ (.I(_0982_),
    .Z(_1641_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3029_ (.I(_0984_),
    .Z(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_8 _3030_ (.I(net1534),
    .ZN(_1643_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _3031_ (.A1(_1640_),
    .A2(_1641_),
    .B1(_1642_),
    .B2(_1643_),
    .ZN(_1644_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3032_ (.A1(net1028),
    .A2(_1638_),
    .B1(_1639_),
    .B2(net1618),
    .C(_1644_),
    .ZN(_1645_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3033_ (.I(_0989_),
    .Z(_1646_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3034_ (.I(_0991_),
    .Z(_1647_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _3035_ (.I(net952),
    .ZN(_1648_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3036_ (.I(_0994_),
    .Z(_1649_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3037_ (.I(_0996_),
    .Z(_1650_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3038_ (.I(net1352),
    .ZN(_1651_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _3039_ (.A1(_1648_),
    .A2(_1649_),
    .B1(_1650_),
    .B2(_1651_),
    .ZN(_1652_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3040_ (.A1(net1485),
    .A2(_1646_),
    .B1(_1647_),
    .B2(net1521),
    .C(_1652_),
    .ZN(_1653_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3041_ (.A1(net1778),
    .A2(net1777),
    .A3(_1645_),
    .A4(net1776),
    .ZN(_1654_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3042_ (.I(_1002_),
    .Z(_1655_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3043_ (.I(_1004_),
    .Z(_1656_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _3044_ (.A1(net1401),
    .A2(_1655_),
    .B1(_1656_),
    .B2(net1414),
    .ZN(_1657_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3045_ (.I(_1007_),
    .Z(_1658_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3046_ (.I(_1009_),
    .Z(_1659_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3047_ (.A1(net1427),
    .A2(_1658_),
    .B1(_1659_),
    .B2(net1334),
    .ZN(_1660_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3048_ (.I(_1012_),
    .Z(_1661_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3049_ (.I(_1014_),
    .Z(_1662_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _3050_ (.A1(net1348),
    .A2(_1661_),
    .B1(_1662_),
    .B2(net1361),
    .ZN(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3051_ (.I(_1017_),
    .Z(_1664_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3052_ (.I(_1019_),
    .Z(_1665_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3053_ (.A1(net1227),
    .A2(_1664_),
    .B1(_1665_),
    .B2(net1375),
    .ZN(_1666_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _3054_ (.A1(_1657_),
    .A2(_1660_),
    .A3(_1663_),
    .A4(_1666_),
    .ZN(_1667_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3055_ (.I(_1023_),
    .Z(_1668_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3056_ (.I(_1025_),
    .Z(_1669_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3057_ (.A1(net1135),
    .A2(_1668_),
    .B1(_1669_),
    .B2(net922),
    .ZN(_1670_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3058_ (.I(_1028_),
    .Z(_1671_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3059_ (.I(_1030_),
    .Z(_1672_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3060_ (.A1(net1148),
    .A2(_1671_),
    .B1(_1672_),
    .B2(net935),
    .ZN(_1673_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3061_ (.I(_1033_),
    .Z(_1674_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3062_ (.I(_1035_),
    .Z(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3063_ (.A1(net1662),
    .A2(_1674_),
    .B1(_1675_),
    .B2(net909),
    .ZN(_1676_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3064_ (.I(_1038_),
    .Z(_1677_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3065_ (.I(_1040_),
    .Z(_1678_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _3066_ (.A1(net948),
    .A2(_1677_),
    .B1(_1678_),
    .B2(net975),
    .ZN(_1679_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _3067_ (.A1(_1670_),
    .A2(_1673_),
    .A3(_1676_),
    .A4(_1679_),
    .ZN(_1680_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3068_ (.A1(_1654_),
    .A2(_1667_),
    .A3(_1680_),
    .ZN(_1681_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3069_ (.A1(_1551_),
    .A2(_1552_),
    .B1(_1620_),
    .B2(_1681_),
    .ZN(_2327_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _3070_ (.I(net1230),
    .ZN(_1682_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3071_ (.I(net1309),
    .ZN(_1683_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3072_ (.A1(_1683_),
    .A2(_1554_),
    .A3(_1555_),
    .ZN(_1684_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _3073_ (.A1(net1322),
    .A2(_1557_),
    .A3(_1558_),
    .Z(_1685_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3074_ (.I(net1389),
    .ZN(_1686_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _3075_ (.A1(_1686_),
    .A2(_1561_),
    .A3(_1430_),
    .ZN(_1687_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3076_ (.I(net1295),
    .ZN(_1688_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3077_ (.A1(_1688_),
    .A2(_1564_),
    .A3(_1565_),
    .ZN(_1689_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _3078_ (.A1(_1684_),
    .A2(_1685_),
    .A3(_1687_),
    .A4(_1689_),
    .ZN(_1690_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3079_ (.I(net1269),
    .ZN(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3080_ (.I(net1256),
    .ZN(_1692_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _3081_ (.A1(_1691_),
    .A2(_1571_),
    .A3(_1572_),
    .B1(_1573_),
    .B2(_1692_),
    .ZN(_1693_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _3082_ (.A1(net1215),
    .A2(_1568_),
    .B1(_1569_),
    .B2(net1243),
    .C(_1693_),
    .ZN(_1694_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _3083_ (.I(net1123),
    .ZN(_1695_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3084_ (.I(net1202),
    .ZN(_1696_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _3085_ (.A1(_1695_),
    .A2(_1440_),
    .A3(_1580_),
    .B1(_1581_),
    .B2(_1696_),
    .ZN(_1697_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3086_ (.A1(net1056),
    .A2(_1577_),
    .B1(_1578_),
    .B2(net1069),
    .C(_1697_),
    .ZN(_1698_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3087_ (.I(net1016),
    .ZN(_1699_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3088_ (.I(net1002),
    .ZN(_1700_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _3089_ (.A1(_1699_),
    .A2(_1588_),
    .A3(_1589_),
    .B1(_1590_),
    .B2(_1700_),
    .ZN(_1701_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3090_ (.A1(net1095),
    .A2(_1585_),
    .B1(_1586_),
    .B2(net1082),
    .C(_1701_),
    .ZN(_1702_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _3091_ (.A1(net1775),
    .A2(net1774),
    .A3(_1698_),
    .A4(_1702_),
    .ZN(_1703_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _3092_ (.A1(net1229),
    .A2(_1595_),
    .B1(_1596_),
    .B2(net962),
    .ZN(_1704_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3093_ (.A1(net1442),
    .A2(_1598_),
    .B1(_1599_),
    .B2(net989),
    .ZN(_1705_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _3094_ (.A1(net1495),
    .A2(_1601_),
    .B1(_1602_),
    .B2(net1482),
    .ZN(_1706_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _3095_ (.A1(net1456),
    .A2(_1604_),
    .B1(_1605_),
    .B2(net1469),
    .ZN(_1707_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _3096_ (.A1(_1704_),
    .A2(_1705_),
    .A3(_1706_),
    .A4(_1707_),
    .ZN(_1708_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3097_ (.A1(net1176),
    .A2(_1608_),
    .B1(_1609_),
    .B2(net1509),
    .ZN(_1709_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _3098_ (.A1(net1650),
    .A2(_1611_),
    .B1(_1612_),
    .B2(net1096),
    .ZN(_1710_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3099_ (.A1(net1189),
    .A2(_1614_),
    .B1(_1615_),
    .B2(net1109),
    .ZN(_1711_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3100_ (.A1(net1162),
    .A2(_1617_),
    .B(_1457_),
    .ZN(_1712_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3101_ (.A1(_1709_),
    .A2(_1710_),
    .A3(_1711_),
    .A4(_1712_),
    .ZN(_1713_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3102_ (.A1(_1703_),
    .A2(_1708_),
    .A3(_1713_),
    .ZN(_1714_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3103_ (.I(net1602),
    .ZN(_1715_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3104_ (.A1(net1628),
    .A2(_1625_),
    .A3(_1626_),
    .ZN(_1716_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3105_ (.A1(_1715_),
    .A2(_1624_),
    .B(_1716_),
    .ZN(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3106_ (.A1(net1615),
    .A2(_1621_),
    .B1(_1622_),
    .B2(net1548),
    .C(_1717_),
    .ZN(_1718_));
 gf180mcu_fd_sc_mcu7t5v0__inv_4 _3107_ (.I(net1282),
    .ZN(_1719_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3108_ (.I(net1589),
    .ZN(_1720_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _3109_ (.A1(_1719_),
    .A2(_1633_),
    .A3(_1466_),
    .B1(_1634_),
    .B2(_1720_),
    .ZN(_1721_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3110_ (.A1(net1561),
    .A2(_1630_),
    .B1(_1631_),
    .B2(net1576),
    .C(_1721_),
    .ZN(_1722_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3111_ (.I(net1043),
    .ZN(_1723_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_8 _3112_ (.I(net1535),
    .ZN(_1724_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _3113_ (.A1(_1723_),
    .A2(_1641_),
    .B1(_1642_),
    .B2(_1724_),
    .ZN(_1725_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3114_ (.A1(net1029),
    .A2(_1638_),
    .B1(_1639_),
    .B2(net1629),
    .C(_1725_),
    .ZN(_1726_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _3115_ (.I(net963),
    .ZN(_1727_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3116_ (.I(net1363),
    .ZN(_1728_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _3117_ (.A1(_1727_),
    .A2(_1649_),
    .B1(_1650_),
    .B2(_1728_),
    .ZN(_1729_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3118_ (.A1(net1496),
    .A2(_1646_),
    .B1(_1647_),
    .B2(net1522),
    .C(_1729_),
    .ZN(_1730_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3119_ (.A1(net1773),
    .A2(net1772),
    .A3(_1726_),
    .A4(net1771),
    .ZN(_1731_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _3120_ (.A1(net1402),
    .A2(_1655_),
    .B1(_1656_),
    .B2(net1415),
    .ZN(_1732_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3121_ (.A1(net1428),
    .A2(_1658_),
    .B1(_1659_),
    .B2(net1335),
    .ZN(_1733_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3122_ (.A1(net1349),
    .A2(_1661_),
    .B1(_1662_),
    .B2(net1362),
    .ZN(_1734_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3123_ (.A1(net1228),
    .A2(_1664_),
    .B1(_1665_),
    .B2(net1376),
    .ZN(_1735_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _3124_ (.A1(_1732_),
    .A2(_1733_),
    .A3(_1734_),
    .A4(_1735_),
    .ZN(_1736_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3125_ (.A1(net1136),
    .A2(_1668_),
    .B1(_1669_),
    .B2(net923),
    .ZN(_1737_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3126_ (.A1(net1149),
    .A2(_1671_),
    .B1(_1672_),
    .B2(net936),
    .ZN(_1738_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3127_ (.A1(net1663),
    .A2(_1674_),
    .B1(_1675_),
    .B2(net910),
    .ZN(_1739_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _3128_ (.A1(net949),
    .A2(_1677_),
    .B1(_1678_),
    .B2(net976),
    .ZN(_1740_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _3129_ (.A1(_1737_),
    .A2(_1738_),
    .A3(_1739_),
    .A4(_1740_),
    .ZN(_1741_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3130_ (.A1(_1731_),
    .A2(_1736_),
    .A3(_1741_),
    .ZN(_1742_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3131_ (.A1(_1682_),
    .A2(_1552_),
    .B1(_1714_),
    .B2(_1742_),
    .ZN(_2328_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3132_ (.I(net1341),
    .ZN(_1743_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3133_ (.I(net1310),
    .ZN(_1744_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3134_ (.A1(_1744_),
    .A2(_1554_),
    .A3(_1555_),
    .ZN(_1745_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3135_ (.A1(net1323),
    .A2(_1557_),
    .A3(_1558_),
    .Z(_1746_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3136_ (.I(net1390),
    .ZN(_1747_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _3137_ (.I(_0028_),
    .Z(_1748_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _3138_ (.A1(_1747_),
    .A2(_1561_),
    .A3(_1748_),
    .ZN(_1749_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3139_ (.I(net1297),
    .ZN(_1750_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3140_ (.A1(_1750_),
    .A2(_1564_),
    .A3(_1565_),
    .ZN(_1751_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _3141_ (.A1(_1745_),
    .A2(_1746_),
    .A3(_1749_),
    .A4(_1751_),
    .ZN(_1752_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3142_ (.I(net1270),
    .ZN(_1753_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3143_ (.I(net1257),
    .ZN(_1754_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _3144_ (.A1(_1753_),
    .A2(_1571_),
    .A3(_1572_),
    .B1(_1573_),
    .B2(_1754_),
    .ZN(_1755_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3145_ (.A1(net1216),
    .A2(_1568_),
    .B1(_1569_),
    .B2(net1244),
    .C(_1755_),
    .ZN(_1756_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _3146_ (.I(net1124),
    .ZN(_1757_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3147_ (.I(_0735_),
    .Z(_1758_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3148_ (.I(net1203),
    .ZN(_1759_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _3149_ (.A1(_1757_),
    .A2(_1758_),
    .A3(_1580_),
    .B1(_1581_),
    .B2(_1759_),
    .ZN(_1760_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3150_ (.A1(net1057),
    .A2(_1577_),
    .B1(_1578_),
    .B2(net1070),
    .C(_1760_),
    .ZN(_1761_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3151_ (.I(net1017),
    .ZN(_1762_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3152_ (.I(net1003),
    .ZN(_1763_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _3153_ (.A1(_1762_),
    .A2(_1588_),
    .A3(_1589_),
    .B1(_1590_),
    .B2(_1763_),
    .ZN(_1764_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3154_ (.A1(net1097),
    .A2(_1585_),
    .B1(_1586_),
    .B2(net1083),
    .C(_1764_),
    .ZN(_1765_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3155_ (.A1(_1752_),
    .A2(_1756_),
    .A3(_1761_),
    .A4(_1765_),
    .ZN(_1766_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _3156_ (.A1(net1241),
    .A2(_1595_),
    .B1(_1596_),
    .B2(net964),
    .ZN(_1767_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3157_ (.A1(net1443),
    .A2(_1598_),
    .B1(_1599_),
    .B2(net990),
    .ZN(_1768_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _3158_ (.A1(net1497),
    .A2(_1601_),
    .B1(_1602_),
    .B2(net1483),
    .ZN(_1769_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _3159_ (.A1(net1457),
    .A2(_1604_),
    .B1(_1605_),
    .B2(net1470),
    .ZN(_1770_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _3160_ (.A1(_1767_),
    .A2(_1768_),
    .A3(_1769_),
    .A4(_1770_),
    .ZN(_1771_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3161_ (.A1(net1177),
    .A2(_1608_),
    .B1(_1609_),
    .B2(net1510),
    .ZN(_1772_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _3162_ (.A1(net1651),
    .A2(_1611_),
    .B1(_1612_),
    .B2(net1107),
    .ZN(_1773_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3163_ (.A1(net1190),
    .A2(_1614_),
    .B1(_1615_),
    .B2(net1110),
    .ZN(_1774_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3164_ (.I(_0011_),
    .Z(_1775_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3165_ (.A1(net1164),
    .A2(_1617_),
    .B(_1775_),
    .ZN(_1776_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3166_ (.A1(_1772_),
    .A2(_1773_),
    .A3(_1774_),
    .A4(_1776_),
    .ZN(_1777_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3167_ (.A1(_1766_),
    .A2(_1771_),
    .A3(_1777_),
    .ZN(_1778_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3168_ (.I(net1603),
    .ZN(_1779_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3169_ (.A1(net1630),
    .A2(_1625_),
    .A3(_1626_),
    .ZN(_1780_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3170_ (.A1(_1779_),
    .A2(_1624_),
    .B(_1780_),
    .ZN(_1781_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3171_ (.A1(net1616),
    .A2(_1621_),
    .B1(_1622_),
    .B2(net1549),
    .C(_1781_),
    .ZN(_1782_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _3172_ (.I(net1283),
    .ZN(_1783_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3173_ (.I(_1147_),
    .Z(_1784_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3174_ (.I(net1590),
    .ZN(_1785_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _3175_ (.A1(_1783_),
    .A2(_1633_),
    .A3(_1784_),
    .B1(_1634_),
    .B2(_1785_),
    .ZN(_1786_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3176_ (.A1(net1564),
    .A2(_1630_),
    .B1(_1631_),
    .B2(net1577),
    .C(_1786_),
    .ZN(_1787_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3177_ (.I(net1044),
    .ZN(_1788_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_8 _3178_ (.I(net1536),
    .ZN(_1789_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _3179_ (.A1(_1788_),
    .A2(_1641_),
    .B1(_1642_),
    .B2(_1789_),
    .ZN(_1790_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3180_ (.A1(net1031),
    .A2(_1638_),
    .B1(_1639_),
    .B2(net1638),
    .C(_1790_),
    .ZN(_1791_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _3181_ (.I(net974),
    .ZN(_1792_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3182_ (.I(net1374),
    .ZN(_1793_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _3183_ (.A1(_1792_),
    .A2(_1649_),
    .B1(_1650_),
    .B2(_1793_),
    .ZN(_1794_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3184_ (.A1(net1507),
    .A2(_1646_),
    .B1(_1647_),
    .B2(net1523),
    .C(_1794_),
    .ZN(_1795_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3185_ (.A1(net1770),
    .A2(net1769),
    .A3(_1791_),
    .A4(net1768),
    .ZN(_1796_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _3186_ (.A1(net1403),
    .A2(_1655_),
    .B1(_1656_),
    .B2(net1416),
    .ZN(_1797_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3187_ (.A1(net1430),
    .A2(_1658_),
    .B1(_1659_),
    .B2(net1336),
    .ZN(_1798_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3188_ (.A1(net1350),
    .A2(_1661_),
    .B1(_1662_),
    .B2(net1364),
    .ZN(_1799_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3189_ (.A1(net1231),
    .A2(_1664_),
    .B1(_1665_),
    .B2(net1377),
    .ZN(_1800_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _3190_ (.A1(_1797_),
    .A2(_1798_),
    .A3(_1799_),
    .A4(_1800_),
    .ZN(_1801_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3191_ (.A1(net1137),
    .A2(_1668_),
    .B1(_1669_),
    .B2(net924),
    .ZN(_1802_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3192_ (.A1(net1150),
    .A2(_1671_),
    .B1(_1672_),
    .B2(net937),
    .ZN(_1803_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3193_ (.A1(net898),
    .A2(_1674_),
    .B1(_1675_),
    .B2(net911),
    .ZN(_1804_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _3194_ (.A1(net950),
    .A2(_1677_),
    .B1(_1678_),
    .B2(net977),
    .ZN(_1805_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _3195_ (.A1(_1802_),
    .A2(_1803_),
    .A3(_1804_),
    .A4(_1805_),
    .ZN(_1806_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3196_ (.A1(_1796_),
    .A2(_1801_),
    .A3(_1806_),
    .ZN(_1807_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3197_ (.A1(_1743_),
    .A2(_1552_),
    .B1(_1778_),
    .B2(_1807_),
    .ZN(_2329_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3198_ (.I(net1452),
    .ZN(_1808_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3199_ (.I(net1311),
    .ZN(_1809_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3200_ (.A1(_1809_),
    .A2(_1554_),
    .A3(_1555_),
    .ZN(_1810_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3201_ (.A1(net1324),
    .A2(_1557_),
    .A3(_1558_),
    .Z(_1811_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3202_ (.I(net1391),
    .ZN(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _3203_ (.A1(_1812_),
    .A2(_1561_),
    .A3(_1748_),
    .ZN(_1813_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3204_ (.I(net1298),
    .ZN(_1814_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _3205_ (.A1(_1814_),
    .A2(_1564_),
    .A3(_1565_),
    .ZN(_1815_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _3206_ (.A1(_1810_),
    .A2(_1811_),
    .A3(_1813_),
    .A4(_1815_),
    .ZN(_1816_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3207_ (.I(net1271),
    .ZN(_1817_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3208_ (.I(net1258),
    .ZN(_1818_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _3209_ (.A1(_1817_),
    .A2(_1571_),
    .A3(_1572_),
    .B1(_1573_),
    .B2(_1818_),
    .ZN(_1819_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3210_ (.A1(net1217),
    .A2(_1568_),
    .B1(_1569_),
    .B2(net1245),
    .C(_1819_),
    .ZN(_1820_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _3211_ (.I(net1125),
    .ZN(_1821_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3212_ (.I(net1204),
    .ZN(_1822_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _3213_ (.A1(_1821_),
    .A2(_1758_),
    .A3(_1580_),
    .B1(_1581_),
    .B2(_1822_),
    .ZN(_1823_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3214_ (.A1(net1058),
    .A2(_1577_),
    .B1(_1578_),
    .B2(net1071),
    .C(_1823_),
    .ZN(_1824_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3215_ (.I(net1018),
    .ZN(_1825_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3216_ (.I(net1004),
    .ZN(_1826_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _3217_ (.A1(_1825_),
    .A2(_1588_),
    .A3(_1589_),
    .B1(_1590_),
    .B2(_1826_),
    .ZN(_1827_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3218_ (.A1(net1098),
    .A2(_1585_),
    .B1(_1586_),
    .B2(net1084),
    .C(_1827_),
    .ZN(_1828_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3219_ (.A1(_1816_),
    .A2(_1820_),
    .A3(_1824_),
    .A4(_1828_),
    .ZN(_1829_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _3220_ (.A1(net1252),
    .A2(_1595_),
    .B1(_1596_),
    .B2(net965),
    .ZN(_1830_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3221_ (.A1(net1444),
    .A2(_1598_),
    .B1(_1599_),
    .B2(net991),
    .ZN(_1831_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _3222_ (.A1(net1498),
    .A2(_1601_),
    .B1(_1602_),
    .B2(net1484),
    .ZN(_1832_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _3223_ (.A1(net1458),
    .A2(_1604_),
    .B1(_1605_),
    .B2(net1471),
    .ZN(_1833_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _3224_ (.A1(_1830_),
    .A2(_1831_),
    .A3(_1832_),
    .A4(_1833_),
    .ZN(_1834_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3225_ (.A1(net1178),
    .A2(_1608_),
    .B1(_1609_),
    .B2(net1511),
    .ZN(_1835_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _3226_ (.A1(net1652),
    .A2(_1611_),
    .B1(_1612_),
    .B2(net1118),
    .ZN(_1836_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3227_ (.A1(net1191),
    .A2(_1614_),
    .B1(_1615_),
    .B2(net1111),
    .ZN(_1837_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3228_ (.A1(net1165),
    .A2(_1617_),
    .B(_1775_),
    .ZN(_1838_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3229_ (.A1(_1835_),
    .A2(_1836_),
    .A3(_1837_),
    .A4(_1838_),
    .ZN(_1839_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3230_ (.A1(_1829_),
    .A2(_1834_),
    .A3(_1839_),
    .ZN(_1840_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3231_ (.I(net1604),
    .ZN(_1841_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3232_ (.A1(net1631),
    .A2(_1625_),
    .A3(_1626_),
    .ZN(_1842_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3233_ (.A1(_1841_),
    .A2(_1624_),
    .B(_1842_),
    .ZN(_1843_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3234_ (.A1(net1617),
    .A2(_1621_),
    .B1(_1622_),
    .B2(net1550),
    .C(_1843_),
    .ZN(_1844_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _3235_ (.I(net1284),
    .ZN(_1845_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3236_ (.I(net1591),
    .ZN(_1846_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _3237_ (.A1(_1845_),
    .A2(_1633_),
    .A3(_1784_),
    .B1(_1634_),
    .B2(_1846_),
    .ZN(_1847_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3238_ (.A1(net1565),
    .A2(_1630_),
    .B1(_1631_),
    .B2(net1578),
    .C(_1847_),
    .ZN(_1848_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3239_ (.I(net1045),
    .ZN(_1849_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_8 _3240_ (.I(net1537),
    .ZN(_1850_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _3241_ (.A1(_1849_),
    .A2(_1641_),
    .B1(_1642_),
    .B2(_1850_),
    .ZN(_1851_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3242_ (.A1(net1032),
    .A2(_1638_),
    .B1(_1639_),
    .B2(net1639),
    .C(_1851_),
    .ZN(_1852_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _3243_ (.I(net985),
    .ZN(_1853_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3244_ (.I(net1385),
    .ZN(_1854_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _3245_ (.A1(_1853_),
    .A2(_1649_),
    .B1(_1650_),
    .B2(_1854_),
    .ZN(_1855_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3246_ (.A1(net1518),
    .A2(_1646_),
    .B1(_1647_),
    .B2(net1524),
    .C(_1855_),
    .ZN(_1856_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3247_ (.A1(net1767),
    .A2(net1766),
    .A3(_1852_),
    .A4(net1765),
    .ZN(_1857_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _3248_ (.A1(net1404),
    .A2(_1655_),
    .B1(_1656_),
    .B2(net1417),
    .ZN(_1858_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3249_ (.A1(net1431),
    .A2(_1658_),
    .B1(_1659_),
    .B2(net1337),
    .ZN(_1859_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3250_ (.A1(net1351),
    .A2(_1661_),
    .B1(_1662_),
    .B2(net1365),
    .ZN(_1860_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3251_ (.A1(net1232),
    .A2(_1664_),
    .B1(_1665_),
    .B2(net1378),
    .ZN(_1861_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _3252_ (.A1(_1858_),
    .A2(_1859_),
    .A3(_1860_),
    .A4(_1861_),
    .ZN(_1862_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3253_ (.A1(net1138),
    .A2(_1668_),
    .B1(_1669_),
    .B2(net925),
    .ZN(_1863_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3254_ (.A1(net1151),
    .A2(_1671_),
    .B1(_1672_),
    .B2(net938),
    .ZN(_1864_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3255_ (.A1(net899),
    .A2(_1674_),
    .B1(_1675_),
    .B2(net912),
    .ZN(_1865_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _3256_ (.A1(net951),
    .A2(_1677_),
    .B1(_1678_),
    .B2(net978),
    .ZN(_1866_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _3257_ (.A1(_1863_),
    .A2(_1864_),
    .A3(_1865_),
    .A4(_1866_),
    .ZN(_1867_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3258_ (.A1(_1857_),
    .A2(_1862_),
    .A3(_1867_),
    .ZN(_1868_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3259_ (.A1(_1808_),
    .A2(_1552_),
    .B1(_1840_),
    .B2(_1868_),
    .ZN(_2330_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3260_ (.I(net1563),
    .ZN(_1869_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3261_ (.I(_0848_),
    .Z(_1870_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3262_ (.I(net1312),
    .ZN(_1871_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3263_ (.I(_0851_),
    .Z(_1872_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3264_ (.I(_0237_),
    .Z(_1873_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3265_ (.A1(_1871_),
    .A2(_1872_),
    .A3(_1873_),
    .ZN(_1874_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3266_ (.I(_0855_),
    .Z(_1875_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3267_ (.I(_0857_),
    .Z(_1876_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _3268_ (.A1(net1325),
    .A2(_1875_),
    .A3(_1876_),
    .Z(_1877_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3269_ (.I(net1392),
    .ZN(_1878_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _3270_ (.I(_0861_),
    .Z(_1879_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _3271_ (.A1(_1878_),
    .A2(_1879_),
    .A3(_1748_),
    .ZN(_1880_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3272_ (.I(net1299),
    .ZN(_1881_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3273_ (.I(_0865_),
    .Z(_1882_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3274_ (.I(_0867_),
    .Z(_1883_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3275_ (.A1(_1881_),
    .A2(_1882_),
    .A3(_1883_),
    .ZN(_1884_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _3276_ (.A1(_1874_),
    .A2(_1877_),
    .A3(_1880_),
    .A4(_1884_),
    .ZN(_1885_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3277_ (.I(_0871_),
    .Z(_1886_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3278_ (.I(_0873_),
    .Z(_1887_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3279_ (.I(net1272),
    .ZN(_1888_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3280_ (.I(_0876_),
    .Z(_1889_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3281_ (.I(_0288_),
    .Z(_1890_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3282_ (.I(_0879_),
    .Z(_1891_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3283_ (.I(net1259),
    .ZN(_1892_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _3284_ (.A1(_1888_),
    .A2(_1889_),
    .A3(_1890_),
    .B1(_1891_),
    .B2(_1892_),
    .ZN(_1893_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3285_ (.A1(net1219),
    .A2(_1886_),
    .B1(_1887_),
    .B2(net1246),
    .C(_1893_),
    .ZN(_1894_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3286_ (.I(_0884_),
    .Z(_1895_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3287_ (.I(_0886_),
    .Z(_1896_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _3288_ (.I(net1126),
    .ZN(_1897_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3289_ (.I(_0889_),
    .Z(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3290_ (.I(_0891_),
    .Z(_1899_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3291_ (.I(net1205),
    .ZN(_1900_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _3292_ (.A1(_1897_),
    .A2(_1758_),
    .A3(_1898_),
    .B1(_1899_),
    .B2(_1900_),
    .ZN(_1901_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3293_ (.A1(net1059),
    .A2(_1895_),
    .B1(_1896_),
    .B2(net1072),
    .C(_1901_),
    .ZN(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3294_ (.I(_0896_),
    .Z(_1903_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3295_ (.I(_0898_),
    .Z(_1904_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3296_ (.I(net1020),
    .ZN(_1905_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3297_ (.I(_0901_),
    .Z(_1906_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3298_ (.I(_0102_),
    .Z(_1907_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3299_ (.I(_0904_),
    .Z(_1908_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3300_ (.I(net1005),
    .ZN(_1909_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _3301_ (.A1(_1905_),
    .A2(_1906_),
    .A3(_1907_),
    .B1(_1908_),
    .B2(_1909_),
    .ZN(_1910_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3302_ (.A1(net1099),
    .A2(_1903_),
    .B1(_1904_),
    .B2(net1086),
    .C(_1910_),
    .ZN(_1911_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _3303_ (.A1(_1885_),
    .A2(_1894_),
    .A3(_1902_),
    .A4(_1911_),
    .ZN(_1912_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3304_ (.I(_0910_),
    .Z(_1913_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3305_ (.I(_0912_),
    .Z(_1914_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _3306_ (.A1(net1263),
    .A2(_1913_),
    .B1(_1914_),
    .B2(net966),
    .ZN(_1915_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3307_ (.I(_0915_),
    .Z(_1916_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3308_ (.I(_0917_),
    .Z(_1917_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3309_ (.A1(net1445),
    .A2(_1916_),
    .B1(_1917_),
    .B2(net992),
    .ZN(_1918_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3310_ (.I(_0920_),
    .Z(_1919_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3311_ (.I(_0922_),
    .Z(_1920_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _3312_ (.A1(net1499),
    .A2(_1919_),
    .B1(_1920_),
    .B2(net1486),
    .ZN(_1921_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3313_ (.I(_0925_),
    .Z(_1922_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3314_ (.I(_0927_),
    .Z(_1923_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _3315_ (.A1(net1459),
    .A2(_1922_),
    .B1(_1923_),
    .B2(net1472),
    .ZN(_1924_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _3316_ (.A1(_1915_),
    .A2(_1918_),
    .A3(_1921_),
    .A4(_1924_),
    .ZN(_1925_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3317_ (.I(_0931_),
    .Z(_1926_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3318_ (.I(_0933_),
    .Z(_1927_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3319_ (.A1(net1179),
    .A2(_1926_),
    .B1(_1927_),
    .B2(net1512),
    .ZN(_1928_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3320_ (.I(_0936_),
    .Z(_1929_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3321_ (.I(_0938_),
    .Z(_1930_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _3322_ (.A1(net1654),
    .A2(_1929_),
    .B1(_1930_),
    .B2(net1130),
    .ZN(_1931_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3323_ (.I(_0941_),
    .Z(_1932_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3324_ (.I(_0943_),
    .Z(_1933_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3325_ (.A1(net1192),
    .A2(_1932_),
    .B1(_1933_),
    .B2(net1112),
    .ZN(_1934_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3326_ (.I(_0946_),
    .Z(_1935_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3327_ (.A1(net1166),
    .A2(_1935_),
    .B(_1775_),
    .ZN(_1936_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _3328_ (.A1(_1928_),
    .A2(_1931_),
    .A3(_1934_),
    .A4(_1936_),
    .ZN(_1937_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _3329_ (.A1(_1912_),
    .A2(_1925_),
    .A3(_1937_),
    .ZN(_1938_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3330_ (.I(_0951_),
    .Z(_1939_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3331_ (.I(_0953_),
    .Z(_1940_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3332_ (.I(net1605),
    .ZN(_1941_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3333_ (.I(_0956_),
    .Z(_1942_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3334_ (.I(_0958_),
    .Z(_1943_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3335_ (.I(_0960_),
    .Z(_1944_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3336_ (.A1(net1632),
    .A2(_1943_),
    .A3(_1944_),
    .ZN(_1945_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3337_ (.A1(_1941_),
    .A2(_1942_),
    .B(_1945_),
    .ZN(_1946_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3338_ (.A1(net1619),
    .A2(_1939_),
    .B1(_1940_),
    .B2(net1552),
    .C(_1946_),
    .ZN(_1947_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3339_ (.I(_0965_),
    .Z(_1948_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3340_ (.I(_0967_),
    .Z(_1949_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _3341_ (.I(net1286),
    .ZN(_1950_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3342_ (.I(_0970_),
    .Z(_1951_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3343_ (.I(_0972_),
    .Z(_1952_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3344_ (.I(net1592),
    .ZN(_1953_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _3345_ (.A1(_1950_),
    .A2(_1951_),
    .A3(_1784_),
    .B1(_1952_),
    .B2(_1953_),
    .ZN(_1954_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3346_ (.A1(net1566),
    .A2(_1948_),
    .B1(_1949_),
    .B2(net1579),
    .C(_1954_),
    .ZN(_1955_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3347_ (.I(_0977_),
    .Z(_1956_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3348_ (.I(_0979_),
    .Z(_1957_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3349_ (.I(net1046),
    .ZN(_1958_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3350_ (.I(_0982_),
    .Z(_1959_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3351_ (.I(_0984_),
    .Z(_1960_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_8 _3352_ (.I(net1538),
    .ZN(_1961_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _3353_ (.A1(_1958_),
    .A2(_1959_),
    .B1(_1960_),
    .B2(_1961_),
    .ZN(_1962_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3354_ (.A1(net1033),
    .A2(_1956_),
    .B1(_1957_),
    .B2(net1640),
    .C(_1962_),
    .ZN(_1963_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3355_ (.I(_0989_),
    .Z(_1964_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3356_ (.I(_0991_),
    .Z(_1965_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3357_ (.I(net996),
    .ZN(_1966_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3358_ (.I(_0994_),
    .Z(_1967_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3359_ (.I(_0996_),
    .Z(_1968_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3360_ (.I(net1396),
    .ZN(_1969_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _3361_ (.A1(_1966_),
    .A2(_1967_),
    .B1(_1968_),
    .B2(_1969_),
    .ZN(_1970_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3362_ (.A1(net1529),
    .A2(_1964_),
    .B1(_1965_),
    .B2(net1525),
    .C(_1970_),
    .ZN(_1971_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3363_ (.A1(net1764),
    .A2(net1763),
    .A3(_1963_),
    .A4(net1762),
    .ZN(_1972_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3364_ (.I(_1002_),
    .Z(_1973_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3365_ (.I(_1004_),
    .Z(_1974_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _3366_ (.A1(net1405),
    .A2(_1973_),
    .B1(_1974_),
    .B2(net1419),
    .ZN(_1975_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3367_ (.I(_1007_),
    .Z(_1976_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3368_ (.I(_1009_),
    .Z(_1977_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3369_ (.A1(net1432),
    .A2(_1976_),
    .B1(_1977_),
    .B2(net1338),
    .ZN(_1978_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3370_ (.I(_1012_),
    .Z(_1979_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _3371_ (.I(_1014_),
    .Z(_1980_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3372_ (.A1(net1353),
    .A2(_1979_),
    .B1(_1980_),
    .B2(net1366),
    .ZN(_1981_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3373_ (.I(_1017_),
    .Z(_1982_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3374_ (.I(_1019_),
    .Z(_1983_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3375_ (.A1(net1233),
    .A2(_1982_),
    .B1(_1983_),
    .B2(net1379),
    .ZN(_1984_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _3376_ (.A1(_1975_),
    .A2(_1978_),
    .A3(_1981_),
    .A4(_1984_),
    .ZN(_1985_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3377_ (.I(_1023_),
    .Z(_1986_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3378_ (.I(_1025_),
    .Z(_1987_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3379_ (.A1(net1139),
    .A2(_1986_),
    .B1(_1987_),
    .B2(net926),
    .ZN(_1988_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3380_ (.I(_1028_),
    .Z(_1989_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3381_ (.I(_1030_),
    .Z(_1990_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3382_ (.A1(net1153),
    .A2(_1989_),
    .B1(_1990_),
    .B2(net939),
    .ZN(_1991_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3383_ (.I(_1033_),
    .Z(_1992_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3384_ (.I(_1035_),
    .Z(_1993_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3385_ (.A1(net900),
    .A2(_1992_),
    .B1(_1993_),
    .B2(net913),
    .ZN(_1994_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3386_ (.I(_1038_),
    .Z(_1995_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3387_ (.I(_1040_),
    .Z(_1996_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _3388_ (.A1(net953),
    .A2(_1995_),
    .B1(_1996_),
    .B2(net979),
    .ZN(_1997_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _3389_ (.A1(_1988_),
    .A2(_1991_),
    .A3(_1994_),
    .A4(_1997_),
    .ZN(_1998_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3390_ (.A1(_1972_),
    .A2(_1985_),
    .A3(_1998_),
    .ZN(_1999_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3391_ (.A1(_1869_),
    .A2(_1870_),
    .B1(_1938_),
    .B2(_1999_),
    .ZN(_2331_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3392_ (.I(net1642),
    .ZN(_2000_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3393_ (.I(net1313),
    .ZN(_2001_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3394_ (.A1(_2001_),
    .A2(_1872_),
    .A3(_1873_),
    .ZN(_2002_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _3395_ (.A1(net1326),
    .A2(_1875_),
    .A3(_1876_),
    .Z(_2003_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3396_ (.I(net1393),
    .ZN(_2004_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _3397_ (.A1(_2004_),
    .A2(_1879_),
    .A3(_1748_),
    .ZN(_2005_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3398_ (.I(net1300),
    .ZN(_2006_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3399_ (.A1(_2006_),
    .A2(_1882_),
    .A3(_1883_),
    .ZN(_2007_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _3400_ (.A1(_2002_),
    .A2(_2003_),
    .A3(_2005_),
    .A4(_2007_),
    .ZN(_2008_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3401_ (.I(net1273),
    .ZN(_2009_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3402_ (.I(net1260),
    .ZN(_2010_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _3403_ (.A1(_2009_),
    .A2(_1889_),
    .A3(_1890_),
    .B1(_1891_),
    .B2(_2010_),
    .ZN(_2011_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3404_ (.A1(net1220),
    .A2(_1886_),
    .B1(_1887_),
    .B2(net1247),
    .C(_2011_),
    .ZN(_2012_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _3405_ (.I(net1127),
    .ZN(_2013_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3406_ (.I(net1206),
    .ZN(_2014_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _3407_ (.A1(_2013_),
    .A2(_1758_),
    .A3(_1898_),
    .B1(_1899_),
    .B2(_2014_),
    .ZN(_2015_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3408_ (.A1(net1060),
    .A2(_1895_),
    .B1(_1896_),
    .B2(net1073),
    .C(_2015_),
    .ZN(_2016_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3409_ (.I(net1021),
    .ZN(_2017_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3410_ (.I(net1006),
    .ZN(_2018_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _3411_ (.A1(_2017_),
    .A2(_1906_),
    .A3(_1907_),
    .B1(_1908_),
    .B2(_2018_),
    .ZN(_2019_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3412_ (.A1(net1100),
    .A2(_1903_),
    .B1(_1904_),
    .B2(net1087),
    .C(_2019_),
    .ZN(_2020_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3413_ (.A1(_2008_),
    .A2(_2012_),
    .A3(_2016_),
    .A4(_2020_),
    .ZN(_2021_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _3414_ (.A1(net1274),
    .A2(_1913_),
    .B1(_1914_),
    .B2(net967),
    .ZN(_2022_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3415_ (.A1(net1446),
    .A2(_1916_),
    .B1(_1917_),
    .B2(net993),
    .ZN(_2023_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _3416_ (.A1(net1500),
    .A2(_1919_),
    .B1(_1920_),
    .B2(net1487),
    .ZN(_2024_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _3417_ (.A1(net1460),
    .A2(_1922_),
    .B1(_1923_),
    .B2(net1473),
    .ZN(_2025_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _3418_ (.A1(_2022_),
    .A2(_2023_),
    .A3(_2024_),
    .A4(_2025_),
    .ZN(_2026_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3419_ (.A1(net1180),
    .A2(_1926_),
    .B1(_1927_),
    .B2(net1513),
    .ZN(_2027_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _3420_ (.A1(net1655),
    .A2(_1929_),
    .B1(_1930_),
    .B2(net1141),
    .ZN(_2028_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3421_ (.A1(net1193),
    .A2(_1932_),
    .B1(_1933_),
    .B2(net1113),
    .ZN(_2029_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3422_ (.A1(net1167),
    .A2(_1935_),
    .B(_1775_),
    .ZN(_2030_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _3423_ (.A1(_2027_),
    .A2(_2028_),
    .A3(_2029_),
    .A4(_2030_),
    .ZN(_2031_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3424_ (.A1(_2021_),
    .A2(_2026_),
    .A3(_2031_),
    .ZN(_2032_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3425_ (.I(net1606),
    .ZN(_2033_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3426_ (.A1(net1633),
    .A2(_1943_),
    .A3(_1944_),
    .ZN(_2034_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3427_ (.A1(_2033_),
    .A2(_1942_),
    .B(_2034_),
    .ZN(_2035_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3428_ (.A1(net1620),
    .A2(_1939_),
    .B1(_1940_),
    .B2(net1553),
    .C(_2035_),
    .ZN(_2036_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _3429_ (.I(net1287),
    .ZN(_2037_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3430_ (.I(net1593),
    .ZN(_2038_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _3431_ (.A1(_2037_),
    .A2(_1951_),
    .A3(_1784_),
    .B1(_1952_),
    .B2(_2038_),
    .ZN(_2039_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3432_ (.A1(net1567),
    .A2(_1948_),
    .B1(_1949_),
    .B2(net1580),
    .C(_2039_),
    .ZN(_2040_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3433_ (.I(net1047),
    .ZN(_2041_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_8 _3434_ (.I(net1539),
    .ZN(_2042_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _3435_ (.A1(_2041_),
    .A2(_1959_),
    .B1(_1960_),
    .B2(_2042_),
    .ZN(_2043_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3436_ (.A1(net1034),
    .A2(_1956_),
    .B1(_1957_),
    .B2(net1641),
    .C(_2043_),
    .ZN(_2044_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3437_ (.I(net1007),
    .ZN(_2045_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3438_ (.I(net1407),
    .ZN(_2046_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _3439_ (.A1(_2045_),
    .A2(_1967_),
    .B1(_1968_),
    .B2(_2046_),
    .ZN(_2047_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3440_ (.A1(net1540),
    .A2(_1964_),
    .B1(_1965_),
    .B2(net1526),
    .C(_2047_),
    .ZN(_2048_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3441_ (.A1(net1761),
    .A2(net1760),
    .A3(_2044_),
    .A4(net1759),
    .ZN(_2049_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _3442_ (.A1(net1406),
    .A2(_1973_),
    .B1(_1974_),
    .B2(net1420),
    .ZN(_2050_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3443_ (.A1(net1433),
    .A2(_1976_),
    .B1(_1977_),
    .B2(net1339),
    .ZN(_2051_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _3444_ (.A1(net1354),
    .A2(_1979_),
    .B1(_1980_),
    .B2(net1367),
    .ZN(_2052_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3445_ (.A1(net1234),
    .A2(_1982_),
    .B1(_1983_),
    .B2(net1380),
    .ZN(_2053_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _3446_ (.A1(_2050_),
    .A2(_2051_),
    .A3(_2052_),
    .A4(_2053_),
    .ZN(_2054_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3447_ (.A1(net1140),
    .A2(_1986_),
    .B1(_1987_),
    .B2(net927),
    .ZN(_2055_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3448_ (.A1(net1154),
    .A2(_1989_),
    .B1(_1990_),
    .B2(net940),
    .ZN(_2056_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3449_ (.A1(net901),
    .A2(_1992_),
    .B1(_1993_),
    .B2(net914),
    .ZN(_2057_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _3450_ (.A1(net954),
    .A2(_1995_),
    .B1(_1996_),
    .B2(net980),
    .ZN(_2058_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _3451_ (.A1(_2055_),
    .A2(_2056_),
    .A3(_2057_),
    .A4(_2058_),
    .ZN(_2059_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3452_ (.A1(_2049_),
    .A2(_2054_),
    .A3(_2059_),
    .ZN(_2060_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3453_ (.A1(_2000_),
    .A2(_1870_),
    .B1(_2032_),
    .B2(_2060_),
    .ZN(_2332_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3454_ (.I(net1653),
    .ZN(_2061_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3455_ (.I(net1314),
    .ZN(_2062_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3456_ (.A1(_2062_),
    .A2(_1872_),
    .A3(_1873_),
    .ZN(_2063_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _3457_ (.A1(net1327),
    .A2(_1875_),
    .A3(_1876_),
    .Z(_2064_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3458_ (.I(net1394),
    .ZN(_2065_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3459_ (.I(_0028_),
    .Z(_2066_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _3460_ (.A1(_2065_),
    .A2(_1879_),
    .A3(_2066_),
    .ZN(_2067_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3461_ (.I(net1301),
    .ZN(_2068_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3462_ (.A1(_2068_),
    .A2(_1882_),
    .A3(_1883_),
    .ZN(_2069_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _3463_ (.A1(_2063_),
    .A2(_2064_),
    .A3(_2067_),
    .A4(_2069_),
    .ZN(_2070_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3464_ (.I(net1275),
    .ZN(_2071_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3465_ (.I(net1261),
    .ZN(_2072_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _3466_ (.A1(_2071_),
    .A2(_1889_),
    .A3(_1890_),
    .B1(_1891_),
    .B2(_2072_),
    .ZN(_2073_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3467_ (.A1(net1221),
    .A2(_1886_),
    .B1(_1887_),
    .B2(net1248),
    .C(_2073_),
    .ZN(_2074_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _3468_ (.I(net1128),
    .ZN(_2075_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3469_ (.I(_0173_),
    .Z(_2076_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3470_ (.I(net1208),
    .ZN(_2077_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _3471_ (.A1(_2075_),
    .A2(_2076_),
    .A3(_1898_),
    .B1(_1899_),
    .B2(_2077_),
    .ZN(_2078_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3472_ (.A1(net1061),
    .A2(_1895_),
    .B1(_1896_),
    .B2(net1075),
    .C(_2078_),
    .ZN(_2079_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3473_ (.I(net1022),
    .ZN(_2080_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3474_ (.I(net1009),
    .ZN(_2081_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _3475_ (.A1(_2080_),
    .A2(_1906_),
    .A3(_1907_),
    .B1(_1908_),
    .B2(_2081_),
    .ZN(_2082_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3476_ (.A1(net1101),
    .A2(_1903_),
    .B1(_1904_),
    .B2(net1088),
    .C(_2082_),
    .ZN(_2083_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3477_ (.A1(_2070_),
    .A2(_2074_),
    .A3(_2079_),
    .A4(_2083_),
    .ZN(_2084_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _3478_ (.A1(net1285),
    .A2(_1913_),
    .B1(_1914_),
    .B2(net968),
    .ZN(_2085_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3479_ (.A1(net1447),
    .A2(_1916_),
    .B1(_1917_),
    .B2(net994),
    .ZN(_2086_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _3480_ (.A1(net1501),
    .A2(_1919_),
    .B1(_1920_),
    .B2(net1488),
    .ZN(_2087_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _3481_ (.A1(net1461),
    .A2(_1922_),
    .B1(_1923_),
    .B2(net1475),
    .ZN(_2088_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3482_ (.A1(_2085_),
    .A2(_2086_),
    .A3(_2087_),
    .A4(_2088_),
    .ZN(_2089_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3483_ (.A1(net1181),
    .A2(_1926_),
    .B1(_1927_),
    .B2(net1514),
    .ZN(_2090_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _3484_ (.A1(net1656),
    .A2(_1929_),
    .B1(_1930_),
    .B2(net1152),
    .ZN(_2091_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3485_ (.A1(net1194),
    .A2(_1932_),
    .B1(_1933_),
    .B2(net1114),
    .ZN(_2092_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3486_ (.I(_0011_),
    .Z(_2093_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3487_ (.A1(net1168),
    .A2(_1935_),
    .B(_2093_),
    .ZN(_2094_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _3488_ (.A1(_2090_),
    .A2(_2091_),
    .A3(_2092_),
    .A4(_2094_),
    .ZN(_2095_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3489_ (.A1(_2084_),
    .A2(_2089_),
    .A3(_2095_),
    .ZN(_2096_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3490_ (.I(net1608),
    .ZN(_2097_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3491_ (.A1(net1634),
    .A2(_1943_),
    .A3(_1944_),
    .ZN(_2098_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3492_ (.A1(_2097_),
    .A2(_1942_),
    .B(_2098_),
    .ZN(_2099_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3493_ (.A1(net1621),
    .A2(_1939_),
    .B1(_1940_),
    .B2(net1554),
    .C(_2099_),
    .ZN(_2100_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _3494_ (.I(net1288),
    .ZN(_2101_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3495_ (.I(_1147_),
    .Z(_2102_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3496_ (.I(net1594),
    .ZN(_2103_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _3497_ (.A1(_2101_),
    .A2(_1951_),
    .A3(_2102_),
    .B1(_1952_),
    .B2(_2103_),
    .ZN(_2104_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3498_ (.A1(net1568),
    .A2(_1948_),
    .B1(_1949_),
    .B2(net1581),
    .C(_2104_),
    .ZN(_2105_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3499_ (.I(net1048),
    .ZN(_2106_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_8 _3500_ (.I(net1541),
    .ZN(_2107_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _3501_ (.A1(_2106_),
    .A2(_1959_),
    .B1(_1960_),
    .B2(_2107_),
    .ZN(_2108_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3502_ (.A1(net1035),
    .A2(_1956_),
    .B1(_1957_),
    .B2(net1643),
    .C(_2108_),
    .ZN(_2109_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3503_ (.I(net1019),
    .ZN(_2110_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3504_ (.I(net1418),
    .ZN(_2111_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _3505_ (.A1(_2110_),
    .A2(_1967_),
    .B1(_1968_),
    .B2(_2111_),
    .ZN(_2112_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3506_ (.A1(net1551),
    .A2(_1964_),
    .B1(_1965_),
    .B2(net1527),
    .C(_2112_),
    .ZN(_2113_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3507_ (.A1(net1758),
    .A2(net1757),
    .A3(_2109_),
    .A4(net1756),
    .ZN(_2114_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _3508_ (.A1(net1408),
    .A2(_1973_),
    .B1(_1974_),
    .B2(net1421),
    .ZN(_2115_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3509_ (.A1(net1434),
    .A2(_1976_),
    .B1(_1977_),
    .B2(net1342),
    .ZN(_2116_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _3510_ (.A1(net1355),
    .A2(_1979_),
    .B1(_1980_),
    .B2(net1368),
    .ZN(_2117_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3511_ (.A1(net1235),
    .A2(_1982_),
    .B1(_1983_),
    .B2(net1381),
    .ZN(_2118_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _3512_ (.A1(_2115_),
    .A2(_2116_),
    .A3(_2117_),
    .A4(_2118_),
    .ZN(_2119_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3513_ (.A1(net1142),
    .A2(_1986_),
    .B1(_1987_),
    .B2(net928),
    .ZN(_2120_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3514_ (.A1(net1155),
    .A2(_1989_),
    .B1(_1990_),
    .B2(net942),
    .ZN(_2121_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3515_ (.A1(net902),
    .A2(_1992_),
    .B1(_1993_),
    .B2(net915),
    .ZN(_2122_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _3516_ (.A1(net955),
    .A2(_1995_),
    .B1(_1996_),
    .B2(net981),
    .ZN(_2123_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _3517_ (.A1(_2120_),
    .A2(_2121_),
    .A3(_2122_),
    .A4(_2123_),
    .ZN(_2124_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3518_ (.A1(_2114_),
    .A2(_2119_),
    .A3(_2124_),
    .ZN(_2125_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3519_ (.A1(_2061_),
    .A2(_1870_),
    .B1(_2096_),
    .B2(_2125_),
    .ZN(_2333_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3520_ (.I(net1664),
    .ZN(_2126_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3521_ (.I(net1315),
    .ZN(_2127_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3522_ (.A1(_2127_),
    .A2(_1872_),
    .A3(_1873_),
    .ZN(_2128_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _3523_ (.A1(net1328),
    .A2(_1875_),
    .A3(_1876_),
    .Z(_2129_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3524_ (.I(net1395),
    .ZN(_2130_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _3525_ (.A1(_2130_),
    .A2(_1879_),
    .A3(_2066_),
    .ZN(_2131_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3526_ (.I(net1302),
    .ZN(_2132_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _3527_ (.A1(_2132_),
    .A2(_1882_),
    .A3(_1883_),
    .ZN(_2133_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _3528_ (.A1(_2128_),
    .A2(_2129_),
    .A3(_2131_),
    .A4(_2133_),
    .ZN(_2134_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3529_ (.I(net1276),
    .ZN(_2135_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3530_ (.I(net1262),
    .ZN(_2136_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _3531_ (.A1(_2135_),
    .A2(_1889_),
    .A3(_1890_),
    .B1(_1891_),
    .B2(_2136_),
    .ZN(_2137_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3532_ (.A1(net1222),
    .A2(_1886_),
    .B1(_1887_),
    .B2(net1249),
    .C(_2137_),
    .ZN(_2138_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _3533_ (.I(net1129),
    .ZN(_2139_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3534_ (.I(net1209),
    .ZN(_2140_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _3535_ (.A1(_2139_),
    .A2(_2076_),
    .A3(_1898_),
    .B1(_1899_),
    .B2(_2140_),
    .ZN(_2141_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3536_ (.A1(net1062),
    .A2(_1895_),
    .B1(_1896_),
    .B2(net1076),
    .C(_2141_),
    .ZN(_2142_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3537_ (.I(net1023),
    .ZN(_2143_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3538_ (.I(net1010),
    .ZN(_2144_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _3539_ (.A1(_2143_),
    .A2(_1906_),
    .A3(_1907_),
    .B1(_1908_),
    .B2(_2144_),
    .ZN(_2145_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3540_ (.A1(net1102),
    .A2(_1903_),
    .B1(_1904_),
    .B2(net1089),
    .C(_2145_),
    .ZN(_2146_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3541_ (.A1(_2134_),
    .A2(_2138_),
    .A3(_2142_),
    .A4(_2146_),
    .ZN(_2147_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _3542_ (.A1(net1296),
    .A2(_1913_),
    .B1(_1914_),
    .B2(net969),
    .ZN(_2148_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3543_ (.A1(net1448),
    .A2(_1916_),
    .B1(_1917_),
    .B2(net995),
    .ZN(_2149_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _3544_ (.A1(net1502),
    .A2(_1919_),
    .B1(_1920_),
    .B2(net1489),
    .ZN(_2150_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _3545_ (.A1(net1462),
    .A2(_1922_),
    .B1(_1923_),
    .B2(net1476),
    .ZN(_2151_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3546_ (.A1(_2148_),
    .A2(_2149_),
    .A3(_2150_),
    .A4(_2151_),
    .ZN(_2152_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3547_ (.A1(net1182),
    .A2(_1926_),
    .B1(_1927_),
    .B2(net1515),
    .ZN(_2153_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _3548_ (.A1(net1657),
    .A2(_1929_),
    .B1(_1930_),
    .B2(net1163),
    .ZN(_2154_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3549_ (.A1(net1195),
    .A2(_1932_),
    .B1(_1933_),
    .B2(net1115),
    .ZN(_2155_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3550_ (.A1(net1169),
    .A2(_1935_),
    .B(_2093_),
    .ZN(_2156_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _3551_ (.A1(_2153_),
    .A2(_2154_),
    .A3(_2155_),
    .A4(_2156_),
    .ZN(_2157_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3552_ (.A1(_2147_),
    .A2(_2152_),
    .A3(_2157_),
    .ZN(_2158_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3553_ (.I(net1609),
    .ZN(_2159_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3554_ (.A1(net1635),
    .A2(_1943_),
    .A3(_1944_),
    .ZN(_2160_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3555_ (.A1(_2159_),
    .A2(_1942_),
    .B(_2160_),
    .ZN(_2161_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3556_ (.A1(net1622),
    .A2(_1939_),
    .B1(_1940_),
    .B2(net1555),
    .C(_2161_),
    .ZN(_2162_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _3557_ (.I(net1289),
    .ZN(_2163_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3558_ (.I(net1595),
    .ZN(_2164_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _3559_ (.A1(_2163_),
    .A2(_1951_),
    .A3(_2102_),
    .B1(_1952_),
    .B2(_2164_),
    .ZN(_2165_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3560_ (.A1(net1569),
    .A2(_1948_),
    .B1(_1949_),
    .B2(net1582),
    .C(_2165_),
    .ZN(_2166_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3561_ (.I(net1049),
    .ZN(_2167_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_8 _3562_ (.I(net1542),
    .ZN(_2168_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _3563_ (.A1(_2167_),
    .A2(_1959_),
    .B1(_1960_),
    .B2(_2168_),
    .ZN(_2169_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3564_ (.A1(net1036),
    .A2(_1956_),
    .B1(_1957_),
    .B2(net1644),
    .C(_2169_),
    .ZN(_2170_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3565_ (.I(net1030),
    .ZN(_2171_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3566_ (.I(net1429),
    .ZN(_2172_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _3567_ (.A1(_2171_),
    .A2(_1967_),
    .B1(_1968_),
    .B2(_2172_),
    .ZN(_2173_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3568_ (.A1(net1562),
    .A2(_1964_),
    .B1(_1965_),
    .B2(net1528),
    .C(_2173_),
    .ZN(_2174_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3569_ (.A1(net1755),
    .A2(net1754),
    .A3(_2170_),
    .A4(net1753),
    .ZN(_2175_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _3570_ (.A1(net1409),
    .A2(_1973_),
    .B1(_1974_),
    .B2(net1422),
    .ZN(_2176_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3571_ (.A1(net1435),
    .A2(_1976_),
    .B1(_1977_),
    .B2(net1343),
    .ZN(_2177_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _3572_ (.A1(net1356),
    .A2(_1979_),
    .B1(_1980_),
    .B2(net1369),
    .ZN(_2178_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3573_ (.A1(net1236),
    .A2(_1982_),
    .B1(_1983_),
    .B2(net1382),
    .ZN(_2179_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _3574_ (.A1(_2176_),
    .A2(_2177_),
    .A3(_2178_),
    .A4(_2179_),
    .ZN(_2180_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3575_ (.A1(net1143),
    .A2(_1986_),
    .B1(_1987_),
    .B2(net929),
    .ZN(_2181_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3576_ (.A1(net1156),
    .A2(_1989_),
    .B1(_1990_),
    .B2(net943),
    .ZN(_2182_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3577_ (.A1(net903),
    .A2(_1992_),
    .B1(_1993_),
    .B2(net916),
    .ZN(_2183_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _3578_ (.A1(net956),
    .A2(_1995_),
    .B1(_1996_),
    .B2(net982),
    .ZN(_2184_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _3579_ (.A1(_2181_),
    .A2(_2182_),
    .A3(_2183_),
    .A4(_2184_),
    .ZN(_2185_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3580_ (.A1(_2175_),
    .A2(_2180_),
    .A3(_2185_),
    .ZN(_2186_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3581_ (.A1(_2126_),
    .A2(_1870_),
    .B1(_2158_),
    .B2(_2186_),
    .ZN(_2334_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3582_ (.I(net908),
    .ZN(_2187_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3583_ (.I(net1316),
    .ZN(_2188_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3584_ (.A1(_2188_),
    .A2(_0023_),
    .A3(_0238_),
    .ZN(_2189_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3585_ (.A1(net1330),
    .A2(_0033_),
    .A3(_0040_),
    .Z(_2190_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3586_ (.I(net1397),
    .ZN(_2191_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3587_ (.A1(_2191_),
    .A2(_0051_),
    .A3(_2066_),
    .ZN(_2192_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3588_ (.I(net1303),
    .ZN(_2193_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3589_ (.A1(_2193_),
    .A2(_0060_),
    .A3(_0054_),
    .ZN(_2194_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _3590_ (.A1(_2189_),
    .A2(_2190_),
    .A3(_2192_),
    .A4(_2194_),
    .ZN(_2195_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3591_ (.I(net1277),
    .ZN(_2196_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3592_ (.I(net1264),
    .ZN(_2197_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _3593_ (.A1(_2196_),
    .A2(_0077_),
    .A3(_0062_),
    .B1(_0084_),
    .B2(_2197_),
    .ZN(_2198_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3594_ (.A1(net1223),
    .A2(_0068_),
    .B1(_0073_),
    .B2(net1250),
    .C(_2198_),
    .ZN(_2199_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3595_ (.I(net1131),
    .ZN(_2200_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3596_ (.I(net1210),
    .ZN(_2201_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _3597_ (.A1(_2200_),
    .A2(_2076_),
    .A3(_0105_),
    .B1(_0111_),
    .B2(_2201_),
    .ZN(_2202_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3598_ (.A1(net1064),
    .A2(_0092_),
    .B1(_0099_),
    .B2(net1077),
    .C(net1828),
    .ZN(_2203_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3599_ (.I(net1024),
    .ZN(_2204_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3600_ (.I(net1011),
    .ZN(_2205_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _3601_ (.A1(_2204_),
    .A2(_0125_),
    .A3(_0103_),
    .B1(_0130_),
    .B2(_2205_),
    .ZN(_2206_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3602_ (.A1(net1103),
    .A2(_0117_),
    .B1(_0121_),
    .B2(net1090),
    .C(_2206_),
    .ZN(_2207_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3603_ (.A1(_2195_),
    .A2(_2199_),
    .A3(_2203_),
    .A4(_2207_),
    .ZN(_2208_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _3604_ (.A1(net1307),
    .A2(_0138_),
    .B1(_0142_),
    .B2(net970),
    .ZN(_2209_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3605_ (.A1(net1449),
    .A2(_0148_),
    .B1(_0153_),
    .B2(net997),
    .ZN(_2210_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3606_ (.A1(net1503),
    .A2(_0157_),
    .B1(_0162_),
    .B2(net1490),
    .ZN(_2211_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _3607_ (.A1(net1464),
    .A2(_0166_),
    .B1(_0169_),
    .B2(net1477),
    .ZN(_2212_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _3608_ (.A1(net1822),
    .A2(_2210_),
    .A3(_2211_),
    .A4(_2212_),
    .ZN(_2213_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3609_ (.A1(net1183),
    .A2(_0175_),
    .B1(_0178_),
    .B2(net1516),
    .ZN(_2214_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _3610_ (.A1(net1658),
    .A2(_0182_),
    .B1(_0185_),
    .B2(net1174),
    .ZN(_2215_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3611_ (.A1(net1197),
    .A2(_0190_),
    .B1(_0196_),
    .B2(net1116),
    .ZN(_2216_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3612_ (.A1(net1170),
    .A2(_0201_),
    .B(_2093_),
    .ZN(_2217_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3613_ (.A1(_2214_),
    .A2(_2215_),
    .A3(_2216_),
    .A4(_2217_),
    .ZN(_2218_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3614_ (.A1(_2208_),
    .A2(_2213_),
    .A3(_2218_),
    .ZN(_2219_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3615_ (.I(net1610),
    .ZN(_2220_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3616_ (.A1(net1636),
    .A2(_0219_),
    .A3(_0221_),
    .ZN(_2221_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3617_ (.A1(_2220_),
    .A2(_0217_),
    .B(_2221_),
    .ZN(_2222_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3618_ (.A1(net1623),
    .A2(_0209_),
    .B1(_0213_),
    .B2(net1556),
    .C(_2222_),
    .ZN(_2223_));
 gf180mcu_fd_sc_mcu7t5v0__inv_4 _3619_ (.I(net1290),
    .ZN(_2224_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3620_ (.I(net1597),
    .ZN(_2225_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _3621_ (.A1(_2224_),
    .A2(_0235_),
    .A3(_2102_),
    .B1(_0240_),
    .B2(_2225_),
    .ZN(_2226_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3622_ (.A1(net1570),
    .A2(_0228_),
    .B1(_0232_),
    .B2(net1583),
    .C(_2226_),
    .ZN(_2227_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3623_ (.I(net1050),
    .ZN(_2228_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_8 _3624_ (.I(net1543),
    .ZN(_2229_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _3625_ (.A1(_2228_),
    .A2(_0253_),
    .B1(_0256_),
    .B2(_2229_),
    .ZN(_2230_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3626_ (.A1(net1037),
    .A2(_0246_),
    .B1(_0249_),
    .B2(net1645),
    .C(_2230_),
    .ZN(_2231_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _3627_ (.I(net1041),
    .ZN(_2232_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3628_ (.I(net1440),
    .ZN(_2233_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _3629_ (.A1(_2232_),
    .A2(_0269_),
    .B1(_0272_),
    .B2(_2233_),
    .ZN(_2234_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _3630_ (.A1(net1574),
    .A2(_0262_),
    .B1(_0265_),
    .B2(net1530),
    .C(_2234_),
    .ZN(_2235_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3631_ (.A1(net1821),
    .A2(net1820),
    .A3(_2231_),
    .A4(net1819),
    .ZN(_2236_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _3632_ (.A1(net1410),
    .A2(_0279_),
    .B1(_0282_),
    .B2(net1423),
    .ZN(_2237_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3633_ (.A1(net1436),
    .A2(_0286_),
    .B1(_0290_),
    .B2(net1344),
    .ZN(_2238_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3634_ (.A1(net1357),
    .A2(_0295_),
    .B1(_0298_),
    .B2(net1370),
    .ZN(_2239_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3635_ (.A1(net1237),
    .A2(_0302_),
    .B1(_0305_),
    .B2(net1383),
    .ZN(_2240_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _3636_ (.A1(_2237_),
    .A2(_2238_),
    .A3(_2239_),
    .A4(_2240_),
    .ZN(_2241_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3637_ (.A1(net1144),
    .A2(_0310_),
    .B1(_0314_),
    .B2(net931),
    .ZN(_2242_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3638_ (.A1(net1157),
    .A2(_0318_),
    .B1(_0321_),
    .B2(net944),
    .ZN(_2243_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3639_ (.A1(net904),
    .A2(_0325_),
    .B1(_0328_),
    .B2(net917),
    .ZN(_2244_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _3640_ (.A1(net957),
    .A2(_0332_),
    .B1(_0335_),
    .B2(net983),
    .ZN(_2245_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _3641_ (.A1(_2242_),
    .A2(_2243_),
    .A3(_2244_),
    .A4(_2245_),
    .ZN(_2246_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3642_ (.A1(_2236_),
    .A2(_2241_),
    .A3(_2246_),
    .ZN(_2247_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3643_ (.A1(_2187_),
    .A2(_0014_),
    .B1(_2219_),
    .B2(_2247_),
    .ZN(_2324_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3644_ (.I(net919),
    .ZN(_2248_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3645_ (.I(net1317),
    .ZN(_2249_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3646_ (.A1(_2249_),
    .A2(_0023_),
    .A3(_0238_),
    .ZN(_2250_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3647_ (.A1(net1331),
    .A2(_0033_),
    .A3(_0040_),
    .Z(_2251_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3648_ (.I(net1398),
    .ZN(_2252_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3649_ (.A1(_2252_),
    .A2(_0051_),
    .A3(_2066_),
    .ZN(_2253_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3650_ (.I(net1304),
    .ZN(_2254_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3651_ (.A1(_2254_),
    .A2(_0060_),
    .A3(_0054_),
    .ZN(_2255_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _3652_ (.A1(_2250_),
    .A2(_2251_),
    .A3(_2253_),
    .A4(_2255_),
    .ZN(_2256_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3653_ (.I(net1278),
    .ZN(_2257_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3654_ (.I(net1265),
    .ZN(_2258_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _3655_ (.A1(_2257_),
    .A2(_0077_),
    .A3(_0062_),
    .B1(_0084_),
    .B2(_2258_),
    .ZN(_2259_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3656_ (.A1(net1224),
    .A2(_0068_),
    .B1(_0073_),
    .B2(net1251),
    .C(_2259_),
    .ZN(_2260_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3657_ (.I(net1132),
    .ZN(_2261_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3658_ (.I(net1211),
    .ZN(_2262_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _3659_ (.A1(_2261_),
    .A2(_2076_),
    .A3(_0105_),
    .B1(_0111_),
    .B2(_2262_),
    .ZN(_2263_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3660_ (.A1(net1065),
    .A2(_0092_),
    .B1(_0099_),
    .B2(net1078),
    .C(net1827),
    .ZN(_2264_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3661_ (.I(net1025),
    .ZN(_2265_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3662_ (.I(net1012),
    .ZN(_2266_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _3663_ (.A1(_2265_),
    .A2(_0125_),
    .A3(_0103_),
    .B1(_0130_),
    .B2(_2266_),
    .ZN(_2267_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3664_ (.A1(net1104),
    .A2(_0117_),
    .B1(_0121_),
    .B2(net1091),
    .C(_2267_),
    .ZN(_2268_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3665_ (.A1(_2256_),
    .A2(_2260_),
    .A3(_2264_),
    .A4(_2268_),
    .ZN(_2269_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _3666_ (.A1(net1318),
    .A2(_0138_),
    .B1(_0142_),
    .B2(net971),
    .ZN(_2270_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3667_ (.A1(net1450),
    .A2(_0148_),
    .B1(_0153_),
    .B2(net998),
    .ZN(_2271_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3668_ (.A1(net1504),
    .A2(_0157_),
    .B1(_0162_),
    .B2(net1491),
    .ZN(_2272_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _3669_ (.A1(net1465),
    .A2(_0166_),
    .B1(_0169_),
    .B2(net1478),
    .ZN(_2273_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _3670_ (.A1(net1818),
    .A2(_2271_),
    .A3(_2272_),
    .A4(_2273_),
    .ZN(_2274_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3671_ (.A1(net1184),
    .A2(_0175_),
    .B1(_0178_),
    .B2(net1517),
    .ZN(_2275_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _3672_ (.A1(net1659),
    .A2(_0182_),
    .B1(_0185_),
    .B2(net1185),
    .ZN(_2276_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3673_ (.A1(net1198),
    .A2(_0190_),
    .B1(_0196_),
    .B2(net1117),
    .ZN(_2277_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3674_ (.A1(net1171),
    .A2(_0201_),
    .B(_2093_),
    .ZN(_2278_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3675_ (.A1(_2275_),
    .A2(_2276_),
    .A3(_2277_),
    .A4(_2278_),
    .ZN(_2279_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3676_ (.A1(_2269_),
    .A2(_2274_),
    .A3(_2279_),
    .ZN(_2280_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3677_ (.I(net1611),
    .ZN(_2281_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3678_ (.A1(net1637),
    .A2(_0219_),
    .A3(_0221_),
    .ZN(_2282_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3679_ (.A1(_2281_),
    .A2(_0217_),
    .B(_2282_),
    .ZN(_2283_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3680_ (.A1(net1624),
    .A2(_0209_),
    .B1(_0213_),
    .B2(net1557),
    .C(_2283_),
    .ZN(_2284_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _3681_ (.I(net1291),
    .ZN(_2285_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3682_ (.I(net1598),
    .ZN(_2286_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _3683_ (.A1(_2285_),
    .A2(_0235_),
    .A3(_2102_),
    .B1(_0240_),
    .B2(_2286_),
    .ZN(_2287_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3684_ (.A1(net1571),
    .A2(_0228_),
    .B1(_0232_),
    .B2(net1584),
    .C(_2287_),
    .ZN(_2288_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3685_ (.I(net1051),
    .ZN(_2289_));
 gf180mcu_fd_sc_mcu7t5v0__inv_4 _3686_ (.I(net1544),
    .ZN(_2290_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _3687_ (.A1(_2289_),
    .A2(_0253_),
    .B1(_0256_),
    .B2(_2290_),
    .ZN(_2291_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3688_ (.A1(net1038),
    .A2(_0246_),
    .B1(_0249_),
    .B2(net1646),
    .C(_2291_),
    .ZN(_2292_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _3689_ (.I(net1052),
    .ZN(_2293_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3690_ (.I(net1451),
    .ZN(_2294_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _3691_ (.A1(_2293_),
    .A2(_0269_),
    .B1(_0272_),
    .B2(_2294_),
    .ZN(_2295_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3692_ (.A1(net1585),
    .A2(_0262_),
    .B1(_0265_),
    .B2(net1531),
    .C(_2295_),
    .ZN(_2296_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3693_ (.A1(net1817),
    .A2(net1816),
    .A3(_2292_),
    .A4(net1815),
    .ZN(_2297_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _3694_ (.A1(net1411),
    .A2(_0279_),
    .B1(_0282_),
    .B2(net1424),
    .ZN(_2298_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _3695_ (.A1(net1437),
    .A2(_0286_),
    .B1(_0290_),
    .B2(net1345),
    .ZN(_2299_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3696_ (.A1(net1358),
    .A2(_0295_),
    .B1(_0298_),
    .B2(net1371),
    .ZN(_2300_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3697_ (.A1(net1238),
    .A2(_0302_),
    .B1(_0305_),
    .B2(net1384),
    .ZN(_2301_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _3698_ (.A1(_2298_),
    .A2(_2299_),
    .A3(_2300_),
    .A4(_2301_),
    .ZN(_2302_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3699_ (.A1(net1145),
    .A2(_0310_),
    .B1(_0314_),
    .B2(net932),
    .ZN(_2303_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3700_ (.A1(net1158),
    .A2(_0318_),
    .B1(_0321_),
    .B2(net945),
    .ZN(_2304_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3701_ (.A1(net905),
    .A2(_0325_),
    .B1(_0328_),
    .B2(net918),
    .ZN(_2305_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _3702_ (.A1(net958),
    .A2(_0332_),
    .B1(_0335_),
    .B2(net984),
    .ZN(_2306_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _3703_ (.A1(_2303_),
    .A2(_2304_),
    .A3(_2305_),
    .A4(_2306_),
    .ZN(_2307_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3704_ (.A1(_2297_),
    .A2(_2302_),
    .A3(_2307_),
    .ZN(_2308_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3705_ (.A1(_2248_),
    .A2(_0014_),
    .B1(_2280_),
    .B2(_2308_),
    .ZN(_2325_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3706_ (.I(net1),
    .ZN(_0000_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3707_ (.I(net1666),
    .Z(_0001_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3708_ (.A1(net1665),
    .A2(_0001_),
    .ZN(_0002_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3709_ (.I(_0002_),
    .Z(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3710_ (.A1(net1668),
    .A2(net1667),
    .ZN(_0004_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3711_ (.I(_0004_),
    .Z(_0005_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _3712_ (.A1(_0003_),
    .A2(_0005_),
    .ZN(_0006_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _3713_ (.I(net1670),
    .ZN(_0007_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _3714_ (.I(net1669),
    .ZN(_0008_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _3715_ (.A1(_0007_),
    .A2(_0008_),
    .ZN(_0009_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _3716_ (.I(_0009_),
    .Z(_0010_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3717_ (.A1(_0006_),
    .A2(_0010_),
    .ZN(_0011_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3718_ (.I(_0011_),
    .Z(_0012_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3719_ (.I(_0012_),
    .Z(_0013_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3720_ (.I(_0013_),
    .Z(_0014_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _3721_ (.I(_0014_),
    .Z(_0015_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3722_ (.I(net496),
    .ZN(_0016_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3723_ (.I(net1668),
    .ZN(_0017_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3724_ (.I(_0017_),
    .Z(_0018_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3725_ (.I(net1667),
    .Z(_0019_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3726_ (.A1(net1665),
    .A2(_0001_),
    .Z(_0020_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _3727_ (.A1(_0018_),
    .A2(_0019_),
    .A3(_0020_),
    .ZN(_0021_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _3728_ (.I(_0021_),
    .Z(_0022_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3729_ (.I(_0022_),
    .Z(_0023_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3730_ (.I(_0023_),
    .Z(_0024_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3731_ (.A1(net1670),
    .A2(_0008_),
    .ZN(_0025_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3732_ (.I(_0025_),
    .Z(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3733_ (.I(_0026_),
    .Z(_0027_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3734_ (.I(_0027_),
    .Z(_0028_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3735_ (.I(_0028_),
    .Z(_0029_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3736_ (.A1(_0016_),
    .A2(_0024_),
    .A3(_0029_),
    .ZN(_0030_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3737_ (.I(net1669),
    .Z(_0031_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3738_ (.A1(_0007_),
    .A2(_0031_),
    .ZN(_0032_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3739_ (.I(_0032_),
    .Z(_0033_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3740_ (.I(_0033_),
    .Z(_0034_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3741_ (.I(net1668),
    .Z(_0035_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3742_ (.I(net1667),
    .Z(_0036_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _3743_ (.I(_0036_),
    .ZN(_0037_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _3744_ (.I(_0002_),
    .Z(_0038_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3745_ (.A1(_0035_),
    .A2(_0037_),
    .A3(_0038_),
    .Z(_0039_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3746_ (.I(_0039_),
    .Z(_0040_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3747_ (.I(_0040_),
    .Z(_0041_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3748_ (.A1(net512),
    .A2(_0034_),
    .A3(_0041_),
    .Z(_0042_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3749_ (.I(net590),
    .ZN(_0043_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3750_ (.I(net1665),
    .Z(_0044_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3751_ (.I(_0044_),
    .Z(_0045_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _3752_ (.I(net1666),
    .ZN(_0046_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3753_ (.I(_0046_),
    .Z(_0047_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3754_ (.A1(_0035_),
    .A2(_0036_),
    .Z(_0048_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3755_ (.I(_0048_),
    .Z(_0049_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _3756_ (.A1(_0045_),
    .A2(_0047_),
    .A3(_0049_),
    .ZN(_0050_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3757_ (.I(_0050_),
    .Z(_0051_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _3758_ (.I(_0051_),
    .Z(_0052_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3759_ (.I(_0027_),
    .Z(_0053_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3760_ (.I(_0053_),
    .Z(_0054_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _3761_ (.A1(_0043_),
    .A2(_0052_),
    .A3(_0054_),
    .ZN(_0055_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3762_ (.I(net481),
    .ZN(_0056_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _3763_ (.I(_0044_),
    .ZN(_0057_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _3764_ (.I(_0001_),
    .Z(_0058_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _3765_ (.A1(_0018_),
    .A2(_0019_),
    .A3(_0057_),
    .A4(_0058_),
    .ZN(_0059_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3766_ (.I(_0059_),
    .Z(_0060_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _3767_ (.I(_0060_),
    .Z(_0061_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _3768_ (.I(_0027_),
    .Z(_0062_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _3769_ (.I(_0062_),
    .Z(_0063_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _3770_ (.A1(_0056_),
    .A2(_0061_),
    .A3(_0063_),
    .ZN(_0064_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _3771_ (.A1(_0030_),
    .A2(_0042_),
    .A3(_0055_),
    .A4(_0064_),
    .ZN(_0065_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3772_ (.I(_0025_),
    .Z(_0066_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3773_ (.A1(_0006_),
    .A2(_0066_),
    .ZN(_0067_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3774_ (.I(_0067_),
    .Z(_0068_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3775_ (.I(_0068_),
    .Z(_0069_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3776_ (.I(_0004_),
    .Z(_0070_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _3777_ (.A1(_0057_),
    .A2(_0058_),
    .A3(_0070_),
    .ZN(_0071_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3778_ (.A1(_0071_),
    .A2(_0066_),
    .ZN(_0072_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3779_ (.I(_0072_),
    .Z(_0073_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3780_ (.I(_0073_),
    .Z(_0074_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3781_ (.I(net450),
    .ZN(_0075_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _3782_ (.A1(_0018_),
    .A2(_0019_),
    .A3(_0002_),
    .ZN(_0076_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3783_ (.I(_0076_),
    .Z(_0077_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3784_ (.I(_0077_),
    .Z(_0078_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _3785_ (.I(_0026_),
    .Z(_0079_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3786_ (.I(_0079_),
    .Z(_0080_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3787_ (.I(net1670),
    .Z(_0081_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3788_ (.I(_0020_),
    .Z(_0082_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _3789_ (.A1(_0081_),
    .A2(_0008_),
    .A3(_0070_),
    .A4(_0082_),
    .ZN(_0083_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3790_ (.I(_0083_),
    .Z(_0084_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3791_ (.I(_0084_),
    .Z(_0085_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3792_ (.I(net434),
    .ZN(_0086_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _3793_ (.A1(_0075_),
    .A2(_0078_),
    .A3(_0080_),
    .B1(_0085_),
    .B2(_0086_),
    .ZN(_0087_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3794_ (.A1(net387),
    .A2(_0069_),
    .B1(_0074_),
    .B2(net418),
    .C(_0087_),
    .ZN(_0088_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _3795_ (.A1(_0007_),
    .A2(net1669),
    .ZN(_0089_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3796_ (.I(_0089_),
    .Z(_0090_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3797_ (.A1(_0090_),
    .A2(_0076_),
    .ZN(_0091_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _3798_ (.I(_0091_),
    .Z(_0092_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3799_ (.I(_0092_),
    .Z(_0093_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _3800_ (.A1(_0017_),
    .A2(_0036_),
    .A3(_0044_),
    .A4(_0046_),
    .ZN(_0094_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _3801_ (.I(_0094_),
    .Z(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3802_ (.I(_0089_),
    .Z(_0096_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3803_ (.I(_0096_),
    .Z(_0097_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3804_ (.A1(_0095_),
    .A2(_0097_),
    .ZN(_0098_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _3805_ (.I(_0098_),
    .Z(_0099_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3806_ (.I(_0099_),
    .Z(_0100_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3807_ (.I(net279),
    .ZN(_0101_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3808_ (.I(_0096_),
    .Z(_0102_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3809_ (.I(_0102_),
    .Z(_0103_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _3810_ (.A1(_0035_),
    .A2(_0037_),
    .A3(_0044_),
    .A4(_0046_),
    .ZN(_0104_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3811_ (.I(_0104_),
    .Z(_0105_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3812_ (.I(_0105_),
    .Z(_0106_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _3813_ (.I(_0007_),
    .Z(_0107_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _3814_ (.I(_0031_),
    .Z(_0108_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _3815_ (.A1(net1668),
    .A2(_0036_),
    .A3(net1665),
    .A4(_0001_),
    .Z(_0109_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _3816_ (.A1(_0107_),
    .A2(_0108_),
    .A3(_0109_),
    .ZN(_0110_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3817_ (.I(_0110_),
    .Z(_0111_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3818_ (.I(_0111_),
    .Z(_0112_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3819_ (.I(net372),
    .ZN(_0113_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _3820_ (.A1(_0101_),
    .A2(_0103_),
    .A3(_0106_),
    .B1(_0112_),
    .B2(_0113_),
    .ZN(_0114_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3821_ (.A1(net201),
    .A2(_0093_),
    .B1(_0100_),
    .B2(net216),
    .C(_0114_),
    .ZN(_0115_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3822_ (.A1(_0021_),
    .A2(_0090_),
    .ZN(_0116_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3823_ (.I(_0116_),
    .Z(_0117_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3824_ (.I(_0117_),
    .Z(_0118_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _3825_ (.I(_0059_),
    .Z(_0119_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3826_ (.A1(_0090_),
    .A2(_0119_),
    .ZN(_0120_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3827_ (.I(_0120_),
    .Z(_0121_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3828_ (.I(_0121_),
    .Z(_0122_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3829_ (.I(net154),
    .ZN(_0123_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _3830_ (.A1(_0045_),
    .A2(_0047_),
    .A3(_0070_),
    .ZN(_0124_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3831_ (.I(_0124_),
    .Z(_0125_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3832_ (.I(_0125_),
    .Z(_0126_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3833_ (.I(_0090_),
    .Z(_0127_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3834_ (.I(_0127_),
    .Z(_0128_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _3835_ (.A1(_0107_),
    .A2(_0108_),
    .A3(_0038_),
    .A4(_0070_),
    .ZN(_0129_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3836_ (.I(_0129_),
    .Z(_0130_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3837_ (.I(_0130_),
    .Z(_0131_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3838_ (.I(net139),
    .ZN(_0132_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _3839_ (.A1(_0123_),
    .A2(_0126_),
    .A3(_0128_),
    .B1(_0131_),
    .B2(_0132_),
    .ZN(_0133_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3840_ (.A1(net248),
    .A2(_0118_),
    .B1(_0122_),
    .B2(net232),
    .C(_0133_),
    .ZN(_0134_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3841_ (.A1(_0065_),
    .A2(_0088_),
    .A3(_0115_),
    .A4(_0134_),
    .ZN(_0135_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _3842_ (.A1(_0005_),
    .A2(_0082_),
    .ZN(_0136_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3843_ (.A1(_0010_),
    .A2(_0136_),
    .ZN(_0137_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3844_ (.I(_0137_),
    .Z(_0138_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3845_ (.I(_0138_),
    .Z(_0139_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3846_ (.I(_0009_),
    .Z(_0140_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3847_ (.A1(_0140_),
    .A2(_0050_),
    .ZN(_0141_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3848_ (.I(_0141_),
    .Z(_0142_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3849_ (.I(_0142_),
    .Z(_0143_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _3850_ (.A1(net367),
    .A2(_0139_),
    .B1(_0143_),
    .B2(net92),
    .ZN(_0144_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3851_ (.A1(_0081_),
    .A2(net1669),
    .ZN(_0145_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _3852_ (.I(_0145_),
    .Z(_0146_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _3853_ (.A1(_0146_),
    .A2(_0124_),
    .ZN(_0147_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3854_ (.I(_0147_),
    .Z(_0148_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3855_ (.I(_0148_),
    .Z(_0149_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _3856_ (.A1(_0081_),
    .A2(_0031_),
    .ZN(_0150_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3857_ (.I(_0109_),
    .Z(_0151_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3858_ (.A1(_0150_),
    .A2(_0151_),
    .Z(_0152_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3859_ (.I(_0152_),
    .Z(_0153_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3860_ (.I(_0153_),
    .Z(_0154_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3861_ (.A1(net651),
    .A2(_0149_),
    .B1(_0154_),
    .B2(net124),
    .ZN(_0155_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3862_ (.A1(_0146_),
    .A2(_0095_),
    .ZN(_0156_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3863_ (.I(_0156_),
    .Z(_0157_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _3864_ (.I(_0157_),
    .Z(_0158_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _3865_ (.I(_0145_),
    .Z(_0159_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3866_ (.I(_0159_),
    .Z(_0160_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3867_ (.A1(_0160_),
    .A2(_0076_),
    .ZN(_0161_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3868_ (.I(_0161_),
    .Z(_0162_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _3869_ (.I(_0162_),
    .Z(_0163_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3870_ (.A1(net714),
    .A2(_0158_),
    .B1(_0163_),
    .B2(net698),
    .ZN(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3871_ (.A1(_0146_),
    .A2(_0071_),
    .ZN(_0165_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3872_ (.I(_0165_),
    .Z(_0166_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3873_ (.I(_0166_),
    .Z(_0167_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3874_ (.A1(_0136_),
    .A2(_0160_),
    .ZN(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3875_ (.I(_0168_),
    .Z(_0169_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3876_ (.I(_0169_),
    .Z(_0170_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _3877_ (.A1(net668),
    .A2(_0167_),
    .B1(_0170_),
    .B2(net683),
    .ZN(_0171_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _3878_ (.A1(net1752),
    .A2(_0155_),
    .A3(_0164_),
    .A4(_0171_),
    .ZN(_0172_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3879_ (.I(_0096_),
    .Z(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3880_ (.A1(_0050_),
    .A2(_0173_),
    .ZN(_0174_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3881_ (.I(_0174_),
    .Z(_0175_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3882_ (.I(_0175_),
    .Z(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _3883_ (.A1(_0160_),
    .A2(_0119_),
    .ZN(_0177_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3884_ (.I(_0177_),
    .Z(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3885_ (.I(_0178_),
    .Z(_0179_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _3886_ (.A1(net341),
    .A2(_0176_),
    .B1(_0179_),
    .B2(net729),
    .ZN(_0180_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3887_ (.A1(_0140_),
    .A2(_0022_),
    .ZN(_0181_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3888_ (.I(_0181_),
    .Z(_0182_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3889_ (.I(_0182_),
    .Z(_0183_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3890_ (.A1(_0140_),
    .A2(_0071_),
    .ZN(_0184_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3891_ (.I(_0184_),
    .Z(_0185_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3892_ (.I(_0185_),
    .Z(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _3893_ (.A1(net894),
    .A2(_0183_),
    .B1(_0186_),
    .B2(net211),
    .ZN(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _3894_ (.A1(_0057_),
    .A2(_0058_),
    .A3(_0048_),
    .Z(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _3895_ (.A1(_0107_),
    .A2(_0108_),
    .A3(_0188_),
    .Z(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3896_ (.I(_0189_),
    .Z(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3897_ (.I(_0190_),
    .Z(_0191_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3898_ (.I(_0035_),
    .Z(_0192_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3899_ (.I(_0037_),
    .Z(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _3900_ (.A1(_0192_),
    .A2(_0193_),
    .A3(_0003_),
    .ZN(_0194_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3901_ (.A1(_0097_),
    .A2(_0194_),
    .ZN(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3902_ (.I(_0195_),
    .Z(_0196_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3903_ (.I(_0196_),
    .Z(_0197_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3904_ (.A1(net357),
    .A2(_0191_),
    .B1(_0197_),
    .B2(net263),
    .ZN(_0198_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _3905_ (.A1(_0003_),
    .A2(_0049_),
    .ZN(_0199_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3906_ (.A1(_0097_),
    .A2(_0199_),
    .ZN(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3907_ (.I(_0200_),
    .Z(_0201_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3908_ (.I(_0201_),
    .Z(_0202_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3909_ (.A1(net325),
    .A2(_0202_),
    .B(_0013_),
    .ZN(_0203_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _3910_ (.A1(_0180_),
    .A2(_0187_),
    .A3(_0198_),
    .A4(_0203_),
    .ZN(_0204_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _3911_ (.A1(_0135_),
    .A2(_0172_),
    .A3(_0204_),
    .ZN(_0205_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3912_ (.A1(_0081_),
    .A2(_0031_),
    .Z(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3913_ (.I(_0206_),
    .Z(_0207_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3914_ (.A1(_0207_),
    .A2(_0188_),
    .Z(_0208_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3915_ (.I(_0208_),
    .Z(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3916_ (.I(_0209_),
    .Z(_0210_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _3917_ (.I(_0104_),
    .Z(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _3918_ (.A1(_0146_),
    .A2(_0211_),
    .ZN(_0212_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3919_ (.I(_0212_),
    .Z(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3920_ (.I(_0213_),
    .Z(_0214_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3921_ (.I(net838),
    .ZN(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _3922_ (.A1(_0045_),
    .A2(_0047_),
    .A3(_0049_),
    .A4(_0207_),
    .ZN(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3923_ (.I(_0216_),
    .Z(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3924_ (.I(_0217_),
    .Z(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3925_ (.I(_0207_),
    .Z(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3926_ (.I(_0219_),
    .Z(_0220_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3927_ (.I(_0151_),
    .Z(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3928_ (.I(_0221_),
    .Z(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3929_ (.A1(net869),
    .A2(_0220_),
    .A3(_0222_),
    .ZN(_0223_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3930_ (.A1(_0215_),
    .A2(_0218_),
    .B(_0223_),
    .ZN(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3931_ (.A1(net853),
    .A2(_0210_),
    .B1(_0214_),
    .B2(net775),
    .C(_0224_),
    .ZN(_0225_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _3932_ (.A1(_0192_),
    .A2(_0193_),
    .A3(_0057_),
    .A4(_0058_),
    .ZN(_0226_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _3933_ (.A1(_0159_),
    .A2(_0226_),
    .ZN(_0227_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3934_ (.I(_0227_),
    .Z(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3935_ (.I(_0228_),
    .Z(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _3936_ (.A1(_0192_),
    .A2(_0193_),
    .A3(_0082_),
    .ZN(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _3937_ (.A1(_0159_),
    .A2(_0230_),
    .ZN(_0231_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3938_ (.I(_0231_),
    .Z(_0232_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3939_ (.I(_0232_),
    .Z(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _3940_ (.I(net465),
    .ZN(_0234_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _3941_ (.I(_0094_),
    .Z(_0235_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _3942_ (.I(_0235_),
    .Z(_0236_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3943_ (.I(_0066_),
    .Z(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3944_ (.I(_0237_),
    .Z(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3945_ (.A1(_0003_),
    .A2(_0049_),
    .A3(_0206_),
    .ZN(_0239_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _3946_ (.I(_0239_),
    .Z(_0240_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _3947_ (.I(_0240_),
    .Z(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3948_ (.I(net823),
    .ZN(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _3949_ (.A1(_0234_),
    .A2(_0236_),
    .A3(_0238_),
    .B1(_0241_),
    .B2(_0242_),
    .ZN(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3950_ (.A1(net792),
    .A2(_0229_),
    .B1(_0233_),
    .B2(net807),
    .C(_0243_),
    .ZN(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3951_ (.A1(_0071_),
    .A2(_0097_),
    .ZN(_0245_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3952_ (.I(_0245_),
    .Z(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3953_ (.I(_0246_),
    .Z(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3954_ (.A1(_0010_),
    .A2(_0119_),
    .ZN(_0248_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _3955_ (.I(_0248_),
    .Z(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3956_ (.I(_0249_),
    .Z(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3957_ (.I(net185),
    .ZN(_0251_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _3958_ (.A1(_0107_),
    .A2(_0108_),
    .A3(_0005_),
    .A4(_0082_),
    .ZN(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3959_ (.I(_0252_),
    .Z(_0253_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3960_ (.I(_0253_),
    .Z(_0254_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _3961_ (.A1(_0192_),
    .A2(_0193_),
    .A3(_0038_),
    .A4(_0206_),
    .ZN(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3962_ (.I(_0255_),
    .Z(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3963_ (.I(_0256_),
    .Z(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_8 _3964_ (.I(net760),
    .ZN(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _3965_ (.A1(_0251_),
    .A2(_0254_),
    .B1(_0257_),
    .B2(_0258_),
    .ZN(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3966_ (.A1(net170),
    .A2(_0247_),
    .B1(_0250_),
    .B2(net833),
    .C(_0259_),
    .ZN(_0260_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3967_ (.A1(_0010_),
    .A2(_0095_),
    .ZN(_0261_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3968_ (.I(_0261_),
    .Z(_0262_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _3969_ (.I(_0262_),
    .Z(_0263_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _3970_ (.A1(_0159_),
    .A2(_0022_),
    .ZN(_0264_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3971_ (.I(_0264_),
    .Z(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _3972_ (.I(_0265_),
    .Z(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3973_ (.I(net56),
    .ZN(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _3974_ (.A1(_0045_),
    .A2(_0047_),
    .A3(_0005_),
    .A4(_0150_),
    .ZN(_0268_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3975_ (.I(_0268_),
    .Z(_0269_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3976_ (.I(_0269_),
    .Z(_0270_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _3977_ (.A1(_0018_),
    .A2(_0019_),
    .A3(_0038_),
    .A4(_0150_),
    .ZN(_0271_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3978_ (.I(_0271_),
    .Z(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3979_ (.I(_0272_),
    .Z(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3980_ (.I(net522),
    .ZN(_0274_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _3981_ (.A1(_0267_),
    .A2(_0270_),
    .B1(_0273_),
    .B2(_0274_),
    .ZN(_0275_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3982_ (.A1(net678),
    .A2(_0263_),
    .B1(_0266_),
    .B2(net745),
    .C(_0275_),
    .ZN(_0276_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _3983_ (.A1(net1750),
    .A2(net1748),
    .A3(_0260_),
    .A4(net1747),
    .ZN(_0277_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3984_ (.A1(_0188_),
    .A2(_0032_),
    .Z(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _3985_ (.I(_0278_),
    .Z(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3986_ (.I(_0279_),
    .Z(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3987_ (.A1(_0151_),
    .A2(_0032_),
    .Z(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _3988_ (.I(_0281_),
    .Z(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3989_ (.I(_0282_),
    .Z(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _3990_ (.A1(net605),
    .A2(_0280_),
    .B1(_0283_),
    .B2(net620),
    .ZN(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3991_ (.A1(_0006_),
    .A2(_0160_),
    .ZN(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3992_ (.I(_0285_),
    .Z(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3993_ (.I(_0286_),
    .Z(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _3994_ (.I(_0026_),
    .Z(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3995_ (.A1(_0288_),
    .A2(_0211_),
    .ZN(_0289_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3996_ (.I(_0289_),
    .Z(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3997_ (.I(_0290_),
    .Z(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3998_ (.A1(net636),
    .A2(_0287_),
    .B1(_0291_),
    .B2(net527),
    .ZN(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3999_ (.I(_0026_),
    .Z(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4000_ (.A1(_0293_),
    .A2(_0226_),
    .ZN(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4001_ (.I(_0294_),
    .Z(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4002_ (.I(_0295_),
    .Z(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4003_ (.A1(_0293_),
    .A2(_0230_),
    .ZN(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4004_ (.I(_0297_),
    .Z(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4005_ (.I(_0298_),
    .Z(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4006_ (.A1(net542),
    .A2(_0296_),
    .B1(_0299_),
    .B2(net559),
    .ZN(_0300_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4007_ (.A1(_0124_),
    .A2(_0293_),
    .ZN(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4008_ (.I(_0301_),
    .Z(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4009_ (.I(_0302_),
    .Z(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4010_ (.A1(_0199_),
    .A2(_0288_),
    .ZN(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4011_ (.I(_0304_),
    .Z(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4012_ (.I(_0305_),
    .Z(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4013_ (.A1(net403),
    .A2(_0303_),
    .B1(_0306_),
    .B2(net574),
    .ZN(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _4014_ (.A1(_0284_),
    .A2(_0292_),
    .A3(_0300_),
    .A4(_0307_),
    .ZN(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4015_ (.A1(_0173_),
    .A2(_0226_),
    .ZN(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4016_ (.I(_0309_),
    .Z(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4017_ (.I(_0310_),
    .Z(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4018_ (.I(_0009_),
    .Z(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4019_ (.A1(_0312_),
    .A2(_0226_),
    .ZN(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4020_ (.I(_0313_),
    .Z(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4021_ (.I(_0314_),
    .Z(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4022_ (.A1(net294),
    .A2(_0311_),
    .B1(_0315_),
    .B2(net46),
    .ZN(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4023_ (.A1(_0173_),
    .A2(_0230_),
    .ZN(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4024_ (.I(_0317_),
    .Z(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4025_ (.I(_0318_),
    .Z(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4026_ (.A1(_0312_),
    .A2(_0230_),
    .ZN(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4027_ (.I(_0320_),
    .Z(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4028_ (.I(_0321_),
    .Z(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4029_ (.A1(net309),
    .A2(_0319_),
    .B1(_0322_),
    .B2(net61),
    .ZN(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4030_ (.A1(_0140_),
    .A2(_0194_),
    .ZN(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4031_ (.I(_0324_),
    .Z(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4032_ (.I(_0325_),
    .Z(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4033_ (.A1(_0312_),
    .A2(_0211_),
    .ZN(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4034_ (.I(_0327_),
    .Z(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4035_ (.I(_0328_),
    .Z(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4036_ (.A1(net15),
    .A2(_0326_),
    .B1(_0329_),
    .B2(net30),
    .ZN(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4037_ (.A1(_0312_),
    .A2(_0199_),
    .ZN(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4038_ (.I(_0331_),
    .Z(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4039_ (.I(_0332_),
    .Z(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _4040_ (.A1(_0150_),
    .A2(_0188_),
    .Z(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4041_ (.I(_0334_),
    .Z(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4042_ (.I(_0335_),
    .Z(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4043_ (.A1(net76),
    .A2(_0333_),
    .B1(_0336_),
    .B2(net107),
    .ZN(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _4044_ (.A1(_0316_),
    .A2(_0323_),
    .A3(_0330_),
    .A4(_0337_),
    .ZN(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _4045_ (.A1(_0277_),
    .A2(_0308_),
    .A3(_0338_),
    .ZN(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4046_ (.A1(_0000_),
    .A2(_0015_),
    .B1(_0205_),
    .B2(_0339_),
    .ZN(_2309_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4047_ (.I(net112),
    .ZN(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4048_ (.I(net497),
    .ZN(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4049_ (.A1(_0341_),
    .A2(_0024_),
    .A3(_0029_),
    .ZN(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4050_ (.A1(net513),
    .A2(_0034_),
    .A3(_0041_),
    .Z(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4051_ (.I(net591),
    .ZN(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _4052_ (.A1(_0344_),
    .A2(_0052_),
    .A3(_0054_),
    .ZN(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4053_ (.I(net482),
    .ZN(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4054_ (.A1(_0346_),
    .A2(_0061_),
    .A3(_0063_),
    .ZN(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _4055_ (.A1(_0342_),
    .A2(_0343_),
    .A3(_0345_),
    .A4(_0347_),
    .ZN(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4056_ (.I(net451),
    .ZN(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4057_ (.I(net435),
    .ZN(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _4058_ (.A1(_0349_),
    .A2(_0078_),
    .A3(_0080_),
    .B1(_0085_),
    .B2(_0350_),
    .ZN(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _4059_ (.A1(net388),
    .A2(_0069_),
    .B1(_0074_),
    .B2(net419),
    .C(_0351_),
    .ZN(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4060_ (.I(net280),
    .ZN(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4061_ (.I(net373),
    .ZN(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _4062_ (.A1(_0353_),
    .A2(_0103_),
    .A3(_0106_),
    .B1(_0112_),
    .B2(_0354_),
    .ZN(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _4063_ (.A1(net202),
    .A2(_0093_),
    .B1(_0100_),
    .B2(net217),
    .C(_0355_),
    .ZN(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4064_ (.I(net155),
    .ZN(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4065_ (.I(net140),
    .ZN(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _4066_ (.A1(_0357_),
    .A2(_0126_),
    .A3(_0128_),
    .B1(_0131_),
    .B2(_0358_),
    .ZN(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _4067_ (.A1(net249),
    .A2(_0118_),
    .B1(_0122_),
    .B2(net233),
    .C(_0359_),
    .ZN(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4068_ (.A1(_0348_),
    .A2(_0352_),
    .A3(_0356_),
    .A4(_0360_),
    .ZN(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4069_ (.A1(net378),
    .A2(_0139_),
    .B1(_0143_),
    .B2(net93),
    .ZN(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4070_ (.A1(net652),
    .A2(_0149_),
    .B1(_0154_),
    .B2(net125),
    .ZN(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4071_ (.A1(net715),
    .A2(_0158_),
    .B1(_0163_),
    .B2(net699),
    .ZN(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4072_ (.A1(net669),
    .A2(_0167_),
    .B1(_0170_),
    .B2(net684),
    .ZN(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _4073_ (.A1(net1746),
    .A2(_0363_),
    .A3(_0364_),
    .A4(_0365_),
    .ZN(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4074_ (.A1(net342),
    .A2(_0176_),
    .B1(_0179_),
    .B2(net730),
    .ZN(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4075_ (.A1(net895),
    .A2(_0183_),
    .B1(_0186_),
    .B2(net222),
    .ZN(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4076_ (.A1(net358),
    .A2(_0191_),
    .B1(_0197_),
    .B2(net264),
    .ZN(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4077_ (.A1(net326),
    .A2(_0202_),
    .B(_0013_),
    .ZN(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4078_ (.A1(_0367_),
    .A2(_0368_),
    .A3(_0369_),
    .A4(_0370_),
    .ZN(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4079_ (.A1(_0361_),
    .A2(_0366_),
    .A3(_0371_),
    .ZN(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4080_ (.I(net839),
    .ZN(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4081_ (.A1(net870),
    .A2(_0220_),
    .A3(_0222_),
    .ZN(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4082_ (.A1(_0373_),
    .A2(_0218_),
    .B(_0374_),
    .ZN(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _4083_ (.A1(net854),
    .A2(_0210_),
    .B1(_0214_),
    .B2(net776),
    .C(_0375_),
    .ZN(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _4084_ (.I(net466),
    .ZN(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4085_ (.I(net824),
    .ZN(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _4086_ (.A1(_0377_),
    .A2(_0236_),
    .A3(_0238_),
    .B1(_0241_),
    .B2(_0378_),
    .ZN(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _4087_ (.A1(net793),
    .A2(_0229_),
    .B1(_0233_),
    .B2(net808),
    .C(_0379_),
    .ZN(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4088_ (.I(net186),
    .ZN(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_8 _4089_ (.I(net761),
    .ZN(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _4090_ (.A1(_0381_),
    .A2(_0254_),
    .B1(_0257_),
    .B2(_0382_),
    .ZN(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _4091_ (.A1(net171),
    .A2(_0247_),
    .B1(_0250_),
    .B2(net844),
    .C(_0383_),
    .ZN(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4092_ (.I(net67),
    .ZN(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4093_ (.I(net533),
    .ZN(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _4094_ (.A1(_0385_),
    .A2(_0270_),
    .B1(_0273_),
    .B2(_0386_),
    .ZN(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _4095_ (.A1(net689),
    .A2(_0263_),
    .B1(_0266_),
    .B2(net746),
    .C(_0387_),
    .ZN(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _4096_ (.A1(net1744),
    .A2(net1742),
    .A3(_0384_),
    .A4(net1741),
    .ZN(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4097_ (.A1(net606),
    .A2(_0280_),
    .B1(_0283_),
    .B2(net621),
    .ZN(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4098_ (.A1(net637),
    .A2(_0287_),
    .B1(_0291_),
    .B2(net528),
    .ZN(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4099_ (.A1(net543),
    .A2(_0296_),
    .B1(_0299_),
    .B2(net560),
    .ZN(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4100_ (.A1(net404),
    .A2(_0303_),
    .B1(_0306_),
    .B2(net575),
    .ZN(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _4101_ (.A1(_0390_),
    .A2(_0391_),
    .A3(_0392_),
    .A4(_0393_),
    .ZN(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4102_ (.A1(net295),
    .A2(_0311_),
    .B1(_0315_),
    .B2(net47),
    .ZN(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4103_ (.A1(net310),
    .A2(_0319_),
    .B1(_0322_),
    .B2(net62),
    .ZN(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4104_ (.A1(net16),
    .A2(_0326_),
    .B1(_0329_),
    .B2(net31),
    .ZN(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4105_ (.A1(net77),
    .A2(_0333_),
    .B1(_0336_),
    .B2(net108),
    .ZN(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _4106_ (.A1(_0395_),
    .A2(_0396_),
    .A3(_0397_),
    .A4(_0398_),
    .ZN(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _4107_ (.A1(_0389_),
    .A2(_0394_),
    .A3(_0399_),
    .ZN(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4108_ (.A1(_0340_),
    .A2(_0015_),
    .B1(net1703),
    .B2(_0400_),
    .ZN(_2314_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4109_ (.I(net223),
    .ZN(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4110_ (.I(net498),
    .ZN(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4111_ (.A1(_0402_),
    .A2(_0024_),
    .A3(_0029_),
    .ZN(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4112_ (.A1(net514),
    .A2(_0034_),
    .A3(_0041_),
    .Z(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4113_ (.I(net592),
    .ZN(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4114_ (.I(_0053_),
    .Z(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _4115_ (.A1(_0405_),
    .A2(_0052_),
    .A3(_0406_),
    .ZN(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4116_ (.I(net483),
    .ZN(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _4117_ (.A1(_0408_),
    .A2(_0061_),
    .A3(_0063_),
    .ZN(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _4118_ (.A1(_0403_),
    .A2(_0404_),
    .A3(_0407_),
    .A4(_0409_),
    .ZN(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4119_ (.I(net452),
    .ZN(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4120_ (.I(net436),
    .ZN(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _4121_ (.A1(_0411_),
    .A2(_0078_),
    .A3(_0080_),
    .B1(_0085_),
    .B2(_0412_),
    .ZN(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _4122_ (.A1(net390),
    .A2(_0069_),
    .B1(_0074_),
    .B2(net420),
    .C(_0413_),
    .ZN(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4123_ (.I(net281),
    .ZN(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4124_ (.I(_0102_),
    .Z(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4125_ (.I(net374),
    .ZN(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _4126_ (.A1(_0415_),
    .A2(_0416_),
    .A3(_0106_),
    .B1(_0112_),
    .B2(_0417_),
    .ZN(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _4127_ (.A1(net203),
    .A2(_0093_),
    .B1(_0100_),
    .B2(net218),
    .C(_0418_),
    .ZN(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4128_ (.I(net157),
    .ZN(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4129_ (.I(net141),
    .ZN(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _4130_ (.A1(_0420_),
    .A2(_0126_),
    .A3(_0128_),
    .B1(_0131_),
    .B2(_0421_),
    .ZN(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _4131_ (.A1(net250),
    .A2(_0118_),
    .B1(_0122_),
    .B2(net235),
    .C(_0422_),
    .ZN(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4132_ (.A1(_0410_),
    .A2(_0414_),
    .A3(_0419_),
    .A4(_0423_),
    .ZN(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4133_ (.A1(net389),
    .A2(_0139_),
    .B1(_0143_),
    .B2(net94),
    .ZN(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4134_ (.A1(net653),
    .A2(_0149_),
    .B1(_0154_),
    .B2(net126),
    .ZN(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4135_ (.A1(net716),
    .A2(_0158_),
    .B1(_0163_),
    .B2(net701),
    .ZN(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4136_ (.A1(net670),
    .A2(_0167_),
    .B1(_0170_),
    .B2(net685),
    .ZN(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _4137_ (.A1(net1740),
    .A2(_0426_),
    .A3(_0427_),
    .A4(_0428_),
    .ZN(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4138_ (.A1(net343),
    .A2(_0176_),
    .B1(_0179_),
    .B2(net731),
    .ZN(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4139_ (.A1(net2),
    .A2(_0183_),
    .B1(_0186_),
    .B2(net234),
    .ZN(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4140_ (.A1(net359),
    .A2(_0191_),
    .B1(_0197_),
    .B2(net265),
    .ZN(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4141_ (.I(_0012_),
    .Z(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4142_ (.A1(net327),
    .A2(_0202_),
    .B(_0433_),
    .ZN(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4143_ (.A1(_0430_),
    .A2(_0431_),
    .A3(_0432_),
    .A4(_0434_),
    .ZN(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4144_ (.A1(_0424_),
    .A2(_0429_),
    .A3(_0435_),
    .ZN(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4145_ (.I(net840),
    .ZN(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4146_ (.A1(net871),
    .A2(_0220_),
    .A3(_0222_),
    .ZN(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4147_ (.A1(_0437_),
    .A2(_0218_),
    .B(_0438_),
    .ZN(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _4148_ (.A1(net856),
    .A2(_0210_),
    .B1(_0214_),
    .B2(net779),
    .C(_0439_),
    .ZN(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _4149_ (.I(net468),
    .ZN(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4150_ (.I(_0237_),
    .Z(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4151_ (.I(net825),
    .ZN(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _4152_ (.A1(_0441_),
    .A2(_0236_),
    .A3(_0442_),
    .B1(_0241_),
    .B2(_0443_),
    .ZN(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _4153_ (.A1(net794),
    .A2(_0229_),
    .B1(_0233_),
    .B2(net809),
    .C(_0444_),
    .ZN(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4154_ (.I(net187),
    .ZN(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_8 _4155_ (.I(net762),
    .ZN(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _4156_ (.A1(_0446_),
    .A2(_0254_),
    .B1(_0257_),
    .B2(_0447_),
    .ZN(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _4157_ (.A1(net172),
    .A2(_0247_),
    .B1(_0250_),
    .B2(net855),
    .C(_0448_),
    .ZN(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4158_ (.I(net78),
    .ZN(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4159_ (.I(net544),
    .ZN(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _4160_ (.A1(_0450_),
    .A2(_0270_),
    .B1(_0273_),
    .B2(_0451_),
    .ZN(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _4161_ (.A1(net700),
    .A2(_0263_),
    .B1(_0266_),
    .B2(net747),
    .C(_0452_),
    .ZN(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _4162_ (.A1(net1738),
    .A2(net1736),
    .A3(_0449_),
    .A4(net1735),
    .ZN(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4163_ (.A1(net607),
    .A2(_0280_),
    .B1(_0283_),
    .B2(net623),
    .ZN(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4164_ (.A1(net638),
    .A2(_0287_),
    .B1(_0291_),
    .B2(net529),
    .ZN(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4165_ (.A1(net545),
    .A2(_0296_),
    .B1(_0299_),
    .B2(net561),
    .ZN(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4166_ (.A1(net405),
    .A2(_0303_),
    .B1(_0306_),
    .B2(net576),
    .ZN(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _4167_ (.A1(_0455_),
    .A2(_0456_),
    .A3(_0457_),
    .A4(_0458_),
    .ZN(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4168_ (.A1(net296),
    .A2(_0311_),
    .B1(_0315_),
    .B2(net48),
    .ZN(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4169_ (.A1(net312),
    .A2(_0319_),
    .B1(_0322_),
    .B2(net63),
    .ZN(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4170_ (.A1(net17),
    .A2(_0326_),
    .B1(_0329_),
    .B2(net32),
    .ZN(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4171_ (.A1(net79),
    .A2(_0333_),
    .B1(_0336_),
    .B2(net109),
    .ZN(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _4172_ (.A1(_0460_),
    .A2(_0461_),
    .A3(_0462_),
    .A4(_0463_),
    .ZN(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _4173_ (.A1(_0454_),
    .A2(_0459_),
    .A3(_0464_),
    .ZN(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4174_ (.A1(_0401_),
    .A2(_0015_),
    .B1(net1702),
    .B2(_0465_),
    .ZN(_2315_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4175_ (.I(net334),
    .ZN(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4176_ (.I(net499),
    .ZN(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4177_ (.A1(_0467_),
    .A2(_0024_),
    .A3(_0029_),
    .ZN(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4178_ (.A1(net515),
    .A2(_0034_),
    .A3(_0041_),
    .Z(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4179_ (.I(net593),
    .ZN(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _4180_ (.A1(_0470_),
    .A2(_0052_),
    .A3(_0406_),
    .ZN(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4181_ (.I(net484),
    .ZN(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _4182_ (.A1(_0472_),
    .A2(_0061_),
    .A3(_0063_),
    .ZN(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _4183_ (.A1(_0468_),
    .A2(_0469_),
    .A3(_0471_),
    .A4(_0473_),
    .ZN(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4184_ (.I(net453),
    .ZN(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4185_ (.I(net437),
    .ZN(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _4186_ (.A1(_0475_),
    .A2(_0078_),
    .A3(_0080_),
    .B1(_0085_),
    .B2(_0476_),
    .ZN(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _4187_ (.A1(net391),
    .A2(_0069_),
    .B1(_0074_),
    .B2(net421),
    .C(_0477_),
    .ZN(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4188_ (.I(net282),
    .ZN(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4189_ (.I(net375),
    .ZN(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _4190_ (.A1(_0479_),
    .A2(_0416_),
    .A3(_0106_),
    .B1(_0112_),
    .B2(_0480_),
    .ZN(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _4191_ (.A1(net204),
    .A2(_0093_),
    .B1(_0100_),
    .B2(net219),
    .C(_0481_),
    .ZN(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4192_ (.I(net158),
    .ZN(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4193_ (.I(net142),
    .ZN(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _4194_ (.A1(_0483_),
    .A2(_0126_),
    .A3(_0128_),
    .B1(_0131_),
    .B2(_0484_),
    .ZN(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _4195_ (.A1(net251),
    .A2(_0118_),
    .B1(_0122_),
    .B2(net236),
    .C(_0485_),
    .ZN(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4196_ (.A1(_0474_),
    .A2(_0478_),
    .A3(_0482_),
    .A4(_0486_),
    .ZN(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4197_ (.A1(net400),
    .A2(_0139_),
    .B1(_0143_),
    .B2(net95),
    .ZN(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4198_ (.A1(net654),
    .A2(_0149_),
    .B1(_0154_),
    .B2(net127),
    .ZN(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4199_ (.A1(net717),
    .A2(_0158_),
    .B1(_0163_),
    .B2(net702),
    .ZN(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4200_ (.A1(net671),
    .A2(_0167_),
    .B1(_0170_),
    .B2(net686),
    .ZN(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _4201_ (.A1(net1734),
    .A2(_0489_),
    .A3(_0490_),
    .A4(_0491_),
    .ZN(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4202_ (.A1(net344),
    .A2(_0176_),
    .B1(_0179_),
    .B2(net732),
    .ZN(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4203_ (.A1(net3),
    .A2(_0183_),
    .B1(_0186_),
    .B2(net245),
    .ZN(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4204_ (.A1(net360),
    .A2(_0191_),
    .B1(_0197_),
    .B2(net266),
    .ZN(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4205_ (.A1(net328),
    .A2(_0202_),
    .B(_0433_),
    .ZN(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4206_ (.A1(_0493_),
    .A2(_0494_),
    .A3(_0495_),
    .A4(_0496_),
    .ZN(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4207_ (.A1(_0487_),
    .A2(_0492_),
    .A3(_0497_),
    .ZN(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4208_ (.I(net841),
    .ZN(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4209_ (.A1(net872),
    .A2(_0220_),
    .A3(_0222_),
    .ZN(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4210_ (.A1(_0499_),
    .A2(_0218_),
    .B(_0500_),
    .ZN(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _4211_ (.A1(net857),
    .A2(_0210_),
    .B1(_0214_),
    .B2(net780),
    .C(_0501_),
    .ZN(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _4212_ (.I(net469),
    .ZN(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4213_ (.I(net826),
    .ZN(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _4214_ (.A1(_0503_),
    .A2(_0236_),
    .A3(_0442_),
    .B1(_0241_),
    .B2(_0504_),
    .ZN(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _4215_ (.A1(net795),
    .A2(_0229_),
    .B1(_0233_),
    .B2(net810),
    .C(_0505_),
    .ZN(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4216_ (.I(net188),
    .ZN(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_8 _4217_ (.I(net763),
    .ZN(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _4218_ (.A1(_0507_),
    .A2(_0254_),
    .B1(_0257_),
    .B2(_0508_),
    .ZN(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _4219_ (.A1(net173),
    .A2(_0247_),
    .B1(_0250_),
    .B2(net866),
    .C(_0509_),
    .ZN(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4220_ (.I(net89),
    .ZN(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4221_ (.I(net555),
    .ZN(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _4222_ (.A1(_0511_),
    .A2(_0270_),
    .B1(_0273_),
    .B2(_0512_),
    .ZN(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _4223_ (.A1(net711),
    .A2(_0263_),
    .B1(_0266_),
    .B2(net748),
    .C(_0513_),
    .ZN(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _4224_ (.A1(net1732),
    .A2(net1730),
    .A3(_0510_),
    .A4(net1729),
    .ZN(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4225_ (.A1(net608),
    .A2(_0280_),
    .B1(_0283_),
    .B2(net624),
    .ZN(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4226_ (.A1(net639),
    .A2(_0287_),
    .B1(_0291_),
    .B2(net530),
    .ZN(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4227_ (.A1(net546),
    .A2(_0296_),
    .B1(_0299_),
    .B2(net562),
    .ZN(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4228_ (.A1(net406),
    .A2(_0303_),
    .B1(_0306_),
    .B2(net577),
    .ZN(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _4229_ (.A1(_0516_),
    .A2(_0517_),
    .A3(_0518_),
    .A4(_0519_),
    .ZN(_0520_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4230_ (.A1(net297),
    .A2(_0311_),
    .B1(_0315_),
    .B2(net49),
    .ZN(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4231_ (.A1(net313),
    .A2(_0319_),
    .B1(_0322_),
    .B2(net64),
    .ZN(_0522_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4232_ (.A1(net18),
    .A2(_0326_),
    .B1(_0329_),
    .B2(net33),
    .ZN(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4233_ (.A1(net80),
    .A2(_0333_),
    .B1(_0336_),
    .B2(net110),
    .ZN(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _4234_ (.A1(_0521_),
    .A2(_0522_),
    .A3(_0523_),
    .A4(_0524_),
    .ZN(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _4235_ (.A1(_0515_),
    .A2(_0520_),
    .A3(_0525_),
    .ZN(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4236_ (.A1(_0466_),
    .A2(_0015_),
    .B1(net1701),
    .B2(_0526_),
    .ZN(_2316_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4237_ (.I(net445),
    .ZN(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4238_ (.I(_0014_),
    .Z(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4239_ (.I(net501),
    .ZN(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4240_ (.I(_0023_),
    .Z(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4241_ (.I(_0027_),
    .Z(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4242_ (.I(_0531_),
    .Z(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4243_ (.A1(_0529_),
    .A2(_0530_),
    .A3(_0532_),
    .ZN(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4244_ (.I(_0033_),
    .Z(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4245_ (.I(_0040_),
    .Z(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4246_ (.A1(net516),
    .A2(_0534_),
    .A3(_0535_),
    .Z(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4247_ (.I(net594),
    .ZN(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4248_ (.I(_0051_),
    .Z(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4249_ (.A1(_0537_),
    .A2(_0538_),
    .A3(_0406_),
    .ZN(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4250_ (.I(net485),
    .ZN(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4251_ (.I(_0060_),
    .Z(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4252_ (.I(_0062_),
    .Z(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4253_ (.A1(_0540_),
    .A2(_0541_),
    .A3(_0542_),
    .ZN(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _4254_ (.A1(_0533_),
    .A2(_0536_),
    .A3(_0539_),
    .A4(_0543_),
    .ZN(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4255_ (.I(_0068_),
    .Z(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4256_ (.I(_0073_),
    .Z(_0546_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4257_ (.I(net454),
    .ZN(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4258_ (.I(_0077_),
    .Z(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4259_ (.I(_0079_),
    .Z(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4260_ (.I(_0084_),
    .Z(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4261_ (.I(net438),
    .ZN(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _4262_ (.A1(_0547_),
    .A2(_0548_),
    .A3(_0549_),
    .B1(_0550_),
    .B2(_0551_),
    .ZN(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _4263_ (.A1(net392),
    .A2(_0545_),
    .B1(_0546_),
    .B2(net423),
    .C(_0552_),
    .ZN(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4264_ (.I(_0092_),
    .Z(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4265_ (.I(_0099_),
    .Z(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4266_ (.I(net283),
    .ZN(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4267_ (.I(_0105_),
    .Z(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4268_ (.I(_0111_),
    .Z(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4269_ (.I(net376),
    .ZN(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _4270_ (.A1(_0556_),
    .A2(_0416_),
    .A3(_0557_),
    .B1(_0558_),
    .B2(_0559_),
    .ZN(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _4271_ (.A1(net205),
    .A2(_0554_),
    .B1(_0555_),
    .B2(net220),
    .C(net1826),
    .ZN(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4272_ (.I(_0117_),
    .Z(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4273_ (.I(_0121_),
    .Z(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4274_ (.I(net159),
    .ZN(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4275_ (.I(_0125_),
    .Z(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4276_ (.I(_0127_),
    .Z(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4277_ (.I(_0130_),
    .Z(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4278_ (.I(net143),
    .ZN(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _4279_ (.A1(_0564_),
    .A2(_0565_),
    .A3(_0566_),
    .B1(_0567_),
    .B2(_0568_),
    .ZN(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _4280_ (.A1(net252),
    .A2(_0562_),
    .B1(_0563_),
    .B2(net237),
    .C(_0569_),
    .ZN(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _4281_ (.A1(_0544_),
    .A2(_0553_),
    .A3(_0561_),
    .A4(_0570_),
    .ZN(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4282_ (.I(_0138_),
    .Z(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4283_ (.I(_0142_),
    .Z(_0573_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4284_ (.A1(net411),
    .A2(_0572_),
    .B1(_0573_),
    .B2(net96),
    .ZN(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4285_ (.I(_0148_),
    .Z(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4286_ (.I(_0153_),
    .Z(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4287_ (.A1(net656),
    .A2(_0575_),
    .B1(_0576_),
    .B2(net128),
    .ZN(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4288_ (.I(_0157_),
    .Z(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4289_ (.I(_0162_),
    .Z(_0579_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4290_ (.A1(net718),
    .A2(_0578_),
    .B1(_0579_),
    .B2(net703),
    .ZN(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4291_ (.I(_0166_),
    .Z(_0581_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4292_ (.I(_0169_),
    .Z(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4293_ (.A1(net672),
    .A2(_0581_),
    .B1(_0582_),
    .B2(net687),
    .ZN(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _4294_ (.A1(net1728),
    .A2(_0577_),
    .A3(_0580_),
    .A4(_0583_),
    .ZN(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4295_ (.I(_0175_),
    .Z(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4296_ (.I(_0178_),
    .Z(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4297_ (.A1(net346),
    .A2(_0585_),
    .B1(_0586_),
    .B2(net734),
    .ZN(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4298_ (.I(_0182_),
    .Z(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4299_ (.I(_0185_),
    .Z(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4300_ (.A1(net4),
    .A2(_0588_),
    .B1(_0589_),
    .B2(net256),
    .ZN(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4301_ (.I(_0190_),
    .Z(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4302_ (.I(_0196_),
    .Z(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4303_ (.A1(net361),
    .A2(_0591_),
    .B1(_0592_),
    .B2(net268),
    .ZN(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4304_ (.I(_0201_),
    .Z(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4305_ (.A1(net329),
    .A2(_0594_),
    .B(_0433_),
    .ZN(_0595_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _4306_ (.A1(_0587_),
    .A2(_0590_),
    .A3(_0593_),
    .A4(_0595_),
    .ZN(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4307_ (.A1(_0571_),
    .A2(_0584_),
    .A3(_0596_),
    .ZN(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4308_ (.I(_0209_),
    .Z(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4309_ (.I(_0213_),
    .Z(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4310_ (.I(net842),
    .ZN(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4311_ (.I(_0217_),
    .Z(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4312_ (.I(_0219_),
    .Z(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4313_ (.I(_0221_),
    .Z(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4314_ (.A1(net873),
    .A2(_0602_),
    .A3(_0603_),
    .ZN(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4315_ (.A1(_0600_),
    .A2(_0601_),
    .B(_0604_),
    .ZN(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _4316_ (.A1(net858),
    .A2(_0598_),
    .B1(_0599_),
    .B2(net781),
    .C(_0605_),
    .ZN(_0606_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4317_ (.I(_0228_),
    .Z(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4318_ (.I(_0232_),
    .Z(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__inv_4 _4319_ (.I(net470),
    .ZN(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4320_ (.I(_0235_),
    .Z(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4321_ (.I(_0240_),
    .Z(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4322_ (.I(net827),
    .ZN(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _4323_ (.A1(_0609_),
    .A2(_0610_),
    .A3(_0442_),
    .B1(_0611_),
    .B2(_0612_),
    .ZN(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _4324_ (.A1(net796),
    .A2(_0607_),
    .B1(_0608_),
    .B2(net812),
    .C(_0613_),
    .ZN(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4325_ (.I(_0246_),
    .Z(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4326_ (.I(_0249_),
    .Z(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4327_ (.I(net190),
    .ZN(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4328_ (.I(_0253_),
    .Z(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4329_ (.I(_0256_),
    .Z(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_8 _4330_ (.I(net764),
    .ZN(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _4331_ (.A1(_0617_),
    .A2(_0618_),
    .B1(_0619_),
    .B2(_0620_),
    .ZN(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _4332_ (.A1(net174),
    .A2(_0615_),
    .B1(_0616_),
    .B2(net877),
    .C(_0621_),
    .ZN(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4333_ (.I(_0262_),
    .Z(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4334_ (.I(_0265_),
    .Z(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4335_ (.I(net100),
    .ZN(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4336_ (.I(_0269_),
    .Z(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4337_ (.I(_0272_),
    .Z(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4338_ (.I(net567),
    .ZN(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _4339_ (.A1(_0625_),
    .A2(_0626_),
    .B1(_0627_),
    .B2(_0628_),
    .ZN(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _4340_ (.A1(net722),
    .A2(_0623_),
    .B1(_0624_),
    .B2(net749),
    .C(_0629_),
    .ZN(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _4341_ (.A1(net1726),
    .A2(net1724),
    .A3(_0622_),
    .A4(net1723),
    .ZN(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4342_ (.I(_0279_),
    .Z(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4343_ (.I(_0282_),
    .Z(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4344_ (.A1(net609),
    .A2(_0632_),
    .B1(_0633_),
    .B2(net625),
    .ZN(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4345_ (.I(_0286_),
    .Z(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4346_ (.I(_0290_),
    .Z(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4347_ (.A1(net640),
    .A2(_0635_),
    .B1(_0636_),
    .B2(net531),
    .ZN(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4348_ (.I(_0295_),
    .Z(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4349_ (.I(_0298_),
    .Z(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4350_ (.A1(net547),
    .A2(_0638_),
    .B1(_0639_),
    .B2(net563),
    .ZN(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4351_ (.I(_0302_),
    .Z(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4352_ (.I(_0305_),
    .Z(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4353_ (.A1(net407),
    .A2(_0641_),
    .B1(_0642_),
    .B2(net579),
    .ZN(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _4354_ (.A1(_0634_),
    .A2(_0637_),
    .A3(_0640_),
    .A4(_0643_),
    .ZN(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4355_ (.I(_0310_),
    .Z(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4356_ (.I(_0314_),
    .Z(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4357_ (.A1(net298),
    .A2(_0645_),
    .B1(_0646_),
    .B2(net50),
    .ZN(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4358_ (.I(_0318_),
    .Z(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4359_ (.I(_0321_),
    .Z(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4360_ (.A1(net314),
    .A2(_0648_),
    .B1(_0649_),
    .B2(net65),
    .ZN(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4361_ (.I(_0325_),
    .Z(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4362_ (.I(_0328_),
    .Z(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4363_ (.A1(net19),
    .A2(_0651_),
    .B1(_0652_),
    .B2(net35),
    .ZN(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4364_ (.I(_0332_),
    .Z(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4365_ (.I(_0335_),
    .Z(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4366_ (.A1(net81),
    .A2(_0654_),
    .B1(_0655_),
    .B2(net113),
    .ZN(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _4367_ (.A1(_0647_),
    .A2(_0650_),
    .A3(_0653_),
    .A4(_0656_),
    .ZN(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _4368_ (.A1(_0631_),
    .A2(_0644_),
    .A3(_0657_),
    .ZN(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4369_ (.A1(_0527_),
    .A2(_0528_),
    .B1(net1700),
    .B2(_0658_),
    .ZN(_2317_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4370_ (.I(net556),
    .ZN(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4371_ (.I(net502),
    .ZN(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4372_ (.A1(_0660_),
    .A2(_0530_),
    .A3(_0532_),
    .ZN(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4373_ (.A1(net517),
    .A2(_0534_),
    .A3(_0535_),
    .Z(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4374_ (.I(net595),
    .ZN(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _4375_ (.A1(_0663_),
    .A2(_0538_),
    .A3(_0406_),
    .ZN(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4376_ (.I(net486),
    .ZN(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4377_ (.A1(_0665_),
    .A2(_0541_),
    .A3(_0542_),
    .ZN(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _4378_ (.A1(_0661_),
    .A2(_0662_),
    .A3(_0664_),
    .A4(_0666_),
    .ZN(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4379_ (.I(net455),
    .ZN(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4380_ (.I(net439),
    .ZN(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _4381_ (.A1(_0668_),
    .A2(_0548_),
    .A3(_0549_),
    .B1(_0550_),
    .B2(_0669_),
    .ZN(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _4382_ (.A1(net393),
    .A2(_0545_),
    .B1(_0546_),
    .B2(net424),
    .C(_0670_),
    .ZN(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4383_ (.I(net284),
    .ZN(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4384_ (.I(net377),
    .ZN(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _4385_ (.A1(_0672_),
    .A2(_0416_),
    .A3(_0557_),
    .B1(_0558_),
    .B2(_0673_),
    .ZN(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _4386_ (.A1(net206),
    .A2(_0554_),
    .B1(_0555_),
    .B2(net221),
    .C(net1825),
    .ZN(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4387_ (.I(net160),
    .ZN(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4388_ (.I(net144),
    .ZN(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _4389_ (.A1(_0676_),
    .A2(_0565_),
    .A3(_0566_),
    .B1(_0567_),
    .B2(_0677_),
    .ZN(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _4390_ (.A1(net253),
    .A2(_0562_),
    .B1(_0563_),
    .B2(net238),
    .C(_0678_),
    .ZN(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4391_ (.A1(_0667_),
    .A2(_0671_),
    .A3(_0675_),
    .A4(_0679_),
    .ZN(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4392_ (.A1(net422),
    .A2(_0572_),
    .B1(_0573_),
    .B2(net97),
    .ZN(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4393_ (.A1(net657),
    .A2(_0575_),
    .B1(_0576_),
    .B2(net129),
    .ZN(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4394_ (.A1(net719),
    .A2(_0578_),
    .B1(_0579_),
    .B2(net704),
    .ZN(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4395_ (.A1(net673),
    .A2(_0581_),
    .B1(_0582_),
    .B2(net688),
    .ZN(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _4396_ (.A1(net1722),
    .A2(_0682_),
    .A3(_0683_),
    .A4(_0684_),
    .ZN(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4397_ (.A1(net347),
    .A2(_0585_),
    .B1(_0586_),
    .B2(net735),
    .ZN(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4398_ (.A1(net5),
    .A2(_0588_),
    .B1(_0589_),
    .B2(net267),
    .ZN(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4399_ (.A1(net362),
    .A2(_0591_),
    .B1(_0592_),
    .B2(net269),
    .ZN(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4400_ (.A1(net330),
    .A2(_0594_),
    .B(_0433_),
    .ZN(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _4401_ (.A1(_0686_),
    .A2(_0687_),
    .A3(_0688_),
    .A4(_0689_),
    .ZN(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4402_ (.A1(_0680_),
    .A2(_0685_),
    .A3(_0690_),
    .ZN(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4403_ (.I(net843),
    .ZN(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4404_ (.A1(net874),
    .A2(_0602_),
    .A3(_0603_),
    .ZN(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4405_ (.A1(_0692_),
    .A2(_0601_),
    .B(_0693_),
    .ZN(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _4406_ (.A1(net859),
    .A2(_0598_),
    .B1(_0599_),
    .B2(net782),
    .C(_0694_),
    .ZN(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__inv_4 _4407_ (.I(net471),
    .ZN(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4408_ (.I(net828),
    .ZN(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _4409_ (.A1(_0696_),
    .A2(_0610_),
    .A3(_0442_),
    .B1(_0611_),
    .B2(_0697_),
    .ZN(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _4410_ (.A1(net797),
    .A2(_0607_),
    .B1(_0608_),
    .B2(net813),
    .C(_0698_),
    .ZN(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4411_ (.I(net191),
    .ZN(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_8 _4412_ (.I(net765),
    .ZN(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _4413_ (.A1(_0700_),
    .A2(_0618_),
    .B1(_0619_),
    .B2(_0701_),
    .ZN(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _4414_ (.A1(net175),
    .A2(_0615_),
    .B1(_0616_),
    .B2(net884),
    .C(_0702_),
    .ZN(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4415_ (.I(net111),
    .ZN(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4416_ (.I(net578),
    .ZN(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _4417_ (.A1(_0704_),
    .A2(_0626_),
    .B1(_0627_),
    .B2(_0705_),
    .ZN(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _4418_ (.A1(net733),
    .A2(_0623_),
    .B1(_0624_),
    .B2(net750),
    .C(_0706_),
    .ZN(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _4419_ (.A1(net1720),
    .A2(net1718),
    .A3(_0703_),
    .A4(net1717),
    .ZN(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4420_ (.A1(net610),
    .A2(_0632_),
    .B1(_0633_),
    .B2(net626),
    .ZN(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4421_ (.A1(net641),
    .A2(_0635_),
    .B1(_0636_),
    .B2(net532),
    .ZN(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4422_ (.A1(net548),
    .A2(_0638_),
    .B1(_0639_),
    .B2(net564),
    .ZN(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4423_ (.A1(net408),
    .A2(_0641_),
    .B1(_0642_),
    .B2(net580),
    .ZN(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _4424_ (.A1(_0709_),
    .A2(_0710_),
    .A3(_0711_),
    .A4(_0712_),
    .ZN(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4425_ (.A1(net299),
    .A2(_0645_),
    .B1(_0646_),
    .B2(net51),
    .ZN(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4426_ (.A1(net315),
    .A2(_0648_),
    .B1(_0649_),
    .B2(net66),
    .ZN(_0715_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4427_ (.A1(net20),
    .A2(_0651_),
    .B1(_0652_),
    .B2(net36),
    .ZN(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4428_ (.A1(net82),
    .A2(_0654_),
    .B1(_0655_),
    .B2(net114),
    .ZN(_0717_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _4429_ (.A1(_0714_),
    .A2(_0715_),
    .A3(_0716_),
    .A4(_0717_),
    .ZN(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _4430_ (.A1(_0708_),
    .A2(_0713_),
    .A3(_0718_),
    .ZN(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4431_ (.A1(_0659_),
    .A2(_0528_),
    .B1(net1699),
    .B2(_0719_),
    .ZN(_2318_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4432_ (.I(net667),
    .ZN(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4433_ (.I(net503),
    .ZN(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4434_ (.A1(_0721_),
    .A2(_0530_),
    .A3(_0532_),
    .ZN(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4435_ (.A1(net518),
    .A2(_0534_),
    .A3(_0535_),
    .Z(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4436_ (.I(net596),
    .ZN(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4437_ (.I(_0053_),
    .Z(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4438_ (.A1(_0724_),
    .A2(_0538_),
    .A3(_0725_),
    .ZN(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4439_ (.I(net487),
    .ZN(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4440_ (.A1(_0727_),
    .A2(_0541_),
    .A3(_0542_),
    .ZN(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _4441_ (.A1(_0722_),
    .A2(_0723_),
    .A3(_0726_),
    .A4(_0728_),
    .ZN(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4442_ (.I(net457),
    .ZN(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4443_ (.I(net440),
    .ZN(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _4444_ (.A1(_0730_),
    .A2(_0548_),
    .A3(_0549_),
    .B1(_0550_),
    .B2(_0731_),
    .ZN(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _4445_ (.A1(net394),
    .A2(_0545_),
    .B1(_0546_),
    .B2(net425),
    .C(_0732_),
    .ZN(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4446_ (.I(net285),
    .ZN(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4447_ (.I(_0096_),
    .Z(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4448_ (.I(_0735_),
    .Z(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4449_ (.I(net379),
    .ZN(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _4450_ (.A1(_0734_),
    .A2(_0736_),
    .A3(_0557_),
    .B1(_0558_),
    .B2(_0737_),
    .ZN(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _4451_ (.A1(net207),
    .A2(_0554_),
    .B1(_0555_),
    .B2(net224),
    .C(net1824),
    .ZN(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4452_ (.I(net161),
    .ZN(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4453_ (.I(net146),
    .ZN(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _4454_ (.A1(_0740_),
    .A2(_0565_),
    .A3(_0566_),
    .B1(_0567_),
    .B2(_0741_),
    .ZN(_0742_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _4455_ (.A1(net254),
    .A2(_0562_),
    .B1(_0563_),
    .B2(net239),
    .C(_0742_),
    .ZN(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4456_ (.A1(_0729_),
    .A2(_0733_),
    .A3(_0739_),
    .A4(_0743_),
    .ZN(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4457_ (.A1(net433),
    .A2(_0572_),
    .B1(_0573_),
    .B2(net98),
    .ZN(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4458_ (.A1(net658),
    .A2(_0575_),
    .B1(_0576_),
    .B2(net130),
    .ZN(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4459_ (.A1(net720),
    .A2(_0578_),
    .B1(_0579_),
    .B2(net705),
    .ZN(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4460_ (.A1(net674),
    .A2(_0581_),
    .B1(_0582_),
    .B2(net690),
    .ZN(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _4461_ (.A1(net1716),
    .A2(_0746_),
    .A3(_0747_),
    .A4(_0748_),
    .ZN(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4462_ (.A1(net348),
    .A2(_0585_),
    .B1(_0586_),
    .B2(net736),
    .ZN(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4463_ (.A1(net6),
    .A2(_0588_),
    .B1(_0589_),
    .B2(net278),
    .ZN(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4464_ (.A1(net363),
    .A2(_0591_),
    .B1(_0592_),
    .B2(net270),
    .ZN(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4465_ (.I(_0012_),
    .Z(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4466_ (.A1(net331),
    .A2(_0594_),
    .B(_0753_),
    .ZN(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _4467_ (.A1(_0750_),
    .A2(_0751_),
    .A3(_0752_),
    .A4(_0754_),
    .ZN(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4468_ (.A1(_0744_),
    .A2(_0749_),
    .A3(_0755_),
    .ZN(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4469_ (.I(net845),
    .ZN(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4470_ (.A1(net875),
    .A2(_0602_),
    .A3(_0603_),
    .ZN(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4471_ (.A1(_0757_),
    .A2(_0601_),
    .B(_0758_),
    .ZN(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _4472_ (.A1(net860),
    .A2(_0598_),
    .B1(_0599_),
    .B2(net783),
    .C(_0759_),
    .ZN(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _4473_ (.I(net472),
    .ZN(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4474_ (.I(_0237_),
    .Z(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4475_ (.I(net829),
    .ZN(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _4476_ (.A1(_0761_),
    .A2(_0610_),
    .A3(_0762_),
    .B1(_0611_),
    .B2(_0763_),
    .ZN(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _4477_ (.A1(net798),
    .A2(_0607_),
    .B1(_0608_),
    .B2(net814),
    .C(_0764_),
    .ZN(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4478_ (.I(net192),
    .ZN(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_8 _4479_ (.I(net767),
    .ZN(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _4480_ (.A1(_0766_),
    .A2(_0618_),
    .B1(_0619_),
    .B2(_0767_),
    .ZN(_0768_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _4481_ (.A1(net176),
    .A2(_0615_),
    .B1(_0616_),
    .B2(net886),
    .C(_0768_),
    .ZN(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4482_ (.I(net123),
    .ZN(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4483_ (.I(net589),
    .ZN(_0771_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _4484_ (.A1(_0770_),
    .A2(_0626_),
    .B1(_0627_),
    .B2(_0771_),
    .ZN(_0772_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _4485_ (.A1(net744),
    .A2(_0623_),
    .B1(_0624_),
    .B2(net751),
    .C(_0772_),
    .ZN(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _4486_ (.A1(net1714),
    .A2(net1712),
    .A3(_0769_),
    .A4(net1711),
    .ZN(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4487_ (.A1(net612),
    .A2(_0632_),
    .B1(_0633_),
    .B2(net627),
    .ZN(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4488_ (.A1(net642),
    .A2(_0635_),
    .B1(_0636_),
    .B2(net534),
    .ZN(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4489_ (.A1(net549),
    .A2(_0638_),
    .B1(_0639_),
    .B2(net565),
    .ZN(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4490_ (.A1(net409),
    .A2(_0641_),
    .B1(_0642_),
    .B2(net581),
    .ZN(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _4491_ (.A1(_0775_),
    .A2(_0776_),
    .A3(_0777_),
    .A4(_0778_),
    .ZN(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4492_ (.A1(net301),
    .A2(_0645_),
    .B1(_0646_),
    .B2(net52),
    .ZN(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4493_ (.A1(net316),
    .A2(_0648_),
    .B1(_0649_),
    .B2(net68),
    .ZN(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4494_ (.A1(net21),
    .A2(_0651_),
    .B1(_0652_),
    .B2(net37),
    .ZN(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4495_ (.A1(net83),
    .A2(_0654_),
    .B1(_0655_),
    .B2(net115),
    .ZN(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _4496_ (.A1(_0780_),
    .A2(_0781_),
    .A3(_0782_),
    .A4(_0783_),
    .ZN(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _4497_ (.A1(_0774_),
    .A2(_0779_),
    .A3(_0784_),
    .ZN(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4498_ (.A1(_0720_),
    .A2(_0528_),
    .B1(net1698),
    .B2(_0785_),
    .ZN(_2319_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4499_ (.I(net778),
    .ZN(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4500_ (.I(net504),
    .ZN(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4501_ (.A1(_0787_),
    .A2(_0530_),
    .A3(_0532_),
    .ZN(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4502_ (.A1(net519),
    .A2(_0534_),
    .A3(_0535_),
    .Z(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4503_ (.I(net597),
    .ZN(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4504_ (.A1(_0790_),
    .A2(_0538_),
    .A3(_0725_),
    .ZN(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4505_ (.I(net488),
    .ZN(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4506_ (.A1(_0792_),
    .A2(_0541_),
    .A3(_0542_),
    .ZN(_0793_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _4507_ (.A1(_0788_),
    .A2(_0789_),
    .A3(_0791_),
    .A4(_0793_),
    .ZN(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4508_ (.I(net458),
    .ZN(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4509_ (.I(net441),
    .ZN(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _4510_ (.A1(_0795_),
    .A2(_0548_),
    .A3(_0549_),
    .B1(_0550_),
    .B2(_0796_),
    .ZN(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _4511_ (.A1(net395),
    .A2(_0545_),
    .B1(_0546_),
    .B2(net426),
    .C(_0797_),
    .ZN(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4512_ (.I(net286),
    .ZN(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4513_ (.I(net380),
    .ZN(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _4514_ (.A1(_0799_),
    .A2(_0736_),
    .A3(_0557_),
    .B1(_0558_),
    .B2(_0800_),
    .ZN(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _4515_ (.A1(net208),
    .A2(_0554_),
    .B1(_0555_),
    .B2(net225),
    .C(net1823),
    .ZN(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4516_ (.I(net162),
    .ZN(_0803_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4517_ (.I(net147),
    .ZN(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _4518_ (.A1(_0803_),
    .A2(_0565_),
    .A3(_0566_),
    .B1(_0567_),
    .B2(_0804_),
    .ZN(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _4519_ (.A1(net255),
    .A2(_0562_),
    .B1(_0563_),
    .B2(net240),
    .C(_0805_),
    .ZN(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _4520_ (.A1(_0794_),
    .A2(_0798_),
    .A3(_0802_),
    .A4(_0806_),
    .ZN(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4521_ (.A1(net444),
    .A2(_0572_),
    .B1(_0573_),
    .B2(net99),
    .ZN(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4522_ (.A1(net659),
    .A2(_0575_),
    .B1(_0576_),
    .B2(net131),
    .ZN(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4523_ (.A1(net721),
    .A2(_0578_),
    .B1(_0579_),
    .B2(net706),
    .ZN(_0810_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4524_ (.A1(net675),
    .A2(_0581_),
    .B1(_0582_),
    .B2(net691),
    .ZN(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _4525_ (.A1(net1710),
    .A2(_0809_),
    .A3(_0810_),
    .A4(_0811_),
    .ZN(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4526_ (.A1(net349),
    .A2(_0585_),
    .B1(_0586_),
    .B2(net737),
    .ZN(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4527_ (.A1(net7),
    .A2(_0588_),
    .B1(_0589_),
    .B2(net289),
    .ZN(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4528_ (.A1(net364),
    .A2(_0591_),
    .B1(_0592_),
    .B2(net271),
    .ZN(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4529_ (.A1(net332),
    .A2(_0594_),
    .B(_0753_),
    .ZN(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _4530_ (.A1(_0813_),
    .A2(_0814_),
    .A3(_0815_),
    .A4(_0816_),
    .ZN(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4531_ (.A1(_0807_),
    .A2(_0812_),
    .A3(_0817_),
    .ZN(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4532_ (.I(net846),
    .ZN(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4533_ (.A1(net876),
    .A2(_0602_),
    .A3(_0603_),
    .ZN(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4534_ (.A1(_0819_),
    .A2(_0601_),
    .B(_0820_),
    .ZN(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _4535_ (.A1(net861),
    .A2(_0598_),
    .B1(_0599_),
    .B2(net784),
    .C(_0821_),
    .ZN(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__inv_4 _4536_ (.I(net473),
    .ZN(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4537_ (.I(net830),
    .ZN(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _4538_ (.A1(_0823_),
    .A2(_0610_),
    .A3(_0762_),
    .B1(_0611_),
    .B2(_0824_),
    .ZN(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _4539_ (.A1(net799),
    .A2(_0607_),
    .B1(_0608_),
    .B2(net815),
    .C(_0825_),
    .ZN(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4540_ (.I(net193),
    .ZN(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_8 _4541_ (.I(net768),
    .ZN(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _4542_ (.A1(_0827_),
    .A2(_0618_),
    .B1(_0619_),
    .B2(_0828_),
    .ZN(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _4543_ (.A1(net177),
    .A2(_0615_),
    .B1(_0616_),
    .B2(net887),
    .C(_0829_),
    .ZN(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4544_ (.I(net134),
    .ZN(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4545_ (.I(net600),
    .ZN(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _4546_ (.A1(_0831_),
    .A2(_0626_),
    .B1(_0627_),
    .B2(_0832_),
    .ZN(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _4547_ (.A1(net755),
    .A2(_0623_),
    .B1(_0624_),
    .B2(net752),
    .C(_0833_),
    .ZN(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _4548_ (.A1(net1708),
    .A2(net1706),
    .A3(_0830_),
    .A4(net1705),
    .ZN(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4549_ (.A1(net613),
    .A2(_0632_),
    .B1(_0633_),
    .B2(net628),
    .ZN(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4550_ (.A1(net643),
    .A2(_0635_),
    .B1(_0636_),
    .B2(net535),
    .ZN(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4551_ (.A1(net550),
    .A2(_0638_),
    .B1(_0639_),
    .B2(net566),
    .ZN(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4552_ (.A1(net410),
    .A2(_0641_),
    .B1(_0642_),
    .B2(net582),
    .ZN(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _4553_ (.A1(_0836_),
    .A2(_0837_),
    .A3(_0838_),
    .A4(_0839_),
    .ZN(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4554_ (.A1(net302),
    .A2(_0645_),
    .B1(_0646_),
    .B2(net53),
    .ZN(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4555_ (.A1(net317),
    .A2(_0648_),
    .B1(_0649_),
    .B2(net69),
    .ZN(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4556_ (.A1(net22),
    .A2(_0651_),
    .B1(_0652_),
    .B2(net38),
    .ZN(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4557_ (.A1(net84),
    .A2(_0654_),
    .B1(_0655_),
    .B2(net116),
    .ZN(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _4558_ (.A1(_0841_),
    .A2(_0842_),
    .A3(_0843_),
    .A4(_0844_),
    .ZN(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _4559_ (.A1(_0835_),
    .A2(_0840_),
    .A3(_0845_),
    .ZN(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4560_ (.A1(_0786_),
    .A2(_0528_),
    .B1(net1697),
    .B2(_0846_),
    .ZN(_2320_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _4561_ (.I(net885),
    .ZN(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4562_ (.I(_0013_),
    .Z(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4563_ (.I(_0848_),
    .Z(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4564_ (.I(net505),
    .ZN(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4565_ (.I(_0022_),
    .Z(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4566_ (.I(_0851_),
    .Z(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4567_ (.I(_0531_),
    .Z(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4568_ (.A1(_0850_),
    .A2(_0852_),
    .A3(_0853_),
    .ZN(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4569_ (.I(_0032_),
    .Z(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4570_ (.I(_0855_),
    .Z(_0856_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4571_ (.I(_0039_),
    .Z(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4572_ (.I(_0857_),
    .Z(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4573_ (.A1(net520),
    .A2(_0856_),
    .A3(_0858_),
    .Z(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4574_ (.I(net598),
    .ZN(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4575_ (.I(_0050_),
    .Z(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4576_ (.I(_0861_),
    .Z(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _4577_ (.A1(_0860_),
    .A2(_0862_),
    .A3(_0725_),
    .ZN(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4578_ (.I(net490),
    .ZN(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4579_ (.I(_0119_),
    .Z(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4580_ (.I(_0865_),
    .Z(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4581_ (.I(_0293_),
    .Z(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4582_ (.I(_0867_),
    .Z(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _4583_ (.A1(_0864_),
    .A2(_0866_),
    .A3(_0868_),
    .ZN(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _4584_ (.A1(_0854_),
    .A2(_0859_),
    .A3(_0863_),
    .A4(_0869_),
    .ZN(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4585_ (.I(_0067_),
    .Z(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4586_ (.I(_0871_),
    .Z(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4587_ (.I(_0072_),
    .Z(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4588_ (.I(_0873_),
    .Z(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4589_ (.I(net459),
    .ZN(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4590_ (.I(_0076_),
    .Z(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4591_ (.I(_0876_),
    .Z(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4592_ (.I(_0079_),
    .Z(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4593_ (.I(_0083_),
    .Z(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4594_ (.I(_0879_),
    .Z(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4595_ (.I(net442),
    .ZN(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _4596_ (.A1(_0875_),
    .A2(_0877_),
    .A3(_0878_),
    .B1(_0880_),
    .B2(_0881_),
    .ZN(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _4597_ (.A1(net396),
    .A2(_0872_),
    .B1(_0874_),
    .B2(net427),
    .C(_0882_),
    .ZN(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4598_ (.I(_0091_),
    .Z(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4599_ (.I(_0884_),
    .Z(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4600_ (.I(_0098_),
    .Z(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4601_ (.I(_0886_),
    .Z(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _4602_ (.I(net287),
    .ZN(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4603_ (.I(_0211_),
    .Z(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4604_ (.I(_0889_),
    .Z(_0890_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4605_ (.I(_0110_),
    .Z(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4606_ (.I(_0891_),
    .Z(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4607_ (.I(net381),
    .ZN(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _4608_ (.A1(_0888_),
    .A2(_0736_),
    .A3(_0890_),
    .B1(_0892_),
    .B2(_0893_),
    .ZN(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _4609_ (.A1(net209),
    .A2(_0885_),
    .B1(_0887_),
    .B2(net226),
    .C(_0894_),
    .ZN(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4610_ (.I(_0116_),
    .Z(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4611_ (.I(_0896_),
    .Z(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4612_ (.I(_0120_),
    .Z(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4613_ (.I(_0898_),
    .Z(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4614_ (.I(net163),
    .ZN(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4615_ (.I(_0124_),
    .Z(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4616_ (.I(_0901_),
    .Z(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4617_ (.I(_0127_),
    .Z(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4618_ (.I(_0129_),
    .Z(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4619_ (.I(_0904_),
    .Z(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4620_ (.I(net148),
    .ZN(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _4621_ (.A1(_0900_),
    .A2(_0902_),
    .A3(_0903_),
    .B1(_0905_),
    .B2(_0906_),
    .ZN(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _4622_ (.A1(net257),
    .A2(_0897_),
    .B1(_0899_),
    .B2(net241),
    .C(_0907_),
    .ZN(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _4623_ (.A1(_0870_),
    .A2(_0883_),
    .A3(_0895_),
    .A4(_0908_),
    .ZN(_0909_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4624_ (.I(_0137_),
    .Z(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4625_ (.I(_0910_),
    .Z(_0911_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4626_ (.I(_0141_),
    .Z(_0912_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4627_ (.I(_0912_),
    .Z(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4628_ (.A1(net456),
    .A2(_0911_),
    .B1(_0913_),
    .B2(net101),
    .ZN(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4629_ (.I(_0147_),
    .Z(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4630_ (.I(_0915_),
    .Z(_0916_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4631_ (.I(_0152_),
    .Z(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4632_ (.I(_0917_),
    .Z(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4633_ (.A1(net660),
    .A2(_0916_),
    .B1(_0918_),
    .B2(net132),
    .ZN(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4634_ (.I(_0156_),
    .Z(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4635_ (.I(_0920_),
    .Z(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4636_ (.I(_0161_),
    .Z(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4637_ (.I(_0922_),
    .Z(_0923_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4638_ (.A1(net723),
    .A2(_0921_),
    .B1(_0923_),
    .B2(net707),
    .ZN(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4639_ (.I(_0165_),
    .Z(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4640_ (.I(_0925_),
    .Z(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4641_ (.I(_0168_),
    .Z(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4642_ (.I(_0927_),
    .Z(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4643_ (.A1(net676),
    .A2(_0926_),
    .B1(_0928_),
    .B2(net692),
    .ZN(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _4644_ (.A1(_0914_),
    .A2(_0919_),
    .A3(_0924_),
    .A4(_0929_),
    .ZN(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4645_ (.I(_0174_),
    .Z(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _4646_ (.I(_0931_),
    .Z(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4647_ (.I(_0177_),
    .Z(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4648_ (.I(_0933_),
    .Z(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4649_ (.A1(net350),
    .A2(_0932_),
    .B1(_0934_),
    .B2(net738),
    .ZN(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4650_ (.I(_0181_),
    .Z(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4651_ (.I(_0936_),
    .Z(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4652_ (.I(_0184_),
    .Z(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4653_ (.I(_0938_),
    .Z(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4654_ (.A1(net8),
    .A2(_0937_),
    .B1(_0939_),
    .B2(net300),
    .ZN(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4655_ (.I(_0189_),
    .Z(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4656_ (.I(_0941_),
    .Z(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4657_ (.I(_0195_),
    .Z(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4658_ (.I(_0943_),
    .Z(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4659_ (.A1(net365),
    .A2(_0942_),
    .B1(_0944_),
    .B2(net272),
    .ZN(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4660_ (.I(_0200_),
    .Z(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4661_ (.I(_0946_),
    .Z(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4662_ (.A1(net335),
    .A2(_0947_),
    .B(_0753_),
    .ZN(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _4663_ (.A1(_0935_),
    .A2(_0940_),
    .A3(_0945_),
    .A4(_0948_),
    .ZN(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _4664_ (.A1(_0909_),
    .A2(_0930_),
    .A3(_0949_),
    .ZN(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4665_ (.I(_0208_),
    .Z(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4666_ (.I(_0951_),
    .Z(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4667_ (.I(_0212_),
    .Z(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4668_ (.I(_0953_),
    .Z(_0954_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4669_ (.I(net847),
    .ZN(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _4670_ (.D(_2323_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net1685));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _4671_ (.D(_2326_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net1688));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _4672_ (.D(_2327_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net1689));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _4673_ (.D(_2328_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net1690));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _4674_ (.D(_2329_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net1691));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _4675_ (.D(_2330_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net1692));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _4676_ (.D(_2331_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net1693));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _4677_ (.D(_2332_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net1694));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _4678_ (.D(_2333_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net1695));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _4679_ (.D(_2334_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net1696));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _4680_ (.D(_2324_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net1686));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _4681_ (.D(_2325_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net1687));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4682_ (.D(_2309_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net1671));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4683_ (.D(_2314_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net1676));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4684_ (.D(_2315_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net1677));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4685_ (.D(_2316_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net1678));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4686_ (.D(_2317_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net1679));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4687_ (.D(_2318_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net1680));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4688_ (.D(_2319_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net1681));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4689_ (.D(_2320_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net1682));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4690_ (.D(_2321_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net1683));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4691_ (.D(_2322_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net1684));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4692_ (.D(_2310_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net1672));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _4693_ (.D(_2311_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net1673));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4694_ (.D(_2312_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net1674));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4695_ (.D(_2313_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net1675));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_clk (.I(clk),
    .Z(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_1_0__f_clk (.I(clknet_0_clk),
    .Z(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_1_1__f_clk (.I(clknet_0_clk),
    .Z(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1 (.I(itasegm[0]),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input10 (.I(itasegm[108]),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input100 (.I(itasegm[18]),
    .Z(net100));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1000 (.I(itasel[193]),
    .Z(net1000));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1001 (.I(itasel[194]),
    .Z(net1001));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1002 (.I(itasel[195]),
    .Z(net1002));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1003 (.I(itasel[196]),
    .Z(net1003));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1004 (.I(itasel[197]),
    .Z(net1004));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1005 (.I(itasel[198]),
    .Z(net1005));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1006 (.I(itasel[199]),
    .Z(net1006));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1007 (.I(itasel[19]),
    .Z(net1007));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1008 (.I(itasel[1]),
    .Z(net1008));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1009 (.I(itasel[200]),
    .Z(net1009));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input101 (.I(itasegm[190]),
    .Z(net101));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1010 (.I(itasel[201]),
    .Z(net1010));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1011 (.I(itasel[202]),
    .Z(net1011));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1012 (.I(itasel[203]),
    .Z(net1012));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1013 (.I(itasel[204]),
    .Z(net1013));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1014 (.I(itasel[205]),
    .Z(net1014));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1015 (.I(itasel[206]),
    .Z(net1015));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1016 (.I(itasel[207]),
    .Z(net1016));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1017 (.I(itasel[208]),
    .Z(net1017));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1018 (.I(itasel[209]),
    .Z(net1018));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1019 (.I(itasel[20]),
    .Z(net1019));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input102 (.I(itasegm[191]),
    .Z(net102));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1020 (.I(itasel[210]),
    .Z(net1020));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1021 (.I(itasel[211]),
    .Z(net1021));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1022 (.I(itasel[212]),
    .Z(net1022));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1023 (.I(itasel[213]),
    .Z(net1023));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1024 (.I(itasel[214]),
    .Z(net1024));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1025 (.I(itasel[215]),
    .Z(net1025));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input1026 (.I(itasel[216]),
    .Z(net1026));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input1027 (.I(itasel[217]),
    .Z(net1027));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1028 (.I(itasel[218]),
    .Z(net1028));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1029 (.I(itasel[219]),
    .Z(net1029));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input103 (.I(itasegm[192]),
    .Z(net103));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1030 (.I(itasel[21]),
    .Z(net1030));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1031 (.I(itasel[220]),
    .Z(net1031));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1032 (.I(itasel[221]),
    .Z(net1032));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1033 (.I(itasel[222]),
    .Z(net1033));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1034 (.I(itasel[223]),
    .Z(net1034));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1035 (.I(itasel[224]),
    .Z(net1035));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1036 (.I(itasel[225]),
    .Z(net1036));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1037 (.I(itasel[226]),
    .Z(net1037));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1038 (.I(itasel[227]),
    .Z(net1038));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1039 (.I(itasel[228]),
    .Z(net1039));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input104 (.I(itasegm[193]),
    .Z(net104));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1040 (.I(itasel[229]),
    .Z(net1040));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1041 (.I(itasel[22]),
    .Z(net1041));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1042 (.I(itasel[230]),
    .Z(net1042));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1043 (.I(itasel[231]),
    .Z(net1043));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1044 (.I(itasel[232]),
    .Z(net1044));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1045 (.I(itasel[233]),
    .Z(net1045));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1046 (.I(itasel[234]),
    .Z(net1046));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1047 (.I(itasel[235]),
    .Z(net1047));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1048 (.I(itasel[236]),
    .Z(net1048));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1049 (.I(itasel[237]),
    .Z(net1049));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input105 (.I(itasegm[194]),
    .Z(net105));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1050 (.I(itasel[238]),
    .Z(net1050));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1051 (.I(itasel[239]),
    .Z(net1051));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1052 (.I(itasel[23]),
    .Z(net1052));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1053 (.I(itasel[240]),
    .Z(net1053));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1054 (.I(itasel[241]),
    .Z(net1054));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1055 (.I(itasel[242]),
    .Z(net1055));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1056 (.I(itasel[243]),
    .Z(net1056));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1057 (.I(itasel[244]),
    .Z(net1057));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1058 (.I(itasel[245]),
    .Z(net1058));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1059 (.I(itasel[246]),
    .Z(net1059));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input106 (.I(itasegm[195]),
    .Z(net106));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1060 (.I(itasel[247]),
    .Z(net1060));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1061 (.I(itasel[248]),
    .Z(net1061));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1062 (.I(itasel[249]),
    .Z(net1062));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1063 (.I(itasel[24]),
    .Z(net1063));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1064 (.I(itasel[250]),
    .Z(net1064));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1065 (.I(itasel[251]),
    .Z(net1065));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1066 (.I(itasel[252]),
    .Z(net1066));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1067 (.I(itasel[253]),
    .Z(net1067));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1068 (.I(itasel[254]),
    .Z(net1068));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1069 (.I(itasel[255]),
    .Z(net1069));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input107 (.I(itasegm[196]),
    .Z(net107));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1070 (.I(itasel[256]),
    .Z(net1070));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1071 (.I(itasel[257]),
    .Z(net1071));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1072 (.I(itasel[258]),
    .Z(net1072));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1073 (.I(itasel[259]),
    .Z(net1073));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1074 (.I(itasel[25]),
    .Z(net1074));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1075 (.I(itasel[260]),
    .Z(net1075));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1076 (.I(itasel[261]),
    .Z(net1076));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1077 (.I(itasel[262]),
    .Z(net1077));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1078 (.I(itasel[263]),
    .Z(net1078));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1079 (.I(itasel[264]),
    .Z(net1079));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input108 (.I(itasegm[197]),
    .Z(net108));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1080 (.I(itasel[265]),
    .Z(net1080));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1081 (.I(itasel[266]),
    .Z(net1081));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1082 (.I(itasel[267]),
    .Z(net1082));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1083 (.I(itasel[268]),
    .Z(net1083));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1084 (.I(itasel[269]),
    .Z(net1084));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1085 (.I(itasel[26]),
    .Z(net1085));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1086 (.I(itasel[270]),
    .Z(net1086));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1087 (.I(itasel[271]),
    .Z(net1087));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1088 (.I(itasel[272]),
    .Z(net1088));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1089 (.I(itasel[273]),
    .Z(net1089));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input109 (.I(itasegm[198]),
    .Z(net109));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1090 (.I(itasel[274]),
    .Z(net1090));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1091 (.I(itasel[275]),
    .Z(net1091));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1092 (.I(itasel[276]),
    .Z(net1092));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1093 (.I(itasel[277]),
    .Z(net1093));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1094 (.I(itasel[278]),
    .Z(net1094));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1095 (.I(itasel[279]),
    .Z(net1095));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1096 (.I(itasel[27]),
    .Z(net1096));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1097 (.I(itasel[280]),
    .Z(net1097));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1098 (.I(itasel[281]),
    .Z(net1098));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1099 (.I(itasel[282]),
    .Z(net1099));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input11 (.I(itasegm[109]),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input110 (.I(itasegm[199]),
    .Z(net110));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1100 (.I(itasel[283]),
    .Z(net1100));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1101 (.I(itasel[284]),
    .Z(net1101));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1102 (.I(itasel[285]),
    .Z(net1102));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1103 (.I(itasel[286]),
    .Z(net1103));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1104 (.I(itasel[287]),
    .Z(net1104));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1105 (.I(itasel[288]),
    .Z(net1105));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1106 (.I(itasel[289]),
    .Z(net1106));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1107 (.I(itasel[28]),
    .Z(net1107));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1108 (.I(itasel[290]),
    .Z(net1108));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1109 (.I(itasel[291]),
    .Z(net1109));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input111 (.I(itasegm[19]),
    .Z(net111));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1110 (.I(itasel[292]),
    .Z(net1110));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1111 (.I(itasel[293]),
    .Z(net1111));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1112 (.I(itasel[294]),
    .Z(net1112));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1113 (.I(itasel[295]),
    .Z(net1113));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1114 (.I(itasel[296]),
    .Z(net1114));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1115 (.I(itasel[297]),
    .Z(net1115));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1116 (.I(itasel[298]),
    .Z(net1116));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1117 (.I(itasel[299]),
    .Z(net1117));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1118 (.I(itasel[29]),
    .Z(net1118));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1119 (.I(itasel[2]),
    .Z(net1119));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input112 (.I(itasegm[1]),
    .Z(net112));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1120 (.I(itasel[300]),
    .Z(net1120));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1121 (.I(itasel[301]),
    .Z(net1121));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1122 (.I(itasel[302]),
    .Z(net1122));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1123 (.I(itasel[303]),
    .Z(net1123));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1124 (.I(itasel[304]),
    .Z(net1124));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1125 (.I(itasel[305]),
    .Z(net1125));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1126 (.I(itasel[306]),
    .Z(net1126));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1127 (.I(itasel[307]),
    .Z(net1127));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1128 (.I(itasel[308]),
    .Z(net1128));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1129 (.I(itasel[309]),
    .Z(net1129));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input113 (.I(itasegm[200]),
    .Z(net113));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1130 (.I(itasel[30]),
    .Z(net1130));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1131 (.I(itasel[310]),
    .Z(net1131));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1132 (.I(itasel[311]),
    .Z(net1132));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input1133 (.I(itasel[312]),
    .Z(net1133));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input1134 (.I(itasel[313]),
    .Z(net1134));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input1135 (.I(itasel[314]),
    .Z(net1135));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input1136 (.I(itasel[315]),
    .Z(net1136));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input1137 (.I(itasel[316]),
    .Z(net1137));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input1138 (.I(itasel[317]),
    .Z(net1138));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input1139 (.I(itasel[318]),
    .Z(net1139));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input114 (.I(itasegm[201]),
    .Z(net114));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input1140 (.I(itasel[319]),
    .Z(net1140));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1141 (.I(itasel[31]),
    .Z(net1141));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input1142 (.I(itasel[320]),
    .Z(net1142));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input1143 (.I(itasel[321]),
    .Z(net1143));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input1144 (.I(itasel[322]),
    .Z(net1144));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input1145 (.I(itasel[323]),
    .Z(net1145));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input1146 (.I(itasel[324]),
    .Z(net1146));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input1147 (.I(itasel[325]),
    .Z(net1147));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input1148 (.I(itasel[326]),
    .Z(net1148));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input1149 (.I(itasel[327]),
    .Z(net1149));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input115 (.I(itasegm[202]),
    .Z(net115));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input1150 (.I(itasel[328]),
    .Z(net1150));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input1151 (.I(itasel[329]),
    .Z(net1151));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1152 (.I(itasel[32]),
    .Z(net1152));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input1153 (.I(itasel[330]),
    .Z(net1153));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input1154 (.I(itasel[331]),
    .Z(net1154));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input1155 (.I(itasel[332]),
    .Z(net1155));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input1156 (.I(itasel[333]),
    .Z(net1156));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input1157 (.I(itasel[334]),
    .Z(net1157));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input1158 (.I(itasel[335]),
    .Z(net1158));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1159 (.I(itasel[336]),
    .Z(net1159));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input116 (.I(itasegm[203]),
    .Z(net116));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1160 (.I(itasel[337]),
    .Z(net1160));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1161 (.I(itasel[338]),
    .Z(net1161));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1162 (.I(itasel[339]),
    .Z(net1162));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1163 (.I(itasel[33]),
    .Z(net1163));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1164 (.I(itasel[340]),
    .Z(net1164));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1165 (.I(itasel[341]),
    .Z(net1165));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1166 (.I(itasel[342]),
    .Z(net1166));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1167 (.I(itasel[343]),
    .Z(net1167));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1168 (.I(itasel[344]),
    .Z(net1168));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1169 (.I(itasel[345]),
    .Z(net1169));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input117 (.I(itasegm[204]),
    .Z(net117));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1170 (.I(itasel[346]),
    .Z(net1170));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1171 (.I(itasel[347]),
    .Z(net1171));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1172 (.I(itasel[348]),
    .Z(net1172));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1173 (.I(itasel[349]),
    .Z(net1173));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1174 (.I(itasel[34]),
    .Z(net1174));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1175 (.I(itasel[350]),
    .Z(net1175));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1176 (.I(itasel[351]),
    .Z(net1176));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1177 (.I(itasel[352]),
    .Z(net1177));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1178 (.I(itasel[353]),
    .Z(net1178));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1179 (.I(itasel[354]),
    .Z(net1179));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input118 (.I(itasegm[205]),
    .Z(net118));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1180 (.I(itasel[355]),
    .Z(net1180));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1181 (.I(itasel[356]),
    .Z(net1181));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1182 (.I(itasel[357]),
    .Z(net1182));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1183 (.I(itasel[358]),
    .Z(net1183));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1184 (.I(itasel[359]),
    .Z(net1184));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1185 (.I(itasel[35]),
    .Z(net1185));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1186 (.I(itasel[360]),
    .Z(net1186));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1187 (.I(itasel[361]),
    .Z(net1187));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1188 (.I(itasel[362]),
    .Z(net1188));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1189 (.I(itasel[363]),
    .Z(net1189));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input119 (.I(itasegm[206]),
    .Z(net119));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1190 (.I(itasel[364]),
    .Z(net1190));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1191 (.I(itasel[365]),
    .Z(net1191));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1192 (.I(itasel[366]),
    .Z(net1192));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1193 (.I(itasel[367]),
    .Z(net1193));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1194 (.I(itasel[368]),
    .Z(net1194));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1195 (.I(itasel[369]),
    .Z(net1195));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input1196 (.I(itasel[36]),
    .Z(net1196));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1197 (.I(itasel[370]),
    .Z(net1197));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1198 (.I(itasel[371]),
    .Z(net1198));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1199 (.I(itasel[372]),
    .Z(net1199));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input12 (.I(itasegm[10]),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input120 (.I(itasegm[207]),
    .Z(net120));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1200 (.I(itasel[373]),
    .Z(net1200));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1201 (.I(itasel[374]),
    .Z(net1201));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1202 (.I(itasel[375]),
    .Z(net1202));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1203 (.I(itasel[376]),
    .Z(net1203));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1204 (.I(itasel[377]),
    .Z(net1204));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1205 (.I(itasel[378]),
    .Z(net1205));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1206 (.I(itasel[379]),
    .Z(net1206));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input1207 (.I(itasel[37]),
    .Z(net1207));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1208 (.I(itasel[380]),
    .Z(net1208));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1209 (.I(itasel[381]),
    .Z(net1209));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input121 (.I(itasegm[208]),
    .Z(net121));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1210 (.I(itasel[382]),
    .Z(net1210));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1211 (.I(itasel[383]),
    .Z(net1211));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1212 (.I(itasel[384]),
    .Z(net1212));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1213 (.I(itasel[385]),
    .Z(net1213));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1214 (.I(itasel[386]),
    .Z(net1214));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1215 (.I(itasel[387]),
    .Z(net1215));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1216 (.I(itasel[388]),
    .Z(net1216));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1217 (.I(itasel[389]),
    .Z(net1217));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input1218 (.I(itasel[38]),
    .Z(net1218));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1219 (.I(itasel[390]),
    .Z(net1219));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input122 (.I(itasegm[209]),
    .Z(net122));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1220 (.I(itasel[391]),
    .Z(net1220));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1221 (.I(itasel[392]),
    .Z(net1221));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1222 (.I(itasel[393]),
    .Z(net1222));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1223 (.I(itasel[394]),
    .Z(net1223));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1224 (.I(itasel[395]),
    .Z(net1224));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input1225 (.I(itasel[396]),
    .Z(net1225));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input1226 (.I(itasel[397]),
    .Z(net1226));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1227 (.I(itasel[398]),
    .Z(net1227));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1228 (.I(itasel[399]),
    .Z(net1228));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input1229 (.I(itasel[39]),
    .Z(net1229));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input123 (.I(itasegm[20]),
    .Z(net123));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1230 (.I(itasel[3]),
    .Z(net1230));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1231 (.I(itasel[400]),
    .Z(net1231));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1232 (.I(itasel[401]),
    .Z(net1232));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1233 (.I(itasel[402]),
    .Z(net1233));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1234 (.I(itasel[403]),
    .Z(net1234));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1235 (.I(itasel[404]),
    .Z(net1235));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1236 (.I(itasel[405]),
    .Z(net1236));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1237 (.I(itasel[406]),
    .Z(net1237));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1238 (.I(itasel[407]),
    .Z(net1238));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1239 (.I(itasel[408]),
    .Z(net1239));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 input124 (.I(itasegm[210]),
    .Z(net124));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1240 (.I(itasel[409]),
    .Z(net1240));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input1241 (.I(itasel[40]),
    .Z(net1241));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1242 (.I(itasel[410]),
    .Z(net1242));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1243 (.I(itasel[411]),
    .Z(net1243));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1244 (.I(itasel[412]),
    .Z(net1244));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1245 (.I(itasel[413]),
    .Z(net1245));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1246 (.I(itasel[414]),
    .Z(net1246));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1247 (.I(itasel[415]),
    .Z(net1247));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1248 (.I(itasel[416]),
    .Z(net1248));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1249 (.I(itasel[417]),
    .Z(net1249));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 input125 (.I(itasegm[211]),
    .Z(net125));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1250 (.I(itasel[418]),
    .Z(net1250));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1251 (.I(itasel[419]),
    .Z(net1251));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input1252 (.I(itasel[41]),
    .Z(net1252));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1253 (.I(itasel[420]),
    .Z(net1253));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1254 (.I(itasel[421]),
    .Z(net1254));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1255 (.I(itasel[422]),
    .Z(net1255));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1256 (.I(itasel[423]),
    .Z(net1256));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1257 (.I(itasel[424]),
    .Z(net1257));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1258 (.I(itasel[425]),
    .Z(net1258));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1259 (.I(itasel[426]),
    .Z(net1259));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 input126 (.I(itasegm[212]),
    .Z(net126));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1260 (.I(itasel[427]),
    .Z(net1260));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1261 (.I(itasel[428]),
    .Z(net1261));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1262 (.I(itasel[429]),
    .Z(net1262));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input1263 (.I(itasel[42]),
    .Z(net1263));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1264 (.I(itasel[430]),
    .Z(net1264));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1265 (.I(itasel[431]),
    .Z(net1265));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1266 (.I(itasel[432]),
    .Z(net1266));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1267 (.I(itasel[433]),
    .Z(net1267));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1268 (.I(itasel[434]),
    .Z(net1268));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1269 (.I(itasel[435]),
    .Z(net1269));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 input127 (.I(itasegm[213]),
    .Z(net127));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1270 (.I(itasel[436]),
    .Z(net1270));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1271 (.I(itasel[437]),
    .Z(net1271));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1272 (.I(itasel[438]),
    .Z(net1272));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1273 (.I(itasel[439]),
    .Z(net1273));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input1274 (.I(itasel[43]),
    .Z(net1274));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1275 (.I(itasel[440]),
    .Z(net1275));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1276 (.I(itasel[441]),
    .Z(net1276));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1277 (.I(itasel[442]),
    .Z(net1277));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1278 (.I(itasel[443]),
    .Z(net1278));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1279 (.I(itasel[444]),
    .Z(net1279));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 input128 (.I(itasegm[214]),
    .Z(net128));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1280 (.I(itasel[445]),
    .Z(net1280));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1281 (.I(itasel[446]),
    .Z(net1281));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1282 (.I(itasel[447]),
    .Z(net1282));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1283 (.I(itasel[448]),
    .Z(net1283));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1284 (.I(itasel[449]),
    .Z(net1284));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input1285 (.I(itasel[44]),
    .Z(net1285));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1286 (.I(itasel[450]),
    .Z(net1286));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1287 (.I(itasel[451]),
    .Z(net1287));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1288 (.I(itasel[452]),
    .Z(net1288));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1289 (.I(itasel[453]),
    .Z(net1289));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 input129 (.I(itasegm[215]),
    .Z(net129));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1290 (.I(itasel[454]),
    .Z(net1290));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1291 (.I(itasel[455]),
    .Z(net1291));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1292 (.I(itasel[456]),
    .Z(net1292));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1293 (.I(itasel[457]),
    .Z(net1293));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1294 (.I(itasel[458]),
    .Z(net1294));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1295 (.I(itasel[459]),
    .Z(net1295));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input1296 (.I(itasel[45]),
    .Z(net1296));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1297 (.I(itasel[460]),
    .Z(net1297));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1298 (.I(itasel[461]),
    .Z(net1298));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1299 (.I(itasel[462]),
    .Z(net1299));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input13 (.I(itasegm[110]),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 input130 (.I(itasegm[216]),
    .Z(net130));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1300 (.I(itasel[463]),
    .Z(net1300));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1301 (.I(itasel[464]),
    .Z(net1301));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1302 (.I(itasel[465]),
    .Z(net1302));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1303 (.I(itasel[466]),
    .Z(net1303));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1304 (.I(itasel[467]),
    .Z(net1304));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1305 (.I(itasel[468]),
    .Z(net1305));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1306 (.I(itasel[469]),
    .Z(net1306));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input1307 (.I(itasel[46]),
    .Z(net1307));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1308 (.I(itasel[470]),
    .Z(net1308));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1309 (.I(itasel[471]),
    .Z(net1309));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 input131 (.I(itasegm[217]),
    .Z(net131));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1310 (.I(itasel[472]),
    .Z(net1310));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1311 (.I(itasel[473]),
    .Z(net1311));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1312 (.I(itasel[474]),
    .Z(net1312));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1313 (.I(itasel[475]),
    .Z(net1313));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1314 (.I(itasel[476]),
    .Z(net1314));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1315 (.I(itasel[477]),
    .Z(net1315));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1316 (.I(itasel[478]),
    .Z(net1316));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1317 (.I(itasel[479]),
    .Z(net1317));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input1318 (.I(itasel[47]),
    .Z(net1318));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1319 (.I(itasel[480]),
    .Z(net1319));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input132 (.I(itasegm[218]),
    .Z(net132));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1320 (.I(itasel[481]),
    .Z(net1320));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1321 (.I(itasel[482]),
    .Z(net1321));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1322 (.I(itasel[483]),
    .Z(net1322));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1323 (.I(itasel[484]),
    .Z(net1323));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1324 (.I(itasel[485]),
    .Z(net1324));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1325 (.I(itasel[486]),
    .Z(net1325));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1326 (.I(itasel[487]),
    .Z(net1326));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1327 (.I(itasel[488]),
    .Z(net1327));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1328 (.I(itasel[489]),
    .Z(net1328));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1329 (.I(itasel[48]),
    .Z(net1329));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input133 (.I(itasegm[219]),
    .Z(net133));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1330 (.I(itasel[490]),
    .Z(net1330));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1331 (.I(itasel[491]),
    .Z(net1331));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1332 (.I(itasel[492]),
    .Z(net1332));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1333 (.I(itasel[493]),
    .Z(net1333));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1334 (.I(itasel[494]),
    .Z(net1334));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1335 (.I(itasel[495]),
    .Z(net1335));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1336 (.I(itasel[496]),
    .Z(net1336));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1337 (.I(itasel[497]),
    .Z(net1337));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1338 (.I(itasel[498]),
    .Z(net1338));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1339 (.I(itasel[499]),
    .Z(net1339));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input134 (.I(itasegm[21]),
    .Z(net134));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1340 (.I(itasel[49]),
    .Z(net1340));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input1341 (.I(itasel[4]),
    .Z(net1341));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1342 (.I(itasel[500]),
    .Z(net1342));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1343 (.I(itasel[501]),
    .Z(net1343));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1344 (.I(itasel[502]),
    .Z(net1344));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1345 (.I(itasel[503]),
    .Z(net1345));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1346 (.I(itasel[504]),
    .Z(net1346));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1347 (.I(itasel[505]),
    .Z(net1347));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1348 (.I(itasel[506]),
    .Z(net1348));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1349 (.I(itasel[507]),
    .Z(net1349));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input135 (.I(itasegm[220]),
    .Z(net135));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1350 (.I(itasel[508]),
    .Z(net1350));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1351 (.I(itasel[509]),
    .Z(net1351));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1352 (.I(itasel[50]),
    .Z(net1352));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1353 (.I(itasel[510]),
    .Z(net1353));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1354 (.I(itasel[511]),
    .Z(net1354));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1355 (.I(itasel[512]),
    .Z(net1355));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1356 (.I(itasel[513]),
    .Z(net1356));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1357 (.I(itasel[514]),
    .Z(net1357));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1358 (.I(itasel[515]),
    .Z(net1358));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1359 (.I(itasel[516]),
    .Z(net1359));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input136 (.I(itasegm[221]),
    .Z(net136));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1360 (.I(itasel[517]),
    .Z(net1360));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1361 (.I(itasel[518]),
    .Z(net1361));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1362 (.I(itasel[519]),
    .Z(net1362));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1363 (.I(itasel[51]),
    .Z(net1363));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1364 (.I(itasel[520]),
    .Z(net1364));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1365 (.I(itasel[521]),
    .Z(net1365));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1366 (.I(itasel[522]),
    .Z(net1366));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1367 (.I(itasel[523]),
    .Z(net1367));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1368 (.I(itasel[524]),
    .Z(net1368));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1369 (.I(itasel[525]),
    .Z(net1369));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input137 (.I(itasegm[222]),
    .Z(net137));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1370 (.I(itasel[526]),
    .Z(net1370));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1371 (.I(itasel[527]),
    .Z(net1371));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1372 (.I(itasel[528]),
    .Z(net1372));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1373 (.I(itasel[529]),
    .Z(net1373));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1374 (.I(itasel[52]),
    .Z(net1374));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1375 (.I(itasel[530]),
    .Z(net1375));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1376 (.I(itasel[531]),
    .Z(net1376));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1377 (.I(itasel[532]),
    .Z(net1377));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1378 (.I(itasel[533]),
    .Z(net1378));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1379 (.I(itasel[534]),
    .Z(net1379));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input138 (.I(itasegm[223]),
    .Z(net138));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1380 (.I(itasel[535]),
    .Z(net1380));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1381 (.I(itasel[536]),
    .Z(net1381));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1382 (.I(itasel[537]),
    .Z(net1382));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1383 (.I(itasel[538]),
    .Z(net1383));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1384 (.I(itasel[539]),
    .Z(net1384));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1385 (.I(itasel[53]),
    .Z(net1385));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1386 (.I(itasel[540]),
    .Z(net1386));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1387 (.I(itasel[541]),
    .Z(net1387));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1388 (.I(itasel[542]),
    .Z(net1388));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1389 (.I(itasel[543]),
    .Z(net1389));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input139 (.I(itasegm[224]),
    .Z(net139));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1390 (.I(itasel[544]),
    .Z(net1390));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1391 (.I(itasel[545]),
    .Z(net1391));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1392 (.I(itasel[546]),
    .Z(net1392));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1393 (.I(itasel[547]),
    .Z(net1393));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1394 (.I(itasel[548]),
    .Z(net1394));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1395 (.I(itasel[549]),
    .Z(net1395));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1396 (.I(itasel[54]),
    .Z(net1396));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1397 (.I(itasel[550]),
    .Z(net1397));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1398 (.I(itasel[551]),
    .Z(net1398));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1399 (.I(itasel[552]),
    .Z(net1399));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input14 (.I(itasegm[111]),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input140 (.I(itasegm[225]),
    .Z(net140));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1400 (.I(itasel[553]),
    .Z(net1400));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1401 (.I(itasel[554]),
    .Z(net1401));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1402 (.I(itasel[555]),
    .Z(net1402));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1403 (.I(itasel[556]),
    .Z(net1403));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1404 (.I(itasel[557]),
    .Z(net1404));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1405 (.I(itasel[558]),
    .Z(net1405));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1406 (.I(itasel[559]),
    .Z(net1406));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1407 (.I(itasel[55]),
    .Z(net1407));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1408 (.I(itasel[560]),
    .Z(net1408));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1409 (.I(itasel[561]),
    .Z(net1409));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input141 (.I(itasegm[226]),
    .Z(net141));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1410 (.I(itasel[562]),
    .Z(net1410));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1411 (.I(itasel[563]),
    .Z(net1411));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1412 (.I(itasel[564]),
    .Z(net1412));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1413 (.I(itasel[565]),
    .Z(net1413));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1414 (.I(itasel[566]),
    .Z(net1414));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1415 (.I(itasel[567]),
    .Z(net1415));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1416 (.I(itasel[568]),
    .Z(net1416));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1417 (.I(itasel[569]),
    .Z(net1417));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1418 (.I(itasel[56]),
    .Z(net1418));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1419 (.I(itasel[570]),
    .Z(net1419));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input142 (.I(itasegm[227]),
    .Z(net142));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1420 (.I(itasel[571]),
    .Z(net1420));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1421 (.I(itasel[572]),
    .Z(net1421));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1422 (.I(itasel[573]),
    .Z(net1422));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1423 (.I(itasel[574]),
    .Z(net1423));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1424 (.I(itasel[575]),
    .Z(net1424));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1425 (.I(itasel[576]),
    .Z(net1425));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1426 (.I(itasel[577]),
    .Z(net1426));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1427 (.I(itasel[578]),
    .Z(net1427));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1428 (.I(itasel[579]),
    .Z(net1428));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1429 (.I(itasel[57]),
    .Z(net1429));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input143 (.I(itasegm[228]),
    .Z(net143));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1430 (.I(itasel[580]),
    .Z(net1430));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1431 (.I(itasel[581]),
    .Z(net1431));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1432 (.I(itasel[582]),
    .Z(net1432));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1433 (.I(itasel[583]),
    .Z(net1433));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1434 (.I(itasel[584]),
    .Z(net1434));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1435 (.I(itasel[585]),
    .Z(net1435));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1436 (.I(itasel[586]),
    .Z(net1436));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1437 (.I(itasel[587]),
    .Z(net1437));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input1438 (.I(itasel[588]),
    .Z(net1438));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input1439 (.I(itasel[589]),
    .Z(net1439));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input144 (.I(itasegm[229]),
    .Z(net144));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1440 (.I(itasel[58]),
    .Z(net1440));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input1441 (.I(itasel[590]),
    .Z(net1441));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input1442 (.I(itasel[591]),
    .Z(net1442));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input1443 (.I(itasel[592]),
    .Z(net1443));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input1444 (.I(itasel[593]),
    .Z(net1444));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input1445 (.I(itasel[594]),
    .Z(net1445));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 input1446 (.I(itasel[595]),
    .Z(net1446));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input1447 (.I(itasel[596]),
    .Z(net1447));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input1448 (.I(itasel[597]),
    .Z(net1448));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1449 (.I(itasel[598]),
    .Z(net1449));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input145 (.I(itasegm[22]),
    .Z(net145));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1450 (.I(itasel[599]),
    .Z(net1450));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1451 (.I(itasel[59]),
    .Z(net1451));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input1452 (.I(itasel[5]),
    .Z(net1452));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1453 (.I(itasel[600]),
    .Z(net1453));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1454 (.I(itasel[601]),
    .Z(net1454));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1455 (.I(itasel[602]),
    .Z(net1455));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1456 (.I(itasel[603]),
    .Z(net1456));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1457 (.I(itasel[604]),
    .Z(net1457));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1458 (.I(itasel[605]),
    .Z(net1458));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1459 (.I(itasel[606]),
    .Z(net1459));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input146 (.I(itasegm[230]),
    .Z(net146));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1460 (.I(itasel[607]),
    .Z(net1460));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1461 (.I(itasel[608]),
    .Z(net1461));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1462 (.I(itasel[609]),
    .Z(net1462));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1463 (.I(itasel[60]),
    .Z(net1463));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1464 (.I(itasel[610]),
    .Z(net1464));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1465 (.I(itasel[611]),
    .Z(net1465));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1466 (.I(itasel[612]),
    .Z(net1466));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1467 (.I(itasel[613]),
    .Z(net1467));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1468 (.I(itasel[614]),
    .Z(net1468));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1469 (.I(itasel[615]),
    .Z(net1469));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input147 (.I(itasegm[231]),
    .Z(net147));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1470 (.I(itasel[616]),
    .Z(net1470));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1471 (.I(itasel[617]),
    .Z(net1471));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1472 (.I(itasel[618]),
    .Z(net1472));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1473 (.I(itasel[619]),
    .Z(net1473));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1474 (.I(itasel[61]),
    .Z(net1474));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1475 (.I(itasel[620]),
    .Z(net1475));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1476 (.I(itasel[621]),
    .Z(net1476));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1477 (.I(itasel[622]),
    .Z(net1477));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1478 (.I(itasel[623]),
    .Z(net1478));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1479 (.I(itasel[624]),
    .Z(net1479));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input148 (.I(itasegm[232]),
    .Z(net148));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1480 (.I(itasel[625]),
    .Z(net1480));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1481 (.I(itasel[626]),
    .Z(net1481));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1482 (.I(itasel[627]),
    .Z(net1482));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1483 (.I(itasel[628]),
    .Z(net1483));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1484 (.I(itasel[629]),
    .Z(net1484));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1485 (.I(itasel[62]),
    .Z(net1485));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1486 (.I(itasel[630]),
    .Z(net1486));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1487 (.I(itasel[631]),
    .Z(net1487));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1488 (.I(itasel[632]),
    .Z(net1488));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1489 (.I(itasel[633]),
    .Z(net1489));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input149 (.I(itasegm[233]),
    .Z(net149));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1490 (.I(itasel[634]),
    .Z(net1490));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1491 (.I(itasel[635]),
    .Z(net1491));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1492 (.I(itasel[636]),
    .Z(net1492));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1493 (.I(itasel[637]),
    .Z(net1493));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1494 (.I(itasel[638]),
    .Z(net1494));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1495 (.I(itasel[639]),
    .Z(net1495));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1496 (.I(itasel[63]),
    .Z(net1496));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1497 (.I(itasel[640]),
    .Z(net1497));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1498 (.I(itasel[641]),
    .Z(net1498));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1499 (.I(itasel[642]),
    .Z(net1499));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input15 (.I(itasegm[112]),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input150 (.I(itasegm[234]),
    .Z(net150));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1500 (.I(itasel[643]),
    .Z(net1500));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1501 (.I(itasel[644]),
    .Z(net1501));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1502 (.I(itasel[645]),
    .Z(net1502));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1503 (.I(itasel[646]),
    .Z(net1503));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1504 (.I(itasel[647]),
    .Z(net1504));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 input1505 (.I(itasel[648]),
    .Z(net1505));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 input1506 (.I(itasel[649]),
    .Z(net1506));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1507 (.I(itasel[64]),
    .Z(net1507));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 input1508 (.I(itasel[650]),
    .Z(net1508));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 input1509 (.I(itasel[651]),
    .Z(net1509));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input151 (.I(itasegm[235]),
    .Z(net151));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 input1510 (.I(itasel[652]),
    .Z(net1510));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 input1511 (.I(itasel[653]),
    .Z(net1511));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 input1512 (.I(itasel[654]),
    .Z(net1512));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 input1513 (.I(itasel[655]),
    .Z(net1513));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input1514 (.I(itasel[656]),
    .Z(net1514));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 input1515 (.I(itasel[657]),
    .Z(net1515));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input1516 (.I(itasel[658]),
    .Z(net1516));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input1517 (.I(itasel[659]),
    .Z(net1517));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1518 (.I(itasel[65]),
    .Z(net1518));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 input1519 (.I(itasel[660]),
    .Z(net1519));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input152 (.I(itasegm[236]),
    .Z(net152));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 input1520 (.I(itasel[661]),
    .Z(net1520));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 input1521 (.I(itasel[662]),
    .Z(net1521));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 input1522 (.I(itasel[663]),
    .Z(net1522));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 input1523 (.I(itasel[664]),
    .Z(net1523));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 input1524 (.I(itasel[665]),
    .Z(net1524));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 input1525 (.I(itasel[666]),
    .Z(net1525));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 input1526 (.I(itasel[667]),
    .Z(net1526));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 input1527 (.I(itasel[668]),
    .Z(net1527));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 input1528 (.I(itasel[669]),
    .Z(net1528));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1529 (.I(itasel[66]),
    .Z(net1529));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input153 (.I(itasegm[237]),
    .Z(net153));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 input1530 (.I(itasel[670]),
    .Z(net1530));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 input1531 (.I(itasel[671]),
    .Z(net1531));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1532 (.I(itasel[672]),
    .Z(net1532));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1533 (.I(itasel[673]),
    .Z(net1533));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1534 (.I(itasel[674]),
    .Z(net1534));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1535 (.I(itasel[675]),
    .Z(net1535));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1536 (.I(itasel[676]),
    .Z(net1536));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1537 (.I(itasel[677]),
    .Z(net1537));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1538 (.I(itasel[678]),
    .Z(net1538));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1539 (.I(itasel[679]),
    .Z(net1539));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input154 (.I(itasegm[238]),
    .Z(net154));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1540 (.I(itasel[67]),
    .Z(net1540));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1541 (.I(itasel[680]),
    .Z(net1541));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1542 (.I(itasel[681]),
    .Z(net1542));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1543 (.I(itasel[682]),
    .Z(net1543));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1544 (.I(itasel[683]),
    .Z(net1544));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1545 (.I(itasel[684]),
    .Z(net1545));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1546 (.I(itasel[685]),
    .Z(net1546));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1547 (.I(itasel[686]),
    .Z(net1547));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1548 (.I(itasel[687]),
    .Z(net1548));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1549 (.I(itasel[688]),
    .Z(net1549));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input155 (.I(itasegm[239]),
    .Z(net155));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1550 (.I(itasel[689]),
    .Z(net1550));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1551 (.I(itasel[68]),
    .Z(net1551));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1552 (.I(itasel[690]),
    .Z(net1552));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1553 (.I(itasel[691]),
    .Z(net1553));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1554 (.I(itasel[692]),
    .Z(net1554));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1555 (.I(itasel[693]),
    .Z(net1555));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1556 (.I(itasel[694]),
    .Z(net1556));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1557 (.I(itasel[695]),
    .Z(net1557));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1558 (.I(itasel[696]),
    .Z(net1558));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1559 (.I(itasel[697]),
    .Z(net1559));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input156 (.I(itasegm[23]),
    .Z(net156));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1560 (.I(itasel[698]),
    .Z(net1560));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1561 (.I(itasel[699]),
    .Z(net1561));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1562 (.I(itasel[69]),
    .Z(net1562));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 input1563 (.I(itasel[6]),
    .Z(net1563));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1564 (.I(itasel[700]),
    .Z(net1564));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1565 (.I(itasel[701]),
    .Z(net1565));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1566 (.I(itasel[702]),
    .Z(net1566));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1567 (.I(itasel[703]),
    .Z(net1567));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1568 (.I(itasel[704]),
    .Z(net1568));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1569 (.I(itasel[705]),
    .Z(net1569));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input157 (.I(itasegm[240]),
    .Z(net157));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1570 (.I(itasel[706]),
    .Z(net1570));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1571 (.I(itasel[707]),
    .Z(net1571));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1572 (.I(itasel[708]),
    .Z(net1572));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1573 (.I(itasel[709]),
    .Z(net1573));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1574 (.I(itasel[70]),
    .Z(net1574));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1575 (.I(itasel[710]),
    .Z(net1575));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1576 (.I(itasel[711]),
    .Z(net1576));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1577 (.I(itasel[712]),
    .Z(net1577));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1578 (.I(itasel[713]),
    .Z(net1578));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1579 (.I(itasel[714]),
    .Z(net1579));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input158 (.I(itasegm[241]),
    .Z(net158));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1580 (.I(itasel[715]),
    .Z(net1580));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1581 (.I(itasel[716]),
    .Z(net1581));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1582 (.I(itasel[717]),
    .Z(net1582));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1583 (.I(itasel[718]),
    .Z(net1583));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1584 (.I(itasel[719]),
    .Z(net1584));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1585 (.I(itasel[71]),
    .Z(net1585));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1586 (.I(itasel[720]),
    .Z(net1586));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1587 (.I(itasel[721]),
    .Z(net1587));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1588 (.I(itasel[722]),
    .Z(net1588));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1589 (.I(itasel[723]),
    .Z(net1589));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input159 (.I(itasegm[242]),
    .Z(net159));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1590 (.I(itasel[724]),
    .Z(net1590));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1591 (.I(itasel[725]),
    .Z(net1591));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1592 (.I(itasel[726]),
    .Z(net1592));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1593 (.I(itasel[727]),
    .Z(net1593));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1594 (.I(itasel[728]),
    .Z(net1594));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1595 (.I(itasel[729]),
    .Z(net1595));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input1596 (.I(itasel[72]),
    .Z(net1596));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1597 (.I(itasel[730]),
    .Z(net1597));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1598 (.I(itasel[731]),
    .Z(net1598));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1599 (.I(itasel[732]),
    .Z(net1599));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input16 (.I(itasegm[113]),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input160 (.I(itasegm[243]),
    .Z(net160));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1600 (.I(itasel[733]),
    .Z(net1600));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1601 (.I(itasel[734]),
    .Z(net1601));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1602 (.I(itasel[735]),
    .Z(net1602));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1603 (.I(itasel[736]),
    .Z(net1603));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1604 (.I(itasel[737]),
    .Z(net1604));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1605 (.I(itasel[738]),
    .Z(net1605));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1606 (.I(itasel[739]),
    .Z(net1606));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input1607 (.I(itasel[73]),
    .Z(net1607));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1608 (.I(itasel[740]),
    .Z(net1608));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1609 (.I(itasel[741]),
    .Z(net1609));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input161 (.I(itasegm[244]),
    .Z(net161));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1610 (.I(itasel[742]),
    .Z(net1610));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1611 (.I(itasel[743]),
    .Z(net1611));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1612 (.I(itasel[744]),
    .Z(net1612));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1613 (.I(itasel[745]),
    .Z(net1613));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1614 (.I(itasel[746]),
    .Z(net1614));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1615 (.I(itasel[747]),
    .Z(net1615));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1616 (.I(itasel[748]),
    .Z(net1616));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1617 (.I(itasel[749]),
    .Z(net1617));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input1618 (.I(itasel[74]),
    .Z(net1618));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1619 (.I(itasel[750]),
    .Z(net1619));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input162 (.I(itasegm[245]),
    .Z(net162));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1620 (.I(itasel[751]),
    .Z(net1620));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1621 (.I(itasel[752]),
    .Z(net1621));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1622 (.I(itasel[753]),
    .Z(net1622));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1623 (.I(itasel[754]),
    .Z(net1623));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1624 (.I(itasel[755]),
    .Z(net1624));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1625 (.I(itasel[756]),
    .Z(net1625));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1626 (.I(itasel[757]),
    .Z(net1626));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1627 (.I(itasel[758]),
    .Z(net1627));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1628 (.I(itasel[759]),
    .Z(net1628));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input1629 (.I(itasel[75]),
    .Z(net1629));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input163 (.I(itasegm[246]),
    .Z(net163));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1630 (.I(itasel[760]),
    .Z(net1630));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1631 (.I(itasel[761]),
    .Z(net1631));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1632 (.I(itasel[762]),
    .Z(net1632));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1633 (.I(itasel[763]),
    .Z(net1633));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1634 (.I(itasel[764]),
    .Z(net1634));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1635 (.I(itasel[765]),
    .Z(net1635));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1636 (.I(itasel[766]),
    .Z(net1636));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1637 (.I(itasel[767]),
    .Z(net1637));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input1638 (.I(itasel[76]),
    .Z(net1638));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input1639 (.I(itasel[77]),
    .Z(net1639));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input164 (.I(itasegm[247]),
    .Z(net164));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input1640 (.I(itasel[78]),
    .Z(net1640));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input1641 (.I(itasel[79]),
    .Z(net1641));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 input1642 (.I(itasel[7]),
    .Z(net1642));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input1643 (.I(itasel[80]),
    .Z(net1643));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input1644 (.I(itasel[81]),
    .Z(net1644));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input1645 (.I(itasel[82]),
    .Z(net1645));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input1646 (.I(itasel[83]),
    .Z(net1646));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1647 (.I(itasel[84]),
    .Z(net1647));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1648 (.I(itasel[85]),
    .Z(net1648));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1649 (.I(itasel[86]),
    .Z(net1649));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input165 (.I(itasegm[248]),
    .Z(net165));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1650 (.I(itasel[87]),
    .Z(net1650));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1651 (.I(itasel[88]),
    .Z(net1651));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1652 (.I(itasel[89]),
    .Z(net1652));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 input1653 (.I(itasel[8]),
    .Z(net1653));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1654 (.I(itasel[90]),
    .Z(net1654));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1655 (.I(itasel[91]),
    .Z(net1655));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1656 (.I(itasel[92]),
    .Z(net1656));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1657 (.I(itasel[93]),
    .Z(net1657));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1658 (.I(itasel[94]),
    .Z(net1658));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1659 (.I(itasel[95]),
    .Z(net1659));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input166 (.I(itasegm[249]),
    .Z(net166));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1660 (.I(itasel[96]),
    .Z(net1660));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1661 (.I(itasel[97]),
    .Z(net1661));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1662 (.I(itasel[98]),
    .Z(net1662));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1663 (.I(itasel[99]),
    .Z(net1663));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 input1664 (.I(itasel[9]),
    .Z(net1664));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input1665 (.I(nsel[0]),
    .Z(net1665));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input1666 (.I(nsel[1]),
    .Z(net1666));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input1667 (.I(nsel[2]),
    .Z(net1667));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input1668 (.I(nsel[3]),
    .Z(net1668));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 input1669 (.I(nsel[4]),
    .Z(net1669));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input167 (.I(itasegm[24]),
    .Z(net167));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input1670 (.I(nsel[5]),
    .Z(net1670));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input168 (.I(itasegm[250]),
    .Z(net168));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input169 (.I(itasegm[251]),
    .Z(net169));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input17 (.I(itasegm[114]),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input170 (.I(itasegm[252]),
    .Z(net170));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input171 (.I(itasegm[253]),
    .Z(net171));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input172 (.I(itasegm[254]),
    .Z(net172));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input173 (.I(itasegm[255]),
    .Z(net173));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input174 (.I(itasegm[256]),
    .Z(net174));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input175 (.I(itasegm[257]),
    .Z(net175));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input176 (.I(itasegm[258]),
    .Z(net176));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input177 (.I(itasegm[259]),
    .Z(net177));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input178 (.I(itasegm[25]),
    .Z(net178));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input179 (.I(itasegm[260]),
    .Z(net179));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input18 (.I(itasegm[115]),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input180 (.I(itasegm[261]),
    .Z(net180));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input181 (.I(itasegm[262]),
    .Z(net181));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input182 (.I(itasegm[263]),
    .Z(net182));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input183 (.I(itasegm[264]),
    .Z(net183));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input184 (.I(itasegm[265]),
    .Z(net184));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input185 (.I(itasegm[266]),
    .Z(net185));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input186 (.I(itasegm[267]),
    .Z(net186));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input187 (.I(itasegm[268]),
    .Z(net187));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input188 (.I(itasegm[269]),
    .Z(net188));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input189 (.I(itasegm[26]),
    .Z(net189));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input19 (.I(itasegm[116]),
    .Z(net19));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input190 (.I(itasegm[270]),
    .Z(net190));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input191 (.I(itasegm[271]),
    .Z(net191));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input192 (.I(itasegm[272]),
    .Z(net192));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input193 (.I(itasegm[273]),
    .Z(net193));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input194 (.I(itasegm[274]),
    .Z(net194));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input195 (.I(itasegm[275]),
    .Z(net195));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input196 (.I(itasegm[276]),
    .Z(net196));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input197 (.I(itasegm[277]),
    .Z(net197));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input198 (.I(itasegm[278]),
    .Z(net198));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input199 (.I(itasegm[279]),
    .Z(net199));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input2 (.I(itasegm[100]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input20 (.I(itasegm[117]),
    .Z(net20));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input200 (.I(itasegm[27]),
    .Z(net200));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input201 (.I(itasegm[280]),
    .Z(net201));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input202 (.I(itasegm[281]),
    .Z(net202));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input203 (.I(itasegm[282]),
    .Z(net203));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input204 (.I(itasegm[283]),
    .Z(net204));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input205 (.I(itasegm[284]),
    .Z(net205));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input206 (.I(itasegm[285]),
    .Z(net206));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input207 (.I(itasegm[286]),
    .Z(net207));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input208 (.I(itasegm[287]),
    .Z(net208));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input209 (.I(itasegm[288]),
    .Z(net209));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input21 (.I(itasegm[118]),
    .Z(net21));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input210 (.I(itasegm[289]),
    .Z(net210));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input211 (.I(itasegm[28]),
    .Z(net211));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input212 (.I(itasegm[290]),
    .Z(net212));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input213 (.I(itasegm[291]),
    .Z(net213));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input214 (.I(itasegm[292]),
    .Z(net214));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input215 (.I(itasegm[293]),
    .Z(net215));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input216 (.I(itasegm[294]),
    .Z(net216));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input217 (.I(itasegm[295]),
    .Z(net217));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input218 (.I(itasegm[296]),
    .Z(net218));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input219 (.I(itasegm[297]),
    .Z(net219));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input22 (.I(itasegm[119]),
    .Z(net22));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input220 (.I(itasegm[298]),
    .Z(net220));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input221 (.I(itasegm[299]),
    .Z(net221));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input222 (.I(itasegm[29]),
    .Z(net222));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input223 (.I(itasegm[2]),
    .Z(net223));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input224 (.I(itasegm[300]),
    .Z(net224));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input225 (.I(itasegm[301]),
    .Z(net225));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input226 (.I(itasegm[302]),
    .Z(net226));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input227 (.I(itasegm[303]),
    .Z(net227));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input228 (.I(itasegm[304]),
    .Z(net228));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input229 (.I(itasegm[305]),
    .Z(net229));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input23 (.I(itasegm[11]),
    .Z(net23));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input230 (.I(itasegm[306]),
    .Z(net230));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input231 (.I(itasegm[307]),
    .Z(net231));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input232 (.I(itasegm[308]),
    .Z(net232));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input233 (.I(itasegm[309]),
    .Z(net233));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input234 (.I(itasegm[30]),
    .Z(net234));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input235 (.I(itasegm[310]),
    .Z(net235));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input236 (.I(itasegm[311]),
    .Z(net236));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input237 (.I(itasegm[312]),
    .Z(net237));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input238 (.I(itasegm[313]),
    .Z(net238));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input239 (.I(itasegm[314]),
    .Z(net239));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input24 (.I(itasegm[120]),
    .Z(net24));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input240 (.I(itasegm[315]),
    .Z(net240));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input241 (.I(itasegm[316]),
    .Z(net241));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input242 (.I(itasegm[317]),
    .Z(net242));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input243 (.I(itasegm[318]),
    .Z(net243));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input244 (.I(itasegm[319]),
    .Z(net244));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input245 (.I(itasegm[31]),
    .Z(net245));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input246 (.I(itasegm[320]),
    .Z(net246));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input247 (.I(itasegm[321]),
    .Z(net247));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input248 (.I(itasegm[322]),
    .Z(net248));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input249 (.I(itasegm[323]),
    .Z(net249));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input25 (.I(itasegm[121]),
    .Z(net25));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input250 (.I(itasegm[324]),
    .Z(net250));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input251 (.I(itasegm[325]),
    .Z(net251));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input252 (.I(itasegm[326]),
    .Z(net252));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input253 (.I(itasegm[327]),
    .Z(net253));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input254 (.I(itasegm[328]),
    .Z(net254));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input255 (.I(itasegm[329]),
    .Z(net255));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input256 (.I(itasegm[32]),
    .Z(net256));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input257 (.I(itasegm[330]),
    .Z(net257));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input258 (.I(itasegm[331]),
    .Z(net258));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input259 (.I(itasegm[332]),
    .Z(net259));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input26 (.I(itasegm[122]),
    .Z(net26));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input260 (.I(itasegm[333]),
    .Z(net260));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input261 (.I(itasegm[334]),
    .Z(net261));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input262 (.I(itasegm[335]),
    .Z(net262));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input263 (.I(itasegm[336]),
    .Z(net263));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input264 (.I(itasegm[337]),
    .Z(net264));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input265 (.I(itasegm[338]),
    .Z(net265));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input266 (.I(itasegm[339]),
    .Z(net266));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input267 (.I(itasegm[33]),
    .Z(net267));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input268 (.I(itasegm[340]),
    .Z(net268));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input269 (.I(itasegm[341]),
    .Z(net269));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input27 (.I(itasegm[123]),
    .Z(net27));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input270 (.I(itasegm[342]),
    .Z(net270));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input271 (.I(itasegm[343]),
    .Z(net271));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input272 (.I(itasegm[344]),
    .Z(net272));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input273 (.I(itasegm[345]),
    .Z(net273));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input274 (.I(itasegm[346]),
    .Z(net274));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input275 (.I(itasegm[347]),
    .Z(net275));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input276 (.I(itasegm[348]),
    .Z(net276));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input277 (.I(itasegm[349]),
    .Z(net277));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input278 (.I(itasegm[34]),
    .Z(net278));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input279 (.I(itasegm[350]),
    .Z(net279));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input28 (.I(itasegm[124]),
    .Z(net28));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input280 (.I(itasegm[351]),
    .Z(net280));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input281 (.I(itasegm[352]),
    .Z(net281));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input282 (.I(itasegm[353]),
    .Z(net282));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input283 (.I(itasegm[354]),
    .Z(net283));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input284 (.I(itasegm[355]),
    .Z(net284));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input285 (.I(itasegm[356]),
    .Z(net285));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input286 (.I(itasegm[357]),
    .Z(net286));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input287 (.I(itasegm[358]),
    .Z(net287));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input288 (.I(itasegm[359]),
    .Z(net288));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input289 (.I(itasegm[35]),
    .Z(net289));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input29 (.I(itasegm[125]),
    .Z(net29));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input290 (.I(itasegm[360]),
    .Z(net290));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input291 (.I(itasegm[361]),
    .Z(net291));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input292 (.I(itasegm[362]),
    .Z(net292));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input293 (.I(itasegm[363]),
    .Z(net293));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input294 (.I(itasegm[364]),
    .Z(net294));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input295 (.I(itasegm[365]),
    .Z(net295));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input296 (.I(itasegm[366]),
    .Z(net296));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input297 (.I(itasegm[367]),
    .Z(net297));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input298 (.I(itasegm[368]),
    .Z(net298));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input299 (.I(itasegm[369]),
    .Z(net299));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input3 (.I(itasegm[101]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input30 (.I(itasegm[126]),
    .Z(net30));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input300 (.I(itasegm[36]),
    .Z(net300));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input301 (.I(itasegm[370]),
    .Z(net301));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input302 (.I(itasegm[371]),
    .Z(net302));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input303 (.I(itasegm[372]),
    .Z(net303));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input304 (.I(itasegm[373]),
    .Z(net304));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input305 (.I(itasegm[374]),
    .Z(net305));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input306 (.I(itasegm[375]),
    .Z(net306));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input307 (.I(itasegm[376]),
    .Z(net307));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 input308 (.I(itasegm[377]),
    .Z(net308));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input309 (.I(itasegm[378]),
    .Z(net309));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input31 (.I(itasegm[127]),
    .Z(net31));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input310 (.I(itasegm[379]),
    .Z(net310));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input311 (.I(itasegm[37]),
    .Z(net311));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input312 (.I(itasegm[380]),
    .Z(net312));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input313 (.I(itasegm[381]),
    .Z(net313));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input314 (.I(itasegm[382]),
    .Z(net314));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input315 (.I(itasegm[383]),
    .Z(net315));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input316 (.I(itasegm[384]),
    .Z(net316));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input317 (.I(itasegm[385]),
    .Z(net317));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input318 (.I(itasegm[386]),
    .Z(net318));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input319 (.I(itasegm[387]),
    .Z(net319));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input32 (.I(itasegm[128]),
    .Z(net32));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input320 (.I(itasegm[388]),
    .Z(net320));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input321 (.I(itasegm[389]),
    .Z(net321));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input322 (.I(itasegm[38]),
    .Z(net322));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input323 (.I(itasegm[390]),
    .Z(net323));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input324 (.I(itasegm[391]),
    .Z(net324));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input325 (.I(itasegm[392]),
    .Z(net325));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input326 (.I(itasegm[393]),
    .Z(net326));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input327 (.I(itasegm[394]),
    .Z(net327));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input328 (.I(itasegm[395]),
    .Z(net328));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input329 (.I(itasegm[396]),
    .Z(net329));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input33 (.I(itasegm[129]),
    .Z(net33));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input330 (.I(itasegm[397]),
    .Z(net330));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input331 (.I(itasegm[398]),
    .Z(net331));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input332 (.I(itasegm[399]),
    .Z(net332));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input333 (.I(itasegm[39]),
    .Z(net333));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input334 (.I(itasegm[3]),
    .Z(net334));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input335 (.I(itasegm[400]),
    .Z(net335));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input336 (.I(itasegm[401]),
    .Z(net336));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input337 (.I(itasegm[402]),
    .Z(net337));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input338 (.I(itasegm[403]),
    .Z(net338));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input339 (.I(itasegm[404]),
    .Z(net339));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input34 (.I(itasegm[12]),
    .Z(net34));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input340 (.I(itasegm[405]),
    .Z(net340));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input341 (.I(itasegm[406]),
    .Z(net341));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input342 (.I(itasegm[407]),
    .Z(net342));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input343 (.I(itasegm[408]),
    .Z(net343));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input344 (.I(itasegm[409]),
    .Z(net344));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input345 (.I(itasegm[40]),
    .Z(net345));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input346 (.I(itasegm[410]),
    .Z(net346));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input347 (.I(itasegm[411]),
    .Z(net347));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input348 (.I(itasegm[412]),
    .Z(net348));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input349 (.I(itasegm[413]),
    .Z(net349));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input35 (.I(itasegm[130]),
    .Z(net35));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input350 (.I(itasegm[414]),
    .Z(net350));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input351 (.I(itasegm[415]),
    .Z(net351));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input352 (.I(itasegm[416]),
    .Z(net352));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input353 (.I(itasegm[417]),
    .Z(net353));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input354 (.I(itasegm[418]),
    .Z(net354));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input355 (.I(itasegm[419]),
    .Z(net355));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input356 (.I(itasegm[41]),
    .Z(net356));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input357 (.I(itasegm[420]),
    .Z(net357));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input358 (.I(itasegm[421]),
    .Z(net358));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input359 (.I(itasegm[422]),
    .Z(net359));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input36 (.I(itasegm[131]),
    .Z(net36));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input360 (.I(itasegm[423]),
    .Z(net360));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input361 (.I(itasegm[424]),
    .Z(net361));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input362 (.I(itasegm[425]),
    .Z(net362));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input363 (.I(itasegm[426]),
    .Z(net363));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input364 (.I(itasegm[427]),
    .Z(net364));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input365 (.I(itasegm[428]),
    .Z(net365));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input366 (.I(itasegm[429]),
    .Z(net366));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input367 (.I(itasegm[42]),
    .Z(net367));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input368 (.I(itasegm[430]),
    .Z(net368));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input369 (.I(itasegm[431]),
    .Z(net369));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input37 (.I(itasegm[132]),
    .Z(net37));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input370 (.I(itasegm[432]),
    .Z(net370));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input371 (.I(itasegm[433]),
    .Z(net371));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input372 (.I(itasegm[434]),
    .Z(net372));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input373 (.I(itasegm[435]),
    .Z(net373));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input374 (.I(itasegm[436]),
    .Z(net374));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input375 (.I(itasegm[437]),
    .Z(net375));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input376 (.I(itasegm[438]),
    .Z(net376));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input377 (.I(itasegm[439]),
    .Z(net377));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input378 (.I(itasegm[43]),
    .Z(net378));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input379 (.I(itasegm[440]),
    .Z(net379));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input38 (.I(itasegm[133]),
    .Z(net38));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input380 (.I(itasegm[441]),
    .Z(net380));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input381 (.I(itasegm[442]),
    .Z(net381));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input382 (.I(itasegm[443]),
    .Z(net382));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input383 (.I(itasegm[444]),
    .Z(net383));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input384 (.I(itasegm[445]),
    .Z(net384));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input385 (.I(itasegm[446]),
    .Z(net385));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input386 (.I(itasegm[447]),
    .Z(net386));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input387 (.I(itasegm[448]),
    .Z(net387));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input388 (.I(itasegm[449]),
    .Z(net388));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input389 (.I(itasegm[44]),
    .Z(net389));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input39 (.I(itasegm[134]),
    .Z(net39));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input390 (.I(itasegm[450]),
    .Z(net390));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input391 (.I(itasegm[451]),
    .Z(net391));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input392 (.I(itasegm[452]),
    .Z(net392));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input393 (.I(itasegm[453]),
    .Z(net393));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input394 (.I(itasegm[454]),
    .Z(net394));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input395 (.I(itasegm[455]),
    .Z(net395));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input396 (.I(itasegm[456]),
    .Z(net396));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input397 (.I(itasegm[457]),
    .Z(net397));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input398 (.I(itasegm[458]),
    .Z(net398));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input399 (.I(itasegm[459]),
    .Z(net399));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input4 (.I(itasegm[102]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input40 (.I(itasegm[135]),
    .Z(net40));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input400 (.I(itasegm[45]),
    .Z(net400));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input401 (.I(itasegm[460]),
    .Z(net401));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input402 (.I(itasegm[461]),
    .Z(net402));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input403 (.I(itasegm[462]),
    .Z(net403));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input404 (.I(itasegm[463]),
    .Z(net404));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input405 (.I(itasegm[464]),
    .Z(net405));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input406 (.I(itasegm[465]),
    .Z(net406));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input407 (.I(itasegm[466]),
    .Z(net407));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input408 (.I(itasegm[467]),
    .Z(net408));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input409 (.I(itasegm[468]),
    .Z(net409));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input41 (.I(itasegm[136]),
    .Z(net41));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input410 (.I(itasegm[469]),
    .Z(net410));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input411 (.I(itasegm[46]),
    .Z(net411));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input412 (.I(itasegm[470]),
    .Z(net412));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input413 (.I(itasegm[471]),
    .Z(net413));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input414 (.I(itasegm[472]),
    .Z(net414));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input415 (.I(itasegm[473]),
    .Z(net415));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input416 (.I(itasegm[474]),
    .Z(net416));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input417 (.I(itasegm[475]),
    .Z(net417));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input418 (.I(itasegm[476]),
    .Z(net418));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input419 (.I(itasegm[477]),
    .Z(net419));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input42 (.I(itasegm[137]),
    .Z(net42));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input420 (.I(itasegm[478]),
    .Z(net420));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input421 (.I(itasegm[479]),
    .Z(net421));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input422 (.I(itasegm[47]),
    .Z(net422));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input423 (.I(itasegm[480]),
    .Z(net423));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input424 (.I(itasegm[481]),
    .Z(net424));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input425 (.I(itasegm[482]),
    .Z(net425));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input426 (.I(itasegm[483]),
    .Z(net426));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input427 (.I(itasegm[484]),
    .Z(net427));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input428 (.I(itasegm[485]),
    .Z(net428));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input429 (.I(itasegm[486]),
    .Z(net429));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input43 (.I(itasegm[138]),
    .Z(net43));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input430 (.I(itasegm[487]),
    .Z(net430));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input431 (.I(itasegm[488]),
    .Z(net431));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input432 (.I(itasegm[489]),
    .Z(net432));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input433 (.I(itasegm[48]),
    .Z(net433));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input434 (.I(itasegm[490]),
    .Z(net434));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input435 (.I(itasegm[491]),
    .Z(net435));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input436 (.I(itasegm[492]),
    .Z(net436));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input437 (.I(itasegm[493]),
    .Z(net437));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input438 (.I(itasegm[494]),
    .Z(net438));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input439 (.I(itasegm[495]),
    .Z(net439));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input44 (.I(itasegm[139]),
    .Z(net44));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input440 (.I(itasegm[496]),
    .Z(net440));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input441 (.I(itasegm[497]),
    .Z(net441));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input442 (.I(itasegm[498]),
    .Z(net442));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input443 (.I(itasegm[499]),
    .Z(net443));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input444 (.I(itasegm[49]),
    .Z(net444));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input445 (.I(itasegm[4]),
    .Z(net445));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input446 (.I(itasegm[500]),
    .Z(net446));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input447 (.I(itasegm[501]),
    .Z(net447));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input448 (.I(itasegm[502]),
    .Z(net448));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input449 (.I(itasegm[503]),
    .Z(net449));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input45 (.I(itasegm[13]),
    .Z(net45));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input450 (.I(itasegm[504]),
    .Z(net450));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input451 (.I(itasegm[505]),
    .Z(net451));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input452 (.I(itasegm[506]),
    .Z(net452));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input453 (.I(itasegm[507]),
    .Z(net453));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input454 (.I(itasegm[508]),
    .Z(net454));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input455 (.I(itasegm[509]),
    .Z(net455));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input456 (.I(itasegm[50]),
    .Z(net456));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input457 (.I(itasegm[510]),
    .Z(net457));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input458 (.I(itasegm[511]),
    .Z(net458));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input459 (.I(itasegm[512]),
    .Z(net459));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input46 (.I(itasegm[140]),
    .Z(net46));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input460 (.I(itasegm[513]),
    .Z(net460));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input461 (.I(itasegm[514]),
    .Z(net461));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input462 (.I(itasegm[515]),
    .Z(net462));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input463 (.I(itasegm[516]),
    .Z(net463));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input464 (.I(itasegm[517]),
    .Z(net464));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input465 (.I(itasegm[518]),
    .Z(net465));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input466 (.I(itasegm[519]),
    .Z(net466));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input467 (.I(itasegm[51]),
    .Z(net467));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input468 (.I(itasegm[520]),
    .Z(net468));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input469 (.I(itasegm[521]),
    .Z(net469));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input47 (.I(itasegm[141]),
    .Z(net47));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input470 (.I(itasegm[522]),
    .Z(net470));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input471 (.I(itasegm[523]),
    .Z(net471));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input472 (.I(itasegm[524]),
    .Z(net472));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input473 (.I(itasegm[525]),
    .Z(net473));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input474 (.I(itasegm[526]),
    .Z(net474));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input475 (.I(itasegm[527]),
    .Z(net475));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input476 (.I(itasegm[528]),
    .Z(net476));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input477 (.I(itasegm[529]),
    .Z(net477));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input478 (.I(itasegm[52]),
    .Z(net478));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input479 (.I(itasegm[530]),
    .Z(net479));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input48 (.I(itasegm[142]),
    .Z(net48));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input480 (.I(itasegm[531]),
    .Z(net480));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input481 (.I(itasegm[532]),
    .Z(net481));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input482 (.I(itasegm[533]),
    .Z(net482));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input483 (.I(itasegm[534]),
    .Z(net483));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input484 (.I(itasegm[535]),
    .Z(net484));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input485 (.I(itasegm[536]),
    .Z(net485));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input486 (.I(itasegm[537]),
    .Z(net486));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input487 (.I(itasegm[538]),
    .Z(net487));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input488 (.I(itasegm[539]),
    .Z(net488));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input489 (.I(itasegm[53]),
    .Z(net489));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input49 (.I(itasegm[143]),
    .Z(net49));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input490 (.I(itasegm[540]),
    .Z(net490));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input491 (.I(itasegm[541]),
    .Z(net491));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input492 (.I(itasegm[542]),
    .Z(net492));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input493 (.I(itasegm[543]),
    .Z(net493));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input494 (.I(itasegm[544]),
    .Z(net494));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input495 (.I(itasegm[545]),
    .Z(net495));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input496 (.I(itasegm[546]),
    .Z(net496));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input497 (.I(itasegm[547]),
    .Z(net497));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input498 (.I(itasegm[548]),
    .Z(net498));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input499 (.I(itasegm[549]),
    .Z(net499));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input5 (.I(itasegm[103]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input50 (.I(itasegm[144]),
    .Z(net50));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input500 (.I(itasegm[54]),
    .Z(net500));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input501 (.I(itasegm[550]),
    .Z(net501));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input502 (.I(itasegm[551]),
    .Z(net502));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input503 (.I(itasegm[552]),
    .Z(net503));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input504 (.I(itasegm[553]),
    .Z(net504));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input505 (.I(itasegm[554]),
    .Z(net505));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input506 (.I(itasegm[555]),
    .Z(net506));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input507 (.I(itasegm[556]),
    .Z(net507));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input508 (.I(itasegm[557]),
    .Z(net508));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input509 (.I(itasegm[558]),
    .Z(net509));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input51 (.I(itasegm[145]),
    .Z(net51));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input510 (.I(itasegm[559]),
    .Z(net510));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input511 (.I(itasegm[55]),
    .Z(net511));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input512 (.I(itasegm[560]),
    .Z(net512));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input513 (.I(itasegm[561]),
    .Z(net513));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input514 (.I(itasegm[562]),
    .Z(net514));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input515 (.I(itasegm[563]),
    .Z(net515));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input516 (.I(itasegm[564]),
    .Z(net516));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input517 (.I(itasegm[565]),
    .Z(net517));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input518 (.I(itasegm[566]),
    .Z(net518));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input519 (.I(itasegm[567]),
    .Z(net519));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input52 (.I(itasegm[146]),
    .Z(net52));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input520 (.I(itasegm[568]),
    .Z(net520));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input521 (.I(itasegm[569]),
    .Z(net521));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input522 (.I(itasegm[56]),
    .Z(net522));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input523 (.I(itasegm[570]),
    .Z(net523));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input524 (.I(itasegm[571]),
    .Z(net524));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input525 (.I(itasegm[572]),
    .Z(net525));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input526 (.I(itasegm[573]),
    .Z(net526));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input527 (.I(itasegm[574]),
    .Z(net527));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input528 (.I(itasegm[575]),
    .Z(net528));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input529 (.I(itasegm[576]),
    .Z(net529));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input53 (.I(itasegm[147]),
    .Z(net53));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input530 (.I(itasegm[577]),
    .Z(net530));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input531 (.I(itasegm[578]),
    .Z(net531));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input532 (.I(itasegm[579]),
    .Z(net532));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input533 (.I(itasegm[57]),
    .Z(net533));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input534 (.I(itasegm[580]),
    .Z(net534));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input535 (.I(itasegm[581]),
    .Z(net535));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input536 (.I(itasegm[582]),
    .Z(net536));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input537 (.I(itasegm[583]),
    .Z(net537));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input538 (.I(itasegm[584]),
    .Z(net538));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input539 (.I(itasegm[585]),
    .Z(net539));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input54 (.I(itasegm[148]),
    .Z(net54));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input540 (.I(itasegm[586]),
    .Z(net540));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input541 (.I(itasegm[587]),
    .Z(net541));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input542 (.I(itasegm[588]),
    .Z(net542));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input543 (.I(itasegm[589]),
    .Z(net543));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input544 (.I(itasegm[58]),
    .Z(net544));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input545 (.I(itasegm[590]),
    .Z(net545));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input546 (.I(itasegm[591]),
    .Z(net546));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input547 (.I(itasegm[592]),
    .Z(net547));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input548 (.I(itasegm[593]),
    .Z(net548));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input549 (.I(itasegm[594]),
    .Z(net549));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input55 (.I(itasegm[149]),
    .Z(net55));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input550 (.I(itasegm[595]),
    .Z(net550));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input551 (.I(itasegm[596]),
    .Z(net551));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input552 (.I(itasegm[597]),
    .Z(net552));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input553 (.I(itasegm[598]),
    .Z(net553));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input554 (.I(itasegm[599]),
    .Z(net554));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input555 (.I(itasegm[59]),
    .Z(net555));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input556 (.I(itasegm[5]),
    .Z(net556));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input557 (.I(itasegm[600]),
    .Z(net557));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input558 (.I(itasegm[601]),
    .Z(net558));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input559 (.I(itasegm[602]),
    .Z(net559));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input56 (.I(itasegm[14]),
    .Z(net56));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input560 (.I(itasegm[603]),
    .Z(net560));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input561 (.I(itasegm[604]),
    .Z(net561));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input562 (.I(itasegm[605]),
    .Z(net562));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input563 (.I(itasegm[606]),
    .Z(net563));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input564 (.I(itasegm[607]),
    .Z(net564));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input565 (.I(itasegm[608]),
    .Z(net565));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input566 (.I(itasegm[609]),
    .Z(net566));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input567 (.I(itasegm[60]),
    .Z(net567));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input568 (.I(itasegm[610]),
    .Z(net568));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input569 (.I(itasegm[611]),
    .Z(net569));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input57 (.I(itasegm[150]),
    .Z(net57));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input570 (.I(itasegm[612]),
    .Z(net570));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input571 (.I(itasegm[613]),
    .Z(net571));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input572 (.I(itasegm[614]),
    .Z(net572));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input573 (.I(itasegm[615]),
    .Z(net573));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input574 (.I(itasegm[616]),
    .Z(net574));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input575 (.I(itasegm[617]),
    .Z(net575));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input576 (.I(itasegm[618]),
    .Z(net576));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input577 (.I(itasegm[619]),
    .Z(net577));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input578 (.I(itasegm[61]),
    .Z(net578));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input579 (.I(itasegm[620]),
    .Z(net579));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input58 (.I(itasegm[151]),
    .Z(net58));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input580 (.I(itasegm[621]),
    .Z(net580));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input581 (.I(itasegm[622]),
    .Z(net581));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input582 (.I(itasegm[623]),
    .Z(net582));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input583 (.I(itasegm[624]),
    .Z(net583));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input584 (.I(itasegm[625]),
    .Z(net584));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input585 (.I(itasegm[626]),
    .Z(net585));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input586 (.I(itasegm[627]),
    .Z(net586));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input587 (.I(itasegm[628]),
    .Z(net587));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input588 (.I(itasegm[629]),
    .Z(net588));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input589 (.I(itasegm[62]),
    .Z(net589));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input59 (.I(itasegm[152]),
    .Z(net59));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input590 (.I(itasegm[630]),
    .Z(net590));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input591 (.I(itasegm[631]),
    .Z(net591));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input592 (.I(itasegm[632]),
    .Z(net592));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input593 (.I(itasegm[633]),
    .Z(net593));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input594 (.I(itasegm[634]),
    .Z(net594));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input595 (.I(itasegm[635]),
    .Z(net595));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input596 (.I(itasegm[636]),
    .Z(net596));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input597 (.I(itasegm[637]),
    .Z(net597));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input598 (.I(itasegm[638]),
    .Z(net598));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input599 (.I(itasegm[639]),
    .Z(net599));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input6 (.I(itasegm[104]),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input60 (.I(itasegm[153]),
    .Z(net60));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input600 (.I(itasegm[63]),
    .Z(net600));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input601 (.I(itasegm[640]),
    .Z(net601));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input602 (.I(itasegm[641]),
    .Z(net602));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input603 (.I(itasegm[642]),
    .Z(net603));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input604 (.I(itasegm[643]),
    .Z(net604));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input605 (.I(itasegm[644]),
    .Z(net605));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input606 (.I(itasegm[645]),
    .Z(net606));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input607 (.I(itasegm[646]),
    .Z(net607));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input608 (.I(itasegm[647]),
    .Z(net608));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input609 (.I(itasegm[648]),
    .Z(net609));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input61 (.I(itasegm[154]),
    .Z(net61));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input610 (.I(itasegm[649]),
    .Z(net610));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input611 (.I(itasegm[64]),
    .Z(net611));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input612 (.I(itasegm[650]),
    .Z(net612));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input613 (.I(itasegm[651]),
    .Z(net613));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input614 (.I(itasegm[652]),
    .Z(net614));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input615 (.I(itasegm[653]),
    .Z(net615));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input616 (.I(itasegm[654]),
    .Z(net616));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input617 (.I(itasegm[655]),
    .Z(net617));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input618 (.I(itasegm[656]),
    .Z(net618));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input619 (.I(itasegm[657]),
    .Z(net619));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input62 (.I(itasegm[155]),
    .Z(net62));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input620 (.I(itasegm[658]),
    .Z(net620));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input621 (.I(itasegm[659]),
    .Z(net621));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input622 (.I(itasegm[65]),
    .Z(net622));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input623 (.I(itasegm[660]),
    .Z(net623));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input624 (.I(itasegm[661]),
    .Z(net624));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input625 (.I(itasegm[662]),
    .Z(net625));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input626 (.I(itasegm[663]),
    .Z(net626));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input627 (.I(itasegm[664]),
    .Z(net627));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input628 (.I(itasegm[665]),
    .Z(net628));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input629 (.I(itasegm[666]),
    .Z(net629));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input63 (.I(itasegm[156]),
    .Z(net63));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input630 (.I(itasegm[667]),
    .Z(net630));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input631 (.I(itasegm[668]),
    .Z(net631));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input632 (.I(itasegm[669]),
    .Z(net632));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input633 (.I(itasegm[66]),
    .Z(net633));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input634 (.I(itasegm[670]),
    .Z(net634));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input635 (.I(itasegm[671]),
    .Z(net635));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input636 (.I(itasegm[672]),
    .Z(net636));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input637 (.I(itasegm[673]),
    .Z(net637));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input638 (.I(itasegm[674]),
    .Z(net638));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input639 (.I(itasegm[675]),
    .Z(net639));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input64 (.I(itasegm[157]),
    .Z(net64));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input640 (.I(itasegm[676]),
    .Z(net640));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input641 (.I(itasegm[677]),
    .Z(net641));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input642 (.I(itasegm[678]),
    .Z(net642));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input643 (.I(itasegm[679]),
    .Z(net643));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input644 (.I(itasegm[67]),
    .Z(net644));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input645 (.I(itasegm[680]),
    .Z(net645));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input646 (.I(itasegm[681]),
    .Z(net646));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input647 (.I(itasegm[682]),
    .Z(net647));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input648 (.I(itasegm[683]),
    .Z(net648));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input649 (.I(itasegm[684]),
    .Z(net649));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input65 (.I(itasegm[158]),
    .Z(net65));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input650 (.I(itasegm[685]),
    .Z(net650));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input651 (.I(itasegm[686]),
    .Z(net651));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input652 (.I(itasegm[687]),
    .Z(net652));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input653 (.I(itasegm[688]),
    .Z(net653));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input654 (.I(itasegm[689]),
    .Z(net654));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input655 (.I(itasegm[68]),
    .Z(net655));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input656 (.I(itasegm[690]),
    .Z(net656));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input657 (.I(itasegm[691]),
    .Z(net657));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input658 (.I(itasegm[692]),
    .Z(net658));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input659 (.I(itasegm[693]),
    .Z(net659));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input66 (.I(itasegm[159]),
    .Z(net66));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input660 (.I(itasegm[694]),
    .Z(net660));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input661 (.I(itasegm[695]),
    .Z(net661));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input662 (.I(itasegm[696]),
    .Z(net662));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input663 (.I(itasegm[697]),
    .Z(net663));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input664 (.I(itasegm[698]),
    .Z(net664));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input665 (.I(itasegm[699]),
    .Z(net665));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input666 (.I(itasegm[69]),
    .Z(net666));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input667 (.I(itasegm[6]),
    .Z(net667));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input668 (.I(itasegm[700]),
    .Z(net668));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input669 (.I(itasegm[701]),
    .Z(net669));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input67 (.I(itasegm[15]),
    .Z(net67));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input670 (.I(itasegm[702]),
    .Z(net670));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input671 (.I(itasegm[703]),
    .Z(net671));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input672 (.I(itasegm[704]),
    .Z(net672));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input673 (.I(itasegm[705]),
    .Z(net673));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input674 (.I(itasegm[706]),
    .Z(net674));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input675 (.I(itasegm[707]),
    .Z(net675));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input676 (.I(itasegm[708]),
    .Z(net676));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input677 (.I(itasegm[709]),
    .Z(net677));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input678 (.I(itasegm[70]),
    .Z(net678));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input679 (.I(itasegm[710]),
    .Z(net679));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input68 (.I(itasegm[160]),
    .Z(net68));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input680 (.I(itasegm[711]),
    .Z(net680));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input681 (.I(itasegm[712]),
    .Z(net681));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input682 (.I(itasegm[713]),
    .Z(net682));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input683 (.I(itasegm[714]),
    .Z(net683));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input684 (.I(itasegm[715]),
    .Z(net684));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input685 (.I(itasegm[716]),
    .Z(net685));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input686 (.I(itasegm[717]),
    .Z(net686));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input687 (.I(itasegm[718]),
    .Z(net687));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input688 (.I(itasegm[719]),
    .Z(net688));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input689 (.I(itasegm[71]),
    .Z(net689));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input69 (.I(itasegm[161]),
    .Z(net69));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input690 (.I(itasegm[720]),
    .Z(net690));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input691 (.I(itasegm[721]),
    .Z(net691));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input692 (.I(itasegm[722]),
    .Z(net692));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input693 (.I(itasegm[723]),
    .Z(net693));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input694 (.I(itasegm[724]),
    .Z(net694));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input695 (.I(itasegm[725]),
    .Z(net695));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input696 (.I(itasegm[726]),
    .Z(net696));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input697 (.I(itasegm[727]),
    .Z(net697));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input698 (.I(itasegm[728]),
    .Z(net698));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input699 (.I(itasegm[729]),
    .Z(net699));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input7 (.I(itasegm[105]),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input70 (.I(itasegm[162]),
    .Z(net70));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input700 (.I(itasegm[72]),
    .Z(net700));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input701 (.I(itasegm[730]),
    .Z(net701));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input702 (.I(itasegm[731]),
    .Z(net702));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input703 (.I(itasegm[732]),
    .Z(net703));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input704 (.I(itasegm[733]),
    .Z(net704));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input705 (.I(itasegm[734]),
    .Z(net705));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input706 (.I(itasegm[735]),
    .Z(net706));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input707 (.I(itasegm[736]),
    .Z(net707));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input708 (.I(itasegm[737]),
    .Z(net708));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input709 (.I(itasegm[738]),
    .Z(net709));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input71 (.I(itasegm[163]),
    .Z(net71));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input710 (.I(itasegm[739]),
    .Z(net710));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input711 (.I(itasegm[73]),
    .Z(net711));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input712 (.I(itasegm[740]),
    .Z(net712));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input713 (.I(itasegm[741]),
    .Z(net713));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input714 (.I(itasegm[742]),
    .Z(net714));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input715 (.I(itasegm[743]),
    .Z(net715));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input716 (.I(itasegm[744]),
    .Z(net716));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input717 (.I(itasegm[745]),
    .Z(net717));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input718 (.I(itasegm[746]),
    .Z(net718));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input719 (.I(itasegm[747]),
    .Z(net719));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input72 (.I(itasegm[164]),
    .Z(net72));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input720 (.I(itasegm[748]),
    .Z(net720));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input721 (.I(itasegm[749]),
    .Z(net721));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input722 (.I(itasegm[74]),
    .Z(net722));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input723 (.I(itasegm[750]),
    .Z(net723));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input724 (.I(itasegm[751]),
    .Z(net724));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input725 (.I(itasegm[752]),
    .Z(net725));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input726 (.I(itasegm[753]),
    .Z(net726));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input727 (.I(itasegm[754]),
    .Z(net727));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input728 (.I(itasegm[755]),
    .Z(net728));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 input729 (.I(itasegm[756]),
    .Z(net729));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input73 (.I(itasegm[165]),
    .Z(net73));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 input730 (.I(itasegm[757]),
    .Z(net730));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input731 (.I(itasegm[758]),
    .Z(net731));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input732 (.I(itasegm[759]),
    .Z(net732));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input733 (.I(itasegm[75]),
    .Z(net733));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input734 (.I(itasegm[760]),
    .Z(net734));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 input735 (.I(itasegm[761]),
    .Z(net735));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input736 (.I(itasegm[762]),
    .Z(net736));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input737 (.I(itasegm[763]),
    .Z(net737));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 input738 (.I(itasegm[764]),
    .Z(net738));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input739 (.I(itasegm[765]),
    .Z(net739));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input74 (.I(itasegm[166]),
    .Z(net74));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input740 (.I(itasegm[766]),
    .Z(net740));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input741 (.I(itasegm[767]),
    .Z(net741));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 input742 (.I(itasegm[768]),
    .Z(net742));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input743 (.I(itasegm[769]),
    .Z(net743));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input744 (.I(itasegm[76]),
    .Z(net744));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 input745 (.I(itasegm[770]),
    .Z(net745));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 input746 (.I(itasegm[771]),
    .Z(net746));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 input747 (.I(itasegm[772]),
    .Z(net747));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 input748 (.I(itasegm[773]),
    .Z(net748));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 input749 (.I(itasegm[774]),
    .Z(net749));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input75 (.I(itasegm[167]),
    .Z(net75));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 input750 (.I(itasegm[775]),
    .Z(net750));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 input751 (.I(itasegm[776]),
    .Z(net751));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 input752 (.I(itasegm[777]),
    .Z(net752));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 input753 (.I(itasegm[778]),
    .Z(net753));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 input754 (.I(itasegm[779]),
    .Z(net754));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input755 (.I(itasegm[77]),
    .Z(net755));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 input756 (.I(itasegm[780]),
    .Z(net756));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 input757 (.I(itasegm[781]),
    .Z(net757));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 input758 (.I(itasegm[782]),
    .Z(net758));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 input759 (.I(itasegm[783]),
    .Z(net759));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input76 (.I(itasegm[168]),
    .Z(net76));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input760 (.I(itasegm[784]),
    .Z(net760));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input761 (.I(itasegm[785]),
    .Z(net761));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input762 (.I(itasegm[786]),
    .Z(net762));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input763 (.I(itasegm[787]),
    .Z(net763));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input764 (.I(itasegm[788]),
    .Z(net764));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input765 (.I(itasegm[789]),
    .Z(net765));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input766 (.I(itasegm[78]),
    .Z(net766));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input767 (.I(itasegm[790]),
    .Z(net767));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input768 (.I(itasegm[791]),
    .Z(net768));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input769 (.I(itasegm[792]),
    .Z(net769));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input77 (.I(itasegm[169]),
    .Z(net77));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input770 (.I(itasegm[793]),
    .Z(net770));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input771 (.I(itasegm[794]),
    .Z(net771));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input772 (.I(itasegm[795]),
    .Z(net772));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input773 (.I(itasegm[796]),
    .Z(net773));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input774 (.I(itasegm[797]),
    .Z(net774));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input775 (.I(itasegm[798]),
    .Z(net775));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input776 (.I(itasegm[799]),
    .Z(net776));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input777 (.I(itasegm[79]),
    .Z(net777));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input778 (.I(itasegm[7]),
    .Z(net778));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input779 (.I(itasegm[800]),
    .Z(net779));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input78 (.I(itasegm[16]),
    .Z(net78));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input780 (.I(itasegm[801]),
    .Z(net780));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input781 (.I(itasegm[802]),
    .Z(net781));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input782 (.I(itasegm[803]),
    .Z(net782));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input783 (.I(itasegm[804]),
    .Z(net783));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input784 (.I(itasegm[805]),
    .Z(net784));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input785 (.I(itasegm[806]),
    .Z(net785));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input786 (.I(itasegm[807]),
    .Z(net786));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input787 (.I(itasegm[808]),
    .Z(net787));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input788 (.I(itasegm[809]),
    .Z(net788));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input789 (.I(itasegm[80]),
    .Z(net789));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input79 (.I(itasegm[170]),
    .Z(net79));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input790 (.I(itasegm[810]),
    .Z(net790));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input791 (.I(itasegm[811]),
    .Z(net791));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input792 (.I(itasegm[812]),
    .Z(net792));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input793 (.I(itasegm[813]),
    .Z(net793));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input794 (.I(itasegm[814]),
    .Z(net794));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input795 (.I(itasegm[815]),
    .Z(net795));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input796 (.I(itasegm[816]),
    .Z(net796));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input797 (.I(itasegm[817]),
    .Z(net797));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input798 (.I(itasegm[818]),
    .Z(net798));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input799 (.I(itasegm[819]),
    .Z(net799));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input8 (.I(itasegm[106]),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input80 (.I(itasegm[171]),
    .Z(net80));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input800 (.I(itasegm[81]),
    .Z(net800));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input801 (.I(itasegm[820]),
    .Z(net801));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input802 (.I(itasegm[821]),
    .Z(net802));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input803 (.I(itasegm[822]),
    .Z(net803));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input804 (.I(itasegm[823]),
    .Z(net804));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input805 (.I(itasegm[824]),
    .Z(net805));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input806 (.I(itasegm[825]),
    .Z(net806));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input807 (.I(itasegm[826]),
    .Z(net807));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input808 (.I(itasegm[827]),
    .Z(net808));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input809 (.I(itasegm[828]),
    .Z(net809));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input81 (.I(itasegm[172]),
    .Z(net81));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input810 (.I(itasegm[829]),
    .Z(net810));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input811 (.I(itasegm[82]),
    .Z(net811));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input812 (.I(itasegm[830]),
    .Z(net812));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input813 (.I(itasegm[831]),
    .Z(net813));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input814 (.I(itasegm[832]),
    .Z(net814));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input815 (.I(itasegm[833]),
    .Z(net815));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input816 (.I(itasegm[834]),
    .Z(net816));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input817 (.I(itasegm[835]),
    .Z(net817));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input818 (.I(itasegm[836]),
    .Z(net818));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input819 (.I(itasegm[837]),
    .Z(net819));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input82 (.I(itasegm[173]),
    .Z(net82));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input820 (.I(itasegm[838]),
    .Z(net820));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input821 (.I(itasegm[839]),
    .Z(net821));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input822 (.I(itasegm[83]),
    .Z(net822));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input823 (.I(itasegm[840]),
    .Z(net823));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input824 (.I(itasegm[841]),
    .Z(net824));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input825 (.I(itasegm[842]),
    .Z(net825));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input826 (.I(itasegm[843]),
    .Z(net826));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input827 (.I(itasegm[844]),
    .Z(net827));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input828 (.I(itasegm[845]),
    .Z(net828));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input829 (.I(itasegm[846]),
    .Z(net829));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input83 (.I(itasegm[174]),
    .Z(net83));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input830 (.I(itasegm[847]),
    .Z(net830));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input831 (.I(itasegm[848]),
    .Z(net831));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input832 (.I(itasegm[849]),
    .Z(net832));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input833 (.I(itasegm[84]),
    .Z(net833));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input834 (.I(itasegm[850]),
    .Z(net834));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input835 (.I(itasegm[851]),
    .Z(net835));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input836 (.I(itasegm[852]),
    .Z(net836));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input837 (.I(itasegm[853]),
    .Z(net837));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input838 (.I(itasegm[854]),
    .Z(net838));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input839 (.I(itasegm[855]),
    .Z(net839));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input84 (.I(itasegm[175]),
    .Z(net84));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input840 (.I(itasegm[856]),
    .Z(net840));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input841 (.I(itasegm[857]),
    .Z(net841));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input842 (.I(itasegm[858]),
    .Z(net842));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input843 (.I(itasegm[859]),
    .Z(net843));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input844 (.I(itasegm[85]),
    .Z(net844));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input845 (.I(itasegm[860]),
    .Z(net845));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input846 (.I(itasegm[861]),
    .Z(net846));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input847 (.I(itasegm[862]),
    .Z(net847));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input848 (.I(itasegm[863]),
    .Z(net848));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input849 (.I(itasegm[864]),
    .Z(net849));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input85 (.I(itasegm[176]),
    .Z(net85));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input850 (.I(itasegm[865]),
    .Z(net850));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input851 (.I(itasegm[866]),
    .Z(net851));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input852 (.I(itasegm[867]),
    .Z(net852));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input853 (.I(itasegm[868]),
    .Z(net853));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input854 (.I(itasegm[869]),
    .Z(net854));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input855 (.I(itasegm[86]),
    .Z(net855));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input856 (.I(itasegm[870]),
    .Z(net856));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input857 (.I(itasegm[871]),
    .Z(net857));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input858 (.I(itasegm[872]),
    .Z(net858));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input859 (.I(itasegm[873]),
    .Z(net859));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input86 (.I(itasegm[177]),
    .Z(net86));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input860 (.I(itasegm[874]),
    .Z(net860));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input861 (.I(itasegm[875]),
    .Z(net861));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input862 (.I(itasegm[876]),
    .Z(net862));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input863 (.I(itasegm[877]),
    .Z(net863));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input864 (.I(itasegm[878]),
    .Z(net864));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input865 (.I(itasegm[879]),
    .Z(net865));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input866 (.I(itasegm[87]),
    .Z(net866));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input867 (.I(itasegm[880]),
    .Z(net867));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input868 (.I(itasegm[881]),
    .Z(net868));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input869 (.I(itasegm[882]),
    .Z(net869));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input87 (.I(itasegm[178]),
    .Z(net87));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input870 (.I(itasegm[883]),
    .Z(net870));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input871 (.I(itasegm[884]),
    .Z(net871));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input872 (.I(itasegm[885]),
    .Z(net872));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input873 (.I(itasegm[886]),
    .Z(net873));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input874 (.I(itasegm[887]),
    .Z(net874));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input875 (.I(itasegm[888]),
    .Z(net875));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input876 (.I(itasegm[889]),
    .Z(net876));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input877 (.I(itasegm[88]),
    .Z(net877));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input878 (.I(itasegm[890]),
    .Z(net878));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input879 (.I(itasegm[891]),
    .Z(net879));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input88 (.I(itasegm[179]),
    .Z(net88));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input880 (.I(itasegm[892]),
    .Z(net880));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input881 (.I(itasegm[893]),
    .Z(net881));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input882 (.I(itasegm[894]),
    .Z(net882));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input883 (.I(itasegm[895]),
    .Z(net883));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input884 (.I(itasegm[89]),
    .Z(net884));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input885 (.I(itasegm[8]),
    .Z(net885));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input886 (.I(itasegm[90]),
    .Z(net886));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input887 (.I(itasegm[91]),
    .Z(net887));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input888 (.I(itasegm[92]),
    .Z(net888));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input889 (.I(itasegm[93]),
    .Z(net889));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input89 (.I(itasegm[17]),
    .Z(net89));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input890 (.I(itasegm[94]),
    .Z(net890));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input891 (.I(itasegm[95]),
    .Z(net891));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input892 (.I(itasegm[96]),
    .Z(net892));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input893 (.I(itasegm[97]),
    .Z(net893));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input894 (.I(itasegm[98]),
    .Z(net894));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input895 (.I(itasegm[99]),
    .Z(net895));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input896 (.I(itasegm[9]),
    .Z(net896));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input897 (.I(itasel[0]),
    .Z(net897));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input898 (.I(itasel[100]),
    .Z(net898));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input899 (.I(itasel[101]),
    .Z(net899));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input9 (.I(itasegm[107]),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input90 (.I(itasegm[180]),
    .Z(net90));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input900 (.I(itasel[102]),
    .Z(net900));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input901 (.I(itasel[103]),
    .Z(net901));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input902 (.I(itasel[104]),
    .Z(net902));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input903 (.I(itasel[105]),
    .Z(net903));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input904 (.I(itasel[106]),
    .Z(net904));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input905 (.I(itasel[107]),
    .Z(net905));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input906 (.I(itasel[108]),
    .Z(net906));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input907 (.I(itasel[109]),
    .Z(net907));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input908 (.I(itasel[10]),
    .Z(net908));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input909 (.I(itasel[110]),
    .Z(net909));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input91 (.I(itasegm[181]),
    .Z(net91));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input910 (.I(itasel[111]),
    .Z(net910));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input911 (.I(itasel[112]),
    .Z(net911));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input912 (.I(itasel[113]),
    .Z(net912));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input913 (.I(itasel[114]),
    .Z(net913));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input914 (.I(itasel[115]),
    .Z(net914));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input915 (.I(itasel[116]),
    .Z(net915));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input916 (.I(itasel[117]),
    .Z(net916));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input917 (.I(itasel[118]),
    .Z(net917));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input918 (.I(itasel[119]),
    .Z(net918));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input919 (.I(itasel[11]),
    .Z(net919));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input92 (.I(itasegm[182]),
    .Z(net92));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input920 (.I(itasel[120]),
    .Z(net920));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input921 (.I(itasel[121]),
    .Z(net921));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input922 (.I(itasel[122]),
    .Z(net922));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input923 (.I(itasel[123]),
    .Z(net923));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input924 (.I(itasel[124]),
    .Z(net924));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input925 (.I(itasel[125]),
    .Z(net925));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input926 (.I(itasel[126]),
    .Z(net926));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input927 (.I(itasel[127]),
    .Z(net927));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input928 (.I(itasel[128]),
    .Z(net928));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input929 (.I(itasel[129]),
    .Z(net929));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input93 (.I(itasegm[183]),
    .Z(net93));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input930 (.I(itasel[12]),
    .Z(net930));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input931 (.I(itasel[130]),
    .Z(net931));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input932 (.I(itasel[131]),
    .Z(net932));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input933 (.I(itasel[132]),
    .Z(net933));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input934 (.I(itasel[133]),
    .Z(net934));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input935 (.I(itasel[134]),
    .Z(net935));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input936 (.I(itasel[135]),
    .Z(net936));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input937 (.I(itasel[136]),
    .Z(net937));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input938 (.I(itasel[137]),
    .Z(net938));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input939 (.I(itasel[138]),
    .Z(net939));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input94 (.I(itasegm[184]),
    .Z(net94));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input940 (.I(itasel[139]),
    .Z(net940));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input941 (.I(itasel[13]),
    .Z(net941));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input942 (.I(itasel[140]),
    .Z(net942));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input943 (.I(itasel[141]),
    .Z(net943));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input944 (.I(itasel[142]),
    .Z(net944));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input945 (.I(itasel[143]),
    .Z(net945));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input946 (.I(itasel[144]),
    .Z(net946));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input947 (.I(itasel[145]),
    .Z(net947));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input948 (.I(itasel[146]),
    .Z(net948));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input949 (.I(itasel[147]),
    .Z(net949));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input95 (.I(itasegm[185]),
    .Z(net95));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input950 (.I(itasel[148]),
    .Z(net950));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input951 (.I(itasel[149]),
    .Z(net951));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input952 (.I(itasel[14]),
    .Z(net952));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input953 (.I(itasel[150]),
    .Z(net953));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input954 (.I(itasel[151]),
    .Z(net954));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input955 (.I(itasel[152]),
    .Z(net955));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input956 (.I(itasel[153]),
    .Z(net956));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input957 (.I(itasel[154]),
    .Z(net957));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input958 (.I(itasel[155]),
    .Z(net958));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input959 (.I(itasel[156]),
    .Z(net959));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input96 (.I(itasegm[186]),
    .Z(net96));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input960 (.I(itasel[157]),
    .Z(net960));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input961 (.I(itasel[158]),
    .Z(net961));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input962 (.I(itasel[159]),
    .Z(net962));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input963 (.I(itasel[15]),
    .Z(net963));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input964 (.I(itasel[160]),
    .Z(net964));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input965 (.I(itasel[161]),
    .Z(net965));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input966 (.I(itasel[162]),
    .Z(net966));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input967 (.I(itasel[163]),
    .Z(net967));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input968 (.I(itasel[164]),
    .Z(net968));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input969 (.I(itasel[165]),
    .Z(net969));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input97 (.I(itasegm[187]),
    .Z(net97));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input970 (.I(itasel[166]),
    .Z(net970));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input971 (.I(itasel[167]),
    .Z(net971));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input972 (.I(itasel[168]),
    .Z(net972));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input973 (.I(itasel[169]),
    .Z(net973));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input974 (.I(itasel[16]),
    .Z(net974));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input975 (.I(itasel[170]),
    .Z(net975));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input976 (.I(itasel[171]),
    .Z(net976));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input977 (.I(itasel[172]),
    .Z(net977));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input978 (.I(itasel[173]),
    .Z(net978));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input979 (.I(itasel[174]),
    .Z(net979));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input98 (.I(itasegm[188]),
    .Z(net98));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input980 (.I(itasel[175]),
    .Z(net980));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input981 (.I(itasel[176]),
    .Z(net981));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input982 (.I(itasel[177]),
    .Z(net982));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input983 (.I(itasel[178]),
    .Z(net983));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input984 (.I(itasel[179]),
    .Z(net984));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input985 (.I(itasel[17]),
    .Z(net985));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 input986 (.I(itasel[180]),
    .Z(net986));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 input987 (.I(itasel[181]),
    .Z(net987));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 input988 (.I(itasel[182]),
    .Z(net988));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 input989 (.I(itasel[183]),
    .Z(net989));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input99 (.I(itasegm[189]),
    .Z(net99));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 input990 (.I(itasel[184]),
    .Z(net990));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 input991 (.I(itasel[185]),
    .Z(net991));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input992 (.I(itasel[186]),
    .Z(net992));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input993 (.I(itasel[187]),
    .Z(net993));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input994 (.I(itasel[188]),
    .Z(net994));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input995 (.I(itasel[189]),
    .Z(net995));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input996 (.I(itasel[18]),
    .Z(net996));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 input997 (.I(itasel[190]),
    .Z(net997));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 input998 (.I(itasel[191]),
    .Z(net998));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input999 (.I(itasel[192]),
    .Z(net999));
 gf180mcu_fd_sc_mcu7t5v0__tiel ita_1829 (.ZN(net1829));
 gf180mcu_fd_sc_mcu7t5v0__tiel ita_1830 (.ZN(net1830));
 gf180mcu_fd_sc_mcu7t5v0__tiel ita_1831 (.ZN(net1831));
 gf180mcu_fd_sc_mcu7t5v0__tiel ita_1832 (.ZN(net1832));
 gf180mcu_fd_sc_mcu7t5v0__tiel ita_1833 (.ZN(net1833));
 gf180mcu_fd_sc_mcu7t5v0__tiel ita_1834 (.ZN(net1834));
 gf180mcu_fd_sc_mcu7t5v0__tiel ita_1835 (.ZN(net1835));
 gf180mcu_fd_sc_mcu7t5v0__tiel ita_1836 (.ZN(net1836));
 gf180mcu_fd_sc_mcu7t5v0__tiel ita_1837 (.ZN(net1837));
 gf180mcu_fd_sc_mcu7t5v0__tiel ita_1838 (.ZN(net1838));
 gf180mcu_fd_sc_mcu7t5v0__tiel ita_1839 (.ZN(net1839));
 gf180mcu_fd_sc_mcu7t5v0__tiel ita_1840 (.ZN(net1840));
 gf180mcu_fd_sc_mcu7t5v0__tiel ita_1841 (.ZN(net1841));
 gf180mcu_fd_sc_mcu7t5v0__tiel ita_1842 (.ZN(net1842));
 gf180mcu_fd_sc_mcu7t5v0__tiel ita_1843 (.ZN(net1843));
 gf180mcu_fd_sc_mcu7t5v0__tiel ita_1844 (.ZN(net1844));
 gf180mcu_fd_sc_mcu7t5v0__tiel ita_1845 (.ZN(net1845));
 gf180mcu_fd_sc_mcu7t5v0__tiel ita_1846 (.ZN(net1846));
 gf180mcu_fd_sc_mcu7t5v0__tiel ita_1847 (.ZN(net1847));
 gf180mcu_fd_sc_mcu7t5v0__tiel ita_1848 (.ZN(net1848));
 gf180mcu_fd_sc_mcu7t5v0__tiel ita_1849 (.ZN(net1849));
 gf180mcu_fd_sc_mcu7t5v0__tiel ita_1850 (.ZN(net1850));
 gf180mcu_fd_sc_mcu7t5v0__tiel ita_1851 (.ZN(net1851));
 gf180mcu_fd_sc_mcu7t5v0__tiel ita_1852 (.ZN(net1852));
 gf180mcu_fd_sc_mcu7t5v0__tiel ita_1853 (.ZN(net1853));
 gf180mcu_fd_sc_mcu7t5v0__tiel ita_1854 (.ZN(net1854));
 gf180mcu_fd_sc_mcu7t5v0__tieh ita_1855 (.Z(net1855));
 gf180mcu_fd_sc_mcu7t5v0__tieh ita_1856 (.Z(net1856));
 gf180mcu_fd_sc_mcu7t5v0__tieh ita_1857 (.Z(net1857));
 gf180mcu_fd_sc_mcu7t5v0__tieh ita_1858 (.Z(net1858));
 gf180mcu_fd_sc_mcu7t5v0__tieh ita_1859 (.Z(net1859));
 gf180mcu_fd_sc_mcu7t5v0__tieh ita_1860 (.Z(net1860));
 gf180mcu_fd_sc_mcu7t5v0__tieh ita_1861 (.Z(net1861));
 gf180mcu_fd_sc_mcu7t5v0__tieh ita_1862 (.Z(net1862));
 gf180mcu_fd_sc_mcu7t5v0__tieh ita_1863 (.Z(net1863));
 gf180mcu_fd_sc_mcu7t5v0__tieh ita_1864 (.Z(net1864));
 gf180mcu_fd_sc_mcu7t5v0__tieh ita_1865 (.Z(net1865));
 gf180mcu_fd_sc_mcu7t5v0__tieh ita_1866 (.Z(net1866));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output1671 (.I(net1671),
    .Z(segm[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output1672 (.I(net1672),
    .Z(segm[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output1673 (.I(net1673),
    .Z(segm[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output1674 (.I(net1674),
    .Z(segm[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output1675 (.I(net1675),
    .Z(segm[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output1676 (.I(net1676),
    .Z(segm[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output1677 (.I(net1677),
    .Z(segm[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output1678 (.I(net1678),
    .Z(segm[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output1679 (.I(net1679),
    .Z(segm[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output1680 (.I(net1680),
    .Z(segm[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output1681 (.I(net1681),
    .Z(segm[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output1682 (.I(net1682),
    .Z(segm[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output1683 (.I(net1683),
    .Z(segm[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output1684 (.I(net1684),
    .Z(segm[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output1685 (.I(net1685),
    .Z(sel[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output1686 (.I(net1686),
    .Z(sel[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output1687 (.I(net1687),
    .Z(sel[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output1688 (.I(net1688),
    .Z(sel[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output1689 (.I(net1689),
    .Z(sel[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output1690 (.I(net1690),
    .Z(sel[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output1691 (.I(net1691),
    .Z(sel[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output1692 (.I(net1692),
    .Z(sel[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output1693 (.I(net1693),
    .Z(sel[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output1694 (.I(net1694),
    .Z(sel[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output1695 (.I(net1695),
    .Z(sel[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output1696 (.I(net1696),
    .Z(sel[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire1697 (.I(_0818_),
    .Z(net1697));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire1698 (.I(_0756_),
    .Z(net1698));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire1699 (.I(_0691_),
    .Z(net1699));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire1700 (.I(_0597_),
    .Z(net1700));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 wire1701 (.I(_0498_),
    .Z(net1701));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire1702 (.I(_0436_),
    .Z(net1702));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire1703 (.I(_0372_),
    .Z(net1703));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire1704 (.I(_1302_),
    .Z(net1704));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 wire1705 (.I(_0834_),
    .Z(net1705));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire1706 (.I(net1707),
    .Z(net1706));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire1707 (.I(_0826_),
    .Z(net1707));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire1708 (.I(net1709),
    .Z(net1708));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 wire1709 (.I(_0822_),
    .Z(net1709));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire1710 (.I(_0808_),
    .Z(net1710));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 wire1711 (.I(_0773_),
    .Z(net1711));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire1712 (.I(net1713),
    .Z(net1712));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire1713 (.I(_0765_),
    .Z(net1713));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire1714 (.I(net1715),
    .Z(net1714));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 wire1715 (.I(_0760_),
    .Z(net1715));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire1716 (.I(_0745_),
    .Z(net1716));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 wire1717 (.I(_0707_),
    .Z(net1717));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire1718 (.I(net1719),
    .Z(net1718));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 wire1719 (.I(_0699_),
    .Z(net1719));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire1720 (.I(net1721),
    .Z(net1720));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 wire1721 (.I(_0695_),
    .Z(net1721));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire1722 (.I(_0681_),
    .Z(net1722));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 wire1723 (.I(_0630_),
    .Z(net1723));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire1724 (.I(net1725),
    .Z(net1724));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire1725 (.I(_0614_),
    .Z(net1725));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire1726 (.I(net1727),
    .Z(net1726));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 wire1727 (.I(_0606_),
    .Z(net1727));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire1728 (.I(_0574_),
    .Z(net1728));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 wire1729 (.I(_0514_),
    .Z(net1729));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire1730 (.I(net1731),
    .Z(net1730));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 wire1731 (.I(_0506_),
    .Z(net1731));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire1732 (.I(net1733),
    .Z(net1732));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 wire1733 (.I(_0502_),
    .Z(net1733));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire1734 (.I(_0488_),
    .Z(net1734));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 wire1735 (.I(_0453_),
    .Z(net1735));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire1736 (.I(net1737),
    .Z(net1736));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 wire1737 (.I(_0445_),
    .Z(net1737));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire1738 (.I(net1739),
    .Z(net1738));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 wire1739 (.I(_0440_),
    .Z(net1739));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire1740 (.I(_0425_),
    .Z(net1740));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 wire1741 (.I(_0388_),
    .Z(net1741));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire1742 (.I(net1743),
    .Z(net1742));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 wire1743 (.I(_0380_),
    .Z(net1743));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire1744 (.I(net1745),
    .Z(net1744));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire1745 (.I(_0376_),
    .Z(net1745));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire1746 (.I(_0362_),
    .Z(net1746));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 wire1747 (.I(_0276_),
    .Z(net1747));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire1748 (.I(net1749),
    .Z(net1748));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 wire1749 (.I(_0244_),
    .Z(net1749));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire1750 (.I(net1751),
    .Z(net1750));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 wire1751 (.I(_0225_),
    .Z(net1751));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire1752 (.I(_0144_),
    .Z(net1752));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire1753 (.I(_2174_),
    .Z(net1753));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 wire1754 (.I(_2166_),
    .Z(net1754));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 wire1755 (.I(_2162_),
    .Z(net1755));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire1756 (.I(_2113_),
    .Z(net1756));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 wire1757 (.I(_2105_),
    .Z(net1757));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 wire1758 (.I(_2100_),
    .Z(net1758));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire1759 (.I(_2048_),
    .Z(net1759));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 wire1760 (.I(_2040_),
    .Z(net1760));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire1761 (.I(_2036_),
    .Z(net1761));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire1762 (.I(_1971_),
    .Z(net1762));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 wire1763 (.I(_1955_),
    .Z(net1763));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire1764 (.I(_1947_),
    .Z(net1764));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 wire1765 (.I(_1856_),
    .Z(net1765));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire1766 (.I(_1848_),
    .Z(net1766));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire1767 (.I(_1844_),
    .Z(net1767));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 wire1768 (.I(_1795_),
    .Z(net1768));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire1769 (.I(_1787_),
    .Z(net1769));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire1770 (.I(_1782_),
    .Z(net1770));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 wire1771 (.I(_1730_),
    .Z(net1771));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire1772 (.I(_1722_),
    .Z(net1772));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire1773 (.I(_1718_),
    .Z(net1773));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 wire1774 (.I(_1694_),
    .Z(net1774));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 wire1775 (.I(_1690_),
    .Z(net1775));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 wire1776 (.I(_1653_),
    .Z(net1776));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire1777 (.I(_1637_),
    .Z(net1777));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire1778 (.I(_1629_),
    .Z(net1778));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire1779 (.I(net1780),
    .Z(net1779));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire1780 (.I(_1530_),
    .Z(net1780));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire1781 (.I(net1782),
    .Z(net1781));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire1782 (.I(_1526_),
    .Z(net1782));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 wire1783 (.I(_1502_),
    .Z(net1783));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 wire1784 (.I(_1498_),
    .Z(net1784));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire1785 (.I(net1786),
    .Z(net1785));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire1786 (.I(_1469_),
    .Z(net1786));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire1787 (.I(net1788),
    .Z(net1787));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire1788 (.I(_1464_),
    .Z(net1788));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 wire1789 (.I(_1438_),
    .Z(net1789));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 wire1790 (.I(_1434_),
    .Z(net1790));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire1791 (.I(net1792),
    .Z(net1791));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire1792 (.I(_1404_),
    .Z(net1792));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire1793 (.I(net1794),
    .Z(net1793));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire1794 (.I(_1400_),
    .Z(net1794));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire1795 (.I(net1796),
    .Z(net1795));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire1796 (.I(_1319_),
    .Z(net1796));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire1797 (.I(net1798),
    .Z(net1797));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire1798 (.I(_1311_),
    .Z(net1798));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire1799 (.I(net1800),
    .Z(net1799));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire1800 (.I(_1212_),
    .Z(net1800));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire1801 (.I(net1802),
    .Z(net1801));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire1802 (.I(_1208_),
    .Z(net1802));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire1803 (.I(net1804),
    .Z(net1803));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire1804 (.I(_1151_),
    .Z(net1804));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire1805 (.I(net1806),
    .Z(net1805));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire1806 (.I(_1145_),
    .Z(net1806));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire1807 (.I(net1808),
    .Z(net1807));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire1808 (.I(_1085_),
    .Z(net1808));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire1809 (.I(net1810),
    .Z(net1809));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire1810 (.I(_1081_),
    .Z(net1810));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire1811 (.I(net1812),
    .Z(net1811));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire1812 (.I(_0976_),
    .Z(net1812));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire1813 (.I(net1814),
    .Z(net1813));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire1814 (.I(_0964_),
    .Z(net1814));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 wire1815 (.I(_2296_),
    .Z(net1815));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire1816 (.I(_2288_),
    .Z(net1816));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire1817 (.I(_2284_),
    .Z(net1817));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire1818 (.I(_2270_),
    .Z(net1818));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 wire1819 (.I(_2235_),
    .Z(net1819));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire1820 (.I(_2227_),
    .Z(net1820));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire1821 (.I(_2223_),
    .Z(net1821));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 wire1822 (.I(_2209_),
    .Z(net1822));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 wire1823 (.I(_0801_),
    .Z(net1823));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 wire1824 (.I(_0738_),
    .Z(net1824));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 wire1825 (.I(_0674_),
    .Z(net1825));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 wire1826 (.I(_0560_),
    .Z(net1826));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 wire1827 (.I(_2263_),
    .Z(net1827));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 wire1828 (.I(_2202_),
    .Z(net1828));
 assign io_oeb[0] = net1855;
 assign io_oeb[10] = net1865;
 assign io_oeb[11] = net1866;
 assign io_oeb[12] = net1829;
 assign io_oeb[13] = net1830;
 assign io_oeb[14] = net1831;
 assign io_oeb[15] = net1832;
 assign io_oeb[16] = net1833;
 assign io_oeb[17] = net1834;
 assign io_oeb[18] = net1835;
 assign io_oeb[19] = net1836;
 assign io_oeb[1] = net1856;
 assign io_oeb[20] = net1837;
 assign io_oeb[21] = net1838;
 assign io_oeb[22] = net1839;
 assign io_oeb[23] = net1840;
 assign io_oeb[24] = net1841;
 assign io_oeb[25] = net1842;
 assign io_oeb[26] = net1843;
 assign io_oeb[27] = net1844;
 assign io_oeb[28] = net1845;
 assign io_oeb[29] = net1846;
 assign io_oeb[2] = net1857;
 assign io_oeb[30] = net1847;
 assign io_oeb[31] = net1848;
 assign io_oeb[32] = net1849;
 assign io_oeb[33] = net1850;
 assign io_oeb[34] = net1851;
 assign io_oeb[35] = net1852;
 assign io_oeb[36] = net1853;
 assign io_oeb[37] = net1854;
 assign io_oeb[3] = net1858;
 assign io_oeb[4] = net1859;
 assign io_oeb[5] = net1860;
 assign io_oeb[6] = net1861;
 assign io_oeb[7] = net1862;
 assign io_oeb[8] = net1863;
 assign io_oeb[9] = net1864;
endmodule

