magic
tech gf180mcuD
magscale 1 10
timestamp 1699645458
<< metal1 >>
rect 26898 38558 26910 38610
rect 26962 38607 26974 38610
rect 27458 38607 27470 38610
rect 26962 38561 27470 38607
rect 26962 38558 26974 38561
rect 27458 38558 27470 38561
rect 27522 38558 27534 38610
rect 1344 38442 40656 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 40656 38442
rect 1344 38356 40656 38390
rect 18622 38274 18674 38286
rect 18622 38210 18674 38222
rect 22430 38274 22482 38286
rect 22430 38210 22482 38222
rect 25566 38274 25618 38286
rect 25566 38210 25618 38222
rect 17826 37998 17838 38050
rect 17890 37998 17902 38050
rect 21522 37998 21534 38050
rect 21586 37998 21598 38050
rect 24546 37998 24558 38050
rect 24610 37998 24622 38050
rect 27470 37938 27522 37950
rect 27470 37874 27522 37886
rect 1344 37658 40656 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 40656 37658
rect 1344 37572 40656 37606
rect 18398 37490 18450 37502
rect 18398 37426 18450 37438
rect 20078 37490 20130 37502
rect 20078 37426 20130 37438
rect 26238 37490 26290 37502
rect 26238 37426 26290 37438
rect 19394 37214 19406 37266
rect 19458 37214 19470 37266
rect 25218 37214 25230 37266
rect 25282 37214 25294 37266
rect 1344 36874 40656 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 40656 36874
rect 1344 36788 40656 36822
rect 1710 36370 1762 36382
rect 1710 36306 1762 36318
rect 1344 36090 40656 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 40656 36090
rect 1344 36004 40656 36038
rect 1344 35306 40656 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 40656 35306
rect 1344 35220 40656 35254
rect 1344 34522 40656 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 40656 34522
rect 1344 34436 40656 34470
rect 1344 33738 40656 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 40656 33738
rect 1344 33652 40656 33686
rect 1344 32954 40656 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 40656 32954
rect 1344 32868 40656 32902
rect 1344 32170 40656 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 40656 32170
rect 1344 32084 40656 32118
rect 1344 31386 40656 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 40656 31386
rect 1344 31300 40656 31334
rect 1344 30602 40656 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 40656 30602
rect 1344 30516 40656 30550
rect 1344 29818 40656 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 40656 29818
rect 1344 29732 40656 29766
rect 1344 29034 40656 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 40656 29034
rect 1344 28948 40656 28982
rect 21982 28754 22034 28766
rect 21982 28690 22034 28702
rect 21870 28642 21922 28654
rect 21870 28578 21922 28590
rect 1344 28250 40656 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 40656 28250
rect 1344 28164 40656 28198
rect 19742 27970 19794 27982
rect 20850 27918 20862 27970
rect 20914 27918 20926 27970
rect 19742 27906 19794 27918
rect 23550 27858 23602 27870
rect 19506 27806 19518 27858
rect 19570 27806 19582 27858
rect 20178 27806 20190 27858
rect 20242 27806 20254 27858
rect 23550 27794 23602 27806
rect 22978 27694 22990 27746
rect 23042 27694 23054 27746
rect 1344 27466 40656 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 40656 27466
rect 1344 27380 40656 27414
rect 21646 27298 21698 27310
rect 21646 27234 21698 27246
rect 19854 27186 19906 27198
rect 19394 27134 19406 27186
rect 19458 27134 19470 27186
rect 19854 27122 19906 27134
rect 20302 27186 20354 27198
rect 20302 27122 20354 27134
rect 21870 27074 21922 27086
rect 16482 27022 16494 27074
rect 16546 27022 16558 27074
rect 21870 27010 21922 27022
rect 16158 26962 16210 26974
rect 20190 26962 20242 26974
rect 17266 26910 17278 26962
rect 17330 26910 17342 26962
rect 16158 26898 16210 26910
rect 20190 26898 20242 26910
rect 20526 26962 20578 26974
rect 20526 26898 20578 26910
rect 20750 26962 20802 26974
rect 21298 26910 21310 26962
rect 21362 26910 21374 26962
rect 20750 26898 20802 26910
rect 16046 26850 16098 26862
rect 16046 26786 16098 26798
rect 19742 26850 19794 26862
rect 19742 26786 19794 26798
rect 1344 26682 40656 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 40656 26682
rect 1344 26596 40656 26630
rect 17838 26514 17890 26526
rect 17838 26450 17890 26462
rect 17950 26514 18002 26526
rect 17950 26450 18002 26462
rect 17726 26290 17778 26302
rect 4274 26238 4286 26290
rect 4338 26238 4350 26290
rect 15138 26238 15150 26290
rect 15202 26238 15214 26290
rect 17726 26226 17778 26238
rect 18062 26290 18114 26302
rect 18274 26238 18286 26290
rect 18338 26238 18350 26290
rect 21858 26238 21870 26290
rect 21922 26238 21934 26290
rect 18062 26226 18114 26238
rect 15598 26178 15650 26190
rect 12226 26126 12238 26178
rect 12290 26126 12302 26178
rect 14354 26126 14366 26178
rect 14418 26126 14430 26178
rect 15598 26114 15650 26126
rect 19630 26178 19682 26190
rect 25342 26178 25394 26190
rect 22530 26126 22542 26178
rect 22594 26126 22606 26178
rect 24658 26126 24670 26178
rect 24722 26126 24734 26178
rect 19630 26114 19682 26126
rect 25342 26114 25394 26126
rect 1934 26066 1986 26078
rect 1934 26002 1986 26014
rect 1344 25898 40656 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 40656 25898
rect 1344 25812 40656 25846
rect 14366 25730 14418 25742
rect 14366 25666 14418 25678
rect 18510 25618 18562 25630
rect 15810 25566 15822 25618
rect 15874 25566 15886 25618
rect 17938 25566 17950 25618
rect 18002 25566 18014 25618
rect 18510 25554 18562 25566
rect 18622 25506 18674 25518
rect 15138 25454 15150 25506
rect 15202 25454 15214 25506
rect 18622 25442 18674 25454
rect 18846 25506 18898 25518
rect 18846 25442 18898 25454
rect 18958 25506 19010 25518
rect 18958 25442 19010 25454
rect 19406 25506 19458 25518
rect 19406 25442 19458 25454
rect 14702 25394 14754 25406
rect 14702 25330 14754 25342
rect 18398 25394 18450 25406
rect 18398 25330 18450 25342
rect 14478 25282 14530 25294
rect 14478 25218 14530 25230
rect 1344 25114 40656 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 40656 25114
rect 1344 25028 40656 25062
rect 15486 24946 15538 24958
rect 15486 24882 15538 24894
rect 15598 24946 15650 24958
rect 15598 24882 15650 24894
rect 23662 24946 23714 24958
rect 23662 24882 23714 24894
rect 15262 24834 15314 24846
rect 15262 24770 15314 24782
rect 26798 24834 26850 24846
rect 26798 24770 26850 24782
rect 27694 24834 27746 24846
rect 27694 24770 27746 24782
rect 15710 24722 15762 24734
rect 22654 24722 22706 24734
rect 4274 24670 4286 24722
rect 4338 24670 4350 24722
rect 14914 24670 14926 24722
rect 14978 24670 14990 24722
rect 15922 24670 15934 24722
rect 15986 24670 15998 24722
rect 19394 24670 19406 24722
rect 19458 24670 19470 24722
rect 15710 24658 15762 24670
rect 22654 24658 22706 24670
rect 23102 24722 23154 24734
rect 26462 24722 26514 24734
rect 27358 24722 27410 24734
rect 23426 24670 23438 24722
rect 23490 24670 23502 24722
rect 27010 24670 27022 24722
rect 27074 24670 27086 24722
rect 37874 24670 37886 24722
rect 37938 24670 37950 24722
rect 23102 24658 23154 24670
rect 26462 24658 26514 24670
rect 27358 24658 27410 24670
rect 16382 24610 16434 24622
rect 12002 24558 12014 24610
rect 12066 24558 12078 24610
rect 14130 24558 14142 24610
rect 14194 24558 14206 24610
rect 16382 24546 16434 24558
rect 18174 24610 18226 24622
rect 20066 24558 20078 24610
rect 20130 24558 20142 24610
rect 22194 24558 22206 24610
rect 22258 24558 22270 24610
rect 23538 24558 23550 24610
rect 23602 24558 23614 24610
rect 18174 24546 18226 24558
rect 1934 24498 1986 24510
rect 1934 24434 1986 24446
rect 27134 24498 27186 24510
rect 27134 24434 27186 24446
rect 40014 24498 40066 24510
rect 40014 24434 40066 24446
rect 1344 24330 40656 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 40656 24330
rect 1344 24244 40656 24278
rect 28030 24162 28082 24174
rect 28030 24098 28082 24110
rect 1934 24050 1986 24062
rect 19854 24050 19906 24062
rect 14802 23998 14814 24050
rect 14866 23998 14878 24050
rect 1934 23986 1986 23998
rect 19854 23986 19906 23998
rect 21422 24050 21474 24062
rect 21422 23986 21474 23998
rect 22990 24050 23042 24062
rect 27134 24050 27186 24062
rect 26674 23998 26686 24050
rect 26738 23998 26750 24050
rect 22990 23986 23042 23998
rect 27134 23986 27186 23998
rect 40014 24050 40066 24062
rect 40014 23986 40066 23998
rect 14142 23938 14194 23950
rect 19966 23938 20018 23950
rect 4274 23886 4286 23938
rect 4338 23886 4350 23938
rect 14914 23886 14926 23938
rect 14978 23886 14990 23938
rect 14142 23874 14194 23886
rect 19966 23874 20018 23886
rect 20190 23938 20242 23950
rect 20402 23886 20414 23938
rect 20466 23886 20478 23938
rect 21522 23886 21534 23938
rect 21586 23886 21598 23938
rect 22642 23886 22654 23938
rect 22706 23886 22718 23938
rect 23762 23886 23774 23938
rect 23826 23886 23838 23938
rect 37650 23886 37662 23938
rect 37714 23886 37726 23938
rect 20190 23874 20242 23886
rect 14366 23826 14418 23838
rect 14366 23762 14418 23774
rect 14478 23826 14530 23838
rect 14478 23762 14530 23774
rect 15262 23826 15314 23838
rect 15262 23762 15314 23774
rect 19742 23826 19794 23838
rect 19742 23762 19794 23774
rect 20638 23826 20690 23838
rect 20638 23762 20690 23774
rect 21310 23826 21362 23838
rect 21310 23762 21362 23774
rect 21758 23826 21810 23838
rect 21758 23762 21810 23774
rect 22206 23826 22258 23838
rect 23326 23826 23378 23838
rect 23202 23774 23214 23826
rect 23266 23774 23278 23826
rect 22206 23762 22258 23774
rect 23326 23762 23378 23774
rect 23438 23826 23490 23838
rect 27022 23826 27074 23838
rect 24546 23774 24558 23826
rect 24610 23774 24622 23826
rect 23438 23762 23490 23774
rect 27022 23762 27074 23774
rect 27358 23826 27410 23838
rect 27358 23762 27410 23774
rect 27582 23826 27634 23838
rect 27582 23762 27634 23774
rect 27918 23826 27970 23838
rect 27918 23762 27970 23774
rect 28030 23826 28082 23838
rect 28030 23762 28082 23774
rect 15374 23714 15426 23726
rect 15374 23650 15426 23662
rect 15598 23714 15650 23726
rect 15598 23650 15650 23662
rect 18062 23714 18114 23726
rect 19070 23714 19122 23726
rect 18386 23662 18398 23714
rect 18450 23662 18462 23714
rect 18722 23662 18734 23714
rect 18786 23662 18798 23714
rect 18062 23650 18114 23662
rect 19070 23650 19122 23662
rect 22318 23714 22370 23726
rect 22318 23650 22370 23662
rect 1344 23546 40656 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 40656 23546
rect 1344 23460 40656 23494
rect 17726 23378 17778 23390
rect 12226 23326 12238 23378
rect 12290 23326 12302 23378
rect 17726 23314 17778 23326
rect 18398 23378 18450 23390
rect 18398 23314 18450 23326
rect 21982 23378 22034 23390
rect 21982 23314 22034 23326
rect 22094 23378 22146 23390
rect 25454 23378 25506 23390
rect 22866 23326 22878 23378
rect 22930 23326 22942 23378
rect 22094 23314 22146 23326
rect 25454 23314 25506 23326
rect 26350 23378 26402 23390
rect 26350 23314 26402 23326
rect 15374 23266 15426 23278
rect 23550 23266 23602 23278
rect 18610 23214 18622 23266
rect 18674 23214 18686 23266
rect 20626 23214 20638 23266
rect 20690 23214 20702 23266
rect 15374 23202 15426 23214
rect 23550 23202 23602 23214
rect 24334 23266 24386 23278
rect 24334 23202 24386 23214
rect 26462 23266 26514 23278
rect 27570 23214 27582 23266
rect 27634 23214 27646 23266
rect 26462 23202 26514 23214
rect 15262 23154 15314 23166
rect 4274 23102 4286 23154
rect 4338 23102 4350 23154
rect 12450 23102 12462 23154
rect 12514 23102 12526 23154
rect 15262 23090 15314 23102
rect 15598 23154 15650 23166
rect 15598 23090 15650 23102
rect 17614 23154 17666 23166
rect 17614 23090 17666 23102
rect 17838 23154 17890 23166
rect 17838 23090 17890 23102
rect 18286 23154 18338 23166
rect 20862 23154 20914 23166
rect 18946 23102 18958 23154
rect 19010 23102 19022 23154
rect 19394 23102 19406 23154
rect 19458 23102 19470 23154
rect 19842 23102 19854 23154
rect 19906 23102 19918 23154
rect 18286 23090 18338 23102
rect 20862 23090 20914 23102
rect 22206 23154 22258 23166
rect 22206 23090 22258 23102
rect 22654 23154 22706 23166
rect 22654 23090 22706 23102
rect 22878 23154 22930 23166
rect 22878 23090 22930 23102
rect 23102 23154 23154 23166
rect 23102 23090 23154 23102
rect 23326 23154 23378 23166
rect 23326 23090 23378 23102
rect 23774 23154 23826 23166
rect 24098 23102 24110 23154
rect 24162 23102 24174 23154
rect 26114 23102 26126 23154
rect 26178 23102 26190 23154
rect 26786 23102 26798 23154
rect 26850 23102 26862 23154
rect 37650 23102 37662 23154
rect 37714 23102 37726 23154
rect 23774 23090 23826 23102
rect 13022 23042 13074 23054
rect 13022 22978 13074 22990
rect 25230 23042 25282 23054
rect 25442 22990 25454 23042
rect 25506 22990 25518 23042
rect 29698 22990 29710 23042
rect 29762 22990 29774 23042
rect 25230 22978 25282 22990
rect 1934 22930 1986 22942
rect 1934 22866 1986 22878
rect 24446 22930 24498 22942
rect 24446 22866 24498 22878
rect 40014 22930 40066 22942
rect 40014 22866 40066 22878
rect 1344 22762 40656 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 40656 22762
rect 1344 22676 40656 22710
rect 17278 22594 17330 22606
rect 17278 22530 17330 22542
rect 19630 22594 19682 22606
rect 19630 22530 19682 22542
rect 20414 22594 20466 22606
rect 20414 22530 20466 22542
rect 1934 22482 1986 22494
rect 29262 22482 29314 22494
rect 9874 22430 9886 22482
rect 9938 22430 9950 22482
rect 21858 22430 21870 22482
rect 21922 22430 21934 22482
rect 28578 22430 28590 22482
rect 28642 22430 28654 22482
rect 1934 22418 1986 22430
rect 29262 22418 29314 22430
rect 15150 22370 15202 22382
rect 15822 22370 15874 22382
rect 20078 22370 20130 22382
rect 23438 22370 23490 22382
rect 4274 22318 4286 22370
rect 4338 22318 4350 22370
rect 12786 22318 12798 22370
rect 12850 22318 12862 22370
rect 13682 22318 13694 22370
rect 13746 22318 13758 22370
rect 14466 22318 14478 22370
rect 14530 22318 14542 22370
rect 15586 22318 15598 22370
rect 15650 22318 15662 22370
rect 17826 22318 17838 22370
rect 17890 22318 17902 22370
rect 19058 22318 19070 22370
rect 19122 22318 19134 22370
rect 19282 22318 19294 22370
rect 19346 22318 19358 22370
rect 21298 22318 21310 22370
rect 21362 22318 21374 22370
rect 25778 22318 25790 22370
rect 25842 22318 25854 22370
rect 15150 22306 15202 22318
rect 15822 22306 15874 22318
rect 20078 22306 20130 22318
rect 23438 22306 23490 22318
rect 14926 22258 14978 22270
rect 12002 22206 12014 22258
rect 12066 22206 12078 22258
rect 13458 22206 13470 22258
rect 13522 22206 13534 22258
rect 14926 22194 14978 22206
rect 15038 22258 15090 22270
rect 15038 22194 15090 22206
rect 15262 22258 15314 22270
rect 15262 22194 15314 22206
rect 15934 22258 15986 22270
rect 15934 22194 15986 22206
rect 17166 22258 17218 22270
rect 17166 22194 17218 22206
rect 17278 22258 17330 22270
rect 19518 22258 19570 22270
rect 18722 22206 18734 22258
rect 18786 22206 18798 22258
rect 17278 22194 17330 22206
rect 19518 22194 19570 22206
rect 19854 22258 19906 22270
rect 21410 22206 21422 22258
rect 21474 22206 21486 22258
rect 25106 22206 25118 22258
rect 25170 22206 25182 22258
rect 26450 22206 26462 22258
rect 26514 22206 26526 22258
rect 19854 22194 19906 22206
rect 16046 22146 16098 22158
rect 16046 22082 16098 22094
rect 16158 22146 16210 22158
rect 16158 22082 16210 22094
rect 16830 22146 16882 22158
rect 18398 22146 18450 22158
rect 18050 22094 18062 22146
rect 18114 22094 18126 22146
rect 16830 22082 16882 22094
rect 18398 22082 18450 22094
rect 1344 21978 40656 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 40656 21978
rect 1344 21892 40656 21926
rect 15038 21810 15090 21822
rect 15038 21746 15090 21758
rect 17950 21810 18002 21822
rect 17950 21746 18002 21758
rect 25342 21810 25394 21822
rect 25342 21746 25394 21758
rect 25566 21810 25618 21822
rect 25566 21746 25618 21758
rect 26462 21810 26514 21822
rect 26462 21746 26514 21758
rect 26910 21810 26962 21822
rect 26910 21746 26962 21758
rect 27358 21810 27410 21822
rect 27358 21746 27410 21758
rect 14142 21698 14194 21710
rect 14142 21634 14194 21646
rect 14478 21698 14530 21710
rect 14478 21634 14530 21646
rect 14702 21698 14754 21710
rect 14702 21634 14754 21646
rect 15822 21698 15874 21710
rect 15822 21634 15874 21646
rect 16270 21698 16322 21710
rect 16270 21634 16322 21646
rect 25230 21698 25282 21710
rect 25230 21634 25282 21646
rect 18958 21586 19010 21598
rect 26238 21586 26290 21598
rect 4274 21534 4286 21586
rect 4338 21534 4350 21586
rect 13458 21534 13470 21586
rect 13522 21534 13534 21586
rect 15250 21534 15262 21586
rect 15314 21534 15326 21586
rect 15586 21534 15598 21586
rect 15650 21534 15662 21586
rect 16482 21534 16494 21586
rect 16546 21534 16558 21586
rect 17714 21534 17726 21586
rect 17778 21534 17790 21586
rect 19282 21534 19294 21586
rect 19346 21534 19358 21586
rect 26002 21534 26014 21586
rect 26066 21534 26078 21586
rect 18958 21522 19010 21534
rect 26238 21522 26290 21534
rect 26574 21586 26626 21598
rect 26574 21522 26626 21534
rect 27022 21586 27074 21598
rect 27022 21522 27074 21534
rect 27134 21586 27186 21598
rect 27134 21522 27186 21534
rect 1934 21474 1986 21486
rect 14254 21474 14306 21486
rect 10658 21422 10670 21474
rect 10722 21422 10734 21474
rect 12786 21422 12798 21474
rect 12850 21422 12862 21474
rect 18498 21422 18510 21474
rect 18562 21422 18574 21474
rect 22866 21422 22878 21474
rect 22930 21422 22942 21474
rect 1934 21410 1986 21422
rect 14254 21410 14306 21422
rect 16158 21362 16210 21374
rect 15250 21310 15262 21362
rect 15314 21310 15326 21362
rect 16158 21298 16210 21310
rect 18062 21362 18114 21374
rect 26002 21310 26014 21362
rect 26066 21310 26078 21362
rect 18062 21298 18114 21310
rect 1344 21194 40656 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 40656 21194
rect 1344 21108 40656 21142
rect 22206 21026 22258 21038
rect 22206 20962 22258 20974
rect 40014 20914 40066 20926
rect 26786 20862 26798 20914
rect 26850 20862 26862 20914
rect 40014 20850 40066 20862
rect 13918 20802 13970 20814
rect 13918 20738 13970 20750
rect 14478 20802 14530 20814
rect 15026 20750 15038 20802
rect 15090 20750 15102 20802
rect 20066 20750 20078 20802
rect 20130 20750 20142 20802
rect 21858 20750 21870 20802
rect 21922 20750 21934 20802
rect 22866 20750 22878 20802
rect 22930 20750 22942 20802
rect 37650 20750 37662 20802
rect 37714 20750 37726 20802
rect 14478 20738 14530 20750
rect 21646 20690 21698 20702
rect 14802 20638 14814 20690
rect 14866 20638 14878 20690
rect 17826 20638 17838 20690
rect 17890 20638 17902 20690
rect 21646 20626 21698 20638
rect 22094 20690 22146 20702
rect 22094 20626 22146 20638
rect 13582 20578 13634 20590
rect 13582 20514 13634 20526
rect 13806 20578 13858 20590
rect 13806 20514 13858 20526
rect 14142 20578 14194 20590
rect 14142 20514 14194 20526
rect 14366 20578 14418 20590
rect 14366 20514 14418 20526
rect 1344 20410 40656 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 40656 20410
rect 1344 20324 40656 20358
rect 26350 20242 26402 20254
rect 20178 20190 20190 20242
rect 20242 20190 20254 20242
rect 23538 20190 23550 20242
rect 23602 20190 23614 20242
rect 26350 20178 26402 20190
rect 15822 20130 15874 20142
rect 22430 20130 22482 20142
rect 17938 20078 17950 20130
rect 18002 20078 18014 20130
rect 18722 20078 18734 20130
rect 18786 20078 18798 20130
rect 19842 20078 19854 20130
rect 19906 20078 19918 20130
rect 20514 20078 20526 20130
rect 20578 20078 20590 20130
rect 24210 20078 24222 20130
rect 24274 20078 24286 20130
rect 25554 20078 25566 20130
rect 25618 20078 25630 20130
rect 15822 20066 15874 20078
rect 22430 20066 22482 20078
rect 16382 20018 16434 20030
rect 16034 19966 16046 20018
rect 16098 19966 16110 20018
rect 16382 19954 16434 19966
rect 18286 20018 18338 20030
rect 21534 20018 21586 20030
rect 18610 19966 18622 20018
rect 18674 19966 18686 20018
rect 19618 19966 19630 20018
rect 19682 19966 19694 20018
rect 18286 19954 18338 19966
rect 21534 19954 21586 19966
rect 22094 20018 22146 20030
rect 22990 20018 23042 20030
rect 22642 19966 22654 20018
rect 22706 19966 22718 20018
rect 22094 19954 22146 19966
rect 22990 19954 23042 19966
rect 23214 20018 23266 20030
rect 23214 19954 23266 19966
rect 23886 20018 23938 20030
rect 25778 19966 25790 20018
rect 25842 19966 25854 20018
rect 26786 19966 26798 20018
rect 26850 19966 26862 20018
rect 23886 19954 23938 19966
rect 13806 19906 13858 19918
rect 19282 19854 19294 19906
rect 19346 19854 19358 19906
rect 27458 19854 27470 19906
rect 27522 19854 27534 19906
rect 29586 19854 29598 19906
rect 29650 19854 29662 19906
rect 13806 19842 13858 19854
rect 15710 19794 15762 19806
rect 15710 19730 15762 19742
rect 22766 19794 22818 19806
rect 22766 19730 22818 19742
rect 1344 19626 40656 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 40656 19626
rect 1344 19540 40656 19574
rect 18734 19458 18786 19470
rect 18734 19394 18786 19406
rect 23550 19458 23602 19470
rect 23550 19394 23602 19406
rect 19070 19346 19122 19358
rect 21310 19346 21362 19358
rect 19506 19294 19518 19346
rect 19570 19294 19582 19346
rect 19070 19282 19122 19294
rect 21310 19282 21362 19294
rect 23102 19346 23154 19358
rect 23102 19282 23154 19294
rect 26798 19346 26850 19358
rect 26798 19282 26850 19294
rect 14030 19234 14082 19246
rect 14030 19170 14082 19182
rect 14702 19234 14754 19246
rect 14702 19170 14754 19182
rect 15150 19234 15202 19246
rect 15150 19170 15202 19182
rect 17614 19234 17666 19246
rect 17614 19170 17666 19182
rect 18622 19234 18674 19246
rect 18622 19170 18674 19182
rect 19406 19234 19458 19246
rect 22542 19234 22594 19246
rect 25678 19234 25730 19246
rect 21746 19182 21758 19234
rect 21810 19182 21822 19234
rect 22866 19182 22878 19234
rect 22930 19182 22942 19234
rect 19406 19170 19458 19182
rect 22542 19170 22594 19182
rect 25678 19170 25730 19182
rect 26574 19234 26626 19246
rect 26574 19170 26626 19182
rect 27022 19234 27074 19246
rect 27022 19170 27074 19182
rect 27134 19234 27186 19246
rect 27134 19170 27186 19182
rect 27806 19234 27858 19246
rect 27806 19170 27858 19182
rect 23214 19122 23266 19134
rect 16594 19070 16606 19122
rect 16658 19070 16670 19122
rect 17266 19070 17278 19122
rect 17330 19070 17342 19122
rect 22194 19070 22206 19122
rect 22258 19070 22270 19122
rect 23214 19058 23266 19070
rect 23662 19122 23714 19134
rect 23662 19058 23714 19070
rect 25342 19122 25394 19134
rect 25342 19058 25394 19070
rect 27582 19122 27634 19134
rect 27582 19058 27634 19070
rect 28142 19122 28194 19134
rect 28142 19058 28194 19070
rect 14478 19010 14530 19022
rect 14478 18946 14530 18958
rect 14590 19010 14642 19022
rect 14590 18946 14642 18958
rect 16942 19010 16994 19022
rect 16942 18946 16994 18958
rect 25454 19010 25506 19022
rect 25454 18946 25506 18958
rect 25902 19010 25954 19022
rect 27918 19010 27970 19022
rect 26226 18958 26238 19010
rect 26290 18958 26302 19010
rect 25902 18946 25954 18958
rect 27918 18946 27970 18958
rect 1344 18842 40656 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 40656 18842
rect 1344 18756 40656 18790
rect 15486 18674 15538 18686
rect 15486 18610 15538 18622
rect 17950 18674 18002 18686
rect 23326 18674 23378 18686
rect 21410 18622 21422 18674
rect 21474 18622 21486 18674
rect 17950 18610 18002 18622
rect 23326 18610 23378 18622
rect 25454 18674 25506 18686
rect 25454 18610 25506 18622
rect 26238 18674 26290 18686
rect 26238 18610 26290 18622
rect 14590 18562 14642 18574
rect 25230 18562 25282 18574
rect 16146 18510 16158 18562
rect 16210 18510 16222 18562
rect 20850 18510 20862 18562
rect 20914 18510 20926 18562
rect 27346 18510 27358 18562
rect 27410 18510 27422 18562
rect 14590 18498 14642 18510
rect 25230 18498 25282 18510
rect 14926 18450 14978 18462
rect 4274 18398 4286 18450
rect 4338 18398 4350 18450
rect 11442 18398 11454 18450
rect 11506 18398 11518 18450
rect 12114 18398 12126 18450
rect 12178 18398 12190 18450
rect 14926 18386 14978 18398
rect 15150 18450 15202 18462
rect 16494 18450 16546 18462
rect 18286 18450 18338 18462
rect 15698 18398 15710 18450
rect 15762 18398 15774 18450
rect 17714 18398 17726 18450
rect 17778 18398 17790 18450
rect 15150 18386 15202 18398
rect 16494 18386 16546 18398
rect 18286 18386 18338 18398
rect 18510 18450 18562 18462
rect 18510 18386 18562 18398
rect 19742 18450 19794 18462
rect 21982 18450 22034 18462
rect 20402 18398 20414 18450
rect 20466 18398 20478 18450
rect 21410 18398 21422 18450
rect 21474 18398 21486 18450
rect 19742 18386 19794 18398
rect 21982 18386 22034 18398
rect 22094 18450 22146 18462
rect 22094 18386 22146 18398
rect 22430 18450 22482 18462
rect 24670 18450 24722 18462
rect 23986 18398 23998 18450
rect 24050 18398 24062 18450
rect 22430 18386 22482 18398
rect 24670 18386 24722 18398
rect 25790 18450 25842 18462
rect 26562 18398 26574 18450
rect 26626 18398 26638 18450
rect 37650 18398 37662 18450
rect 37714 18398 37726 18450
rect 25790 18386 25842 18398
rect 14702 18338 14754 18350
rect 14242 18286 14254 18338
rect 14306 18286 14318 18338
rect 19394 18286 19406 18338
rect 19458 18286 19470 18338
rect 23762 18286 23774 18338
rect 23826 18286 23838 18338
rect 29474 18286 29486 18338
rect 29538 18286 29550 18338
rect 14702 18274 14754 18286
rect 1934 18226 1986 18238
rect 22654 18226 22706 18238
rect 18834 18174 18846 18226
rect 18898 18174 18910 18226
rect 19954 18174 19966 18226
rect 20018 18174 20030 18226
rect 1934 18162 1986 18174
rect 22654 18162 22706 18174
rect 22878 18226 22930 18238
rect 22878 18162 22930 18174
rect 25566 18226 25618 18238
rect 25566 18162 25618 18174
rect 40014 18226 40066 18238
rect 40014 18162 40066 18174
rect 1344 18058 40656 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 40656 18058
rect 1344 17972 40656 18006
rect 22206 17778 22258 17790
rect 15250 17726 15262 17778
rect 15314 17726 15326 17778
rect 17378 17726 17390 17778
rect 17442 17726 17454 17778
rect 20402 17726 20414 17778
rect 20466 17726 20478 17778
rect 22206 17714 22258 17726
rect 18734 17666 18786 17678
rect 27918 17666 27970 17678
rect 14466 17614 14478 17666
rect 14530 17614 14542 17666
rect 20626 17614 20638 17666
rect 20690 17614 20702 17666
rect 21746 17614 21758 17666
rect 21810 17614 21822 17666
rect 23202 17614 23214 17666
rect 23266 17614 23278 17666
rect 23986 17614 23998 17666
rect 24050 17614 24062 17666
rect 18734 17602 18786 17614
rect 27918 17602 27970 17614
rect 27582 17554 27634 17566
rect 19730 17502 19742 17554
rect 19794 17502 19806 17554
rect 23426 17502 23438 17554
rect 23490 17502 23502 17554
rect 27582 17490 27634 17502
rect 27694 17554 27746 17566
rect 27694 17490 27746 17502
rect 17838 17442 17890 17454
rect 20078 17442 20130 17454
rect 19058 17390 19070 17442
rect 19122 17390 19134 17442
rect 23762 17390 23774 17442
rect 23826 17390 23838 17442
rect 17838 17378 17890 17390
rect 20078 17378 20130 17390
rect 1344 17274 40656 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 40656 17274
rect 1344 17188 40656 17222
rect 14478 17106 14530 17118
rect 21086 17106 21138 17118
rect 27358 17106 27410 17118
rect 18722 17054 18734 17106
rect 18786 17054 18798 17106
rect 21410 17054 21422 17106
rect 21474 17054 21486 17106
rect 14478 17042 14530 17054
rect 21086 17042 21138 17054
rect 27358 17042 27410 17054
rect 27246 16994 27298 17006
rect 13234 16942 13246 16994
rect 13298 16942 13310 16994
rect 27246 16930 27298 16942
rect 19070 16882 19122 16894
rect 14018 16830 14030 16882
rect 14082 16830 14094 16882
rect 19070 16818 19122 16830
rect 27134 16882 27186 16894
rect 27134 16818 27186 16830
rect 27694 16882 27746 16894
rect 37874 16830 37886 16882
rect 37938 16830 37950 16882
rect 27694 16818 27746 16830
rect 11106 16718 11118 16770
rect 11170 16718 11182 16770
rect 39890 16718 39902 16770
rect 39954 16718 39966 16770
rect 1344 16490 40656 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 40656 16490
rect 1344 16404 40656 16438
rect 27694 16322 27746 16334
rect 27694 16258 27746 16270
rect 19966 16210 20018 16222
rect 19966 16146 20018 16158
rect 40014 16210 40066 16222
rect 40014 16146 40066 16158
rect 18510 16098 18562 16110
rect 18510 16034 18562 16046
rect 18734 16098 18786 16110
rect 18734 16034 18786 16046
rect 19070 16098 19122 16110
rect 19070 16034 19122 16046
rect 19294 16098 19346 16110
rect 19294 16034 19346 16046
rect 19518 16098 19570 16110
rect 19518 16034 19570 16046
rect 20190 16098 20242 16110
rect 20190 16034 20242 16046
rect 24110 16098 24162 16110
rect 24110 16034 24162 16046
rect 26126 16098 26178 16110
rect 26126 16034 26178 16046
rect 26574 16098 26626 16110
rect 26574 16034 26626 16046
rect 27022 16098 27074 16110
rect 27022 16034 27074 16046
rect 27582 16098 27634 16110
rect 37650 16046 37662 16098
rect 37714 16046 37726 16098
rect 27582 16034 27634 16046
rect 18286 15986 18338 15998
rect 18286 15922 18338 15934
rect 24446 15986 24498 15998
rect 24446 15922 24498 15934
rect 25902 15986 25954 15998
rect 25902 15922 25954 15934
rect 26686 15986 26738 15998
rect 26686 15922 26738 15934
rect 18622 15874 18674 15886
rect 18622 15810 18674 15822
rect 19182 15874 19234 15886
rect 26350 15874 26402 15886
rect 20514 15822 20526 15874
rect 20578 15822 20590 15874
rect 19182 15810 19234 15822
rect 26350 15810 26402 15822
rect 26910 15874 26962 15886
rect 26910 15810 26962 15822
rect 27694 15874 27746 15886
rect 27694 15810 27746 15822
rect 1344 15706 40656 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 40656 15706
rect 1344 15620 40656 15654
rect 15598 15538 15650 15550
rect 15598 15474 15650 15486
rect 22878 15538 22930 15550
rect 22878 15474 22930 15486
rect 23102 15538 23154 15550
rect 23102 15474 23154 15486
rect 25230 15538 25282 15550
rect 25230 15474 25282 15486
rect 26238 15538 26290 15550
rect 26238 15474 26290 15486
rect 16382 15426 16434 15438
rect 27346 15374 27358 15426
rect 27410 15374 27422 15426
rect 16382 15362 16434 15374
rect 25342 15314 25394 15326
rect 15810 15262 15822 15314
rect 15874 15262 15886 15314
rect 16146 15262 16158 15314
rect 16210 15262 16222 15314
rect 23426 15262 23438 15314
rect 23490 15262 23502 15314
rect 25342 15250 25394 15262
rect 25454 15314 25506 15326
rect 25778 15262 25790 15314
rect 25842 15262 25854 15314
rect 26562 15262 26574 15314
rect 26626 15262 26638 15314
rect 37650 15262 37662 15314
rect 37714 15262 37726 15314
rect 25454 15250 25506 15262
rect 15150 15202 15202 15214
rect 15150 15138 15202 15150
rect 15262 15202 15314 15214
rect 15262 15138 15314 15150
rect 22990 15202 23042 15214
rect 40014 15202 40066 15214
rect 29474 15150 29486 15202
rect 29538 15150 29550 15202
rect 22990 15138 23042 15150
rect 40014 15138 40066 15150
rect 15934 15090 15986 15102
rect 15934 15026 15986 15038
rect 1344 14922 40656 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 40656 14922
rect 1344 14836 40656 14870
rect 14578 14590 14590 14642
rect 14642 14590 14654 14642
rect 16706 14590 16718 14642
rect 16770 14590 16782 14642
rect 18610 14590 18622 14642
rect 18674 14590 18686 14642
rect 20738 14590 20750 14642
rect 20802 14590 20814 14642
rect 22866 14590 22878 14642
rect 22930 14590 22942 14642
rect 24994 14590 25006 14642
rect 25058 14590 25070 14642
rect 26114 14590 26126 14642
rect 26178 14590 26190 14642
rect 28242 14590 28254 14642
rect 28306 14590 28318 14642
rect 29262 14530 29314 14542
rect 13906 14478 13918 14530
rect 13970 14478 13982 14530
rect 17826 14478 17838 14530
rect 17890 14478 17902 14530
rect 22082 14478 22094 14530
rect 22146 14478 22158 14530
rect 25330 14478 25342 14530
rect 25394 14478 25406 14530
rect 29262 14466 29314 14478
rect 17502 14306 17554 14318
rect 17502 14242 17554 14254
rect 1344 14138 40656 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 40656 14138
rect 1344 14052 40656 14086
rect 16718 13970 16770 13982
rect 16718 13906 16770 13918
rect 14242 13806 14254 13858
rect 14306 13806 14318 13858
rect 27906 13806 27918 13858
rect 27970 13806 27982 13858
rect 19406 13746 19458 13758
rect 23550 13746 23602 13758
rect 13570 13694 13582 13746
rect 13634 13694 13646 13746
rect 20290 13694 20302 13746
rect 20354 13694 20366 13746
rect 19406 13682 19458 13694
rect 23550 13682 23602 13694
rect 25342 13746 25394 13758
rect 27682 13694 27694 13746
rect 27746 13694 27758 13746
rect 25342 13682 25394 13694
rect 16830 13634 16882 13646
rect 16370 13582 16382 13634
rect 16434 13582 16446 13634
rect 16830 13570 16882 13582
rect 17502 13634 17554 13646
rect 17502 13570 17554 13582
rect 19182 13634 19234 13646
rect 20962 13582 20974 13634
rect 21026 13582 21038 13634
rect 23090 13582 23102 13634
rect 23154 13582 23166 13634
rect 19182 13570 19234 13582
rect 19730 13470 19742 13522
rect 19794 13470 19806 13522
rect 1344 13354 40656 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 40656 13354
rect 1344 13268 40656 13302
rect 17166 13074 17218 13086
rect 17166 13010 17218 13022
rect 15822 12962 15874 12974
rect 16594 12910 16606 12962
rect 16658 12910 16670 12962
rect 20178 12910 20190 12962
rect 20242 12910 20254 12962
rect 15822 12898 15874 12910
rect 16158 12850 16210 12862
rect 16158 12786 16210 12798
rect 20414 12850 20466 12862
rect 20414 12786 20466 12798
rect 15934 12738 15986 12750
rect 15934 12674 15986 12686
rect 16046 12738 16098 12750
rect 16046 12674 16098 12686
rect 1344 12570 40656 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 40656 12570
rect 1344 12484 40656 12518
rect 1344 11786 40656 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 40656 11786
rect 1344 11700 40656 11734
rect 1344 11002 40656 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 40656 11002
rect 1344 10916 40656 10950
rect 1344 10218 40656 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 40656 10218
rect 1344 10132 40656 10166
rect 1344 9434 40656 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 40656 9434
rect 1344 9348 40656 9382
rect 1344 8650 40656 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 40656 8650
rect 1344 8564 40656 8598
rect 1344 7866 40656 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 40656 7866
rect 1344 7780 40656 7814
rect 1344 7082 40656 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 40656 7082
rect 1344 6996 40656 7030
rect 1344 6298 40656 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 40656 6298
rect 1344 6212 40656 6246
rect 1344 5514 40656 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 40656 5514
rect 1344 5428 40656 5462
rect 1344 4730 40656 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 40656 4730
rect 1344 4644 40656 4678
rect 17378 4286 17390 4338
rect 17442 4286 17454 4338
rect 18498 4174 18510 4226
rect 18562 4174 18574 4226
rect 1344 3946 40656 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 40656 3946
rect 1344 3860 40656 3894
rect 26126 3666 26178 3678
rect 26126 3602 26178 3614
rect 17042 3502 17054 3554
rect 17106 3502 17118 3554
rect 25218 3502 25230 3554
rect 25282 3502 25294 3554
rect 18062 3330 18114 3342
rect 18062 3266 18114 3278
rect 1344 3162 40656 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 40656 3162
rect 1344 3076 40656 3110
<< via1 >>
rect 26910 38558 26962 38610
rect 27470 38558 27522 38610
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 18622 38222 18674 38274
rect 22430 38222 22482 38274
rect 25566 38222 25618 38274
rect 17838 37998 17890 38050
rect 21534 37998 21586 38050
rect 24558 37998 24610 38050
rect 27470 37886 27522 37938
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 18398 37438 18450 37490
rect 20078 37438 20130 37490
rect 26238 37438 26290 37490
rect 19406 37214 19458 37266
rect 25230 37214 25282 37266
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 1710 36318 1762 36370
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 21982 28702 22034 28754
rect 21870 28590 21922 28642
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 19742 27918 19794 27970
rect 20862 27918 20914 27970
rect 19518 27806 19570 27858
rect 20190 27806 20242 27858
rect 23550 27806 23602 27858
rect 22990 27694 23042 27746
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 21646 27246 21698 27298
rect 19406 27134 19458 27186
rect 19854 27134 19906 27186
rect 20302 27134 20354 27186
rect 16494 27022 16546 27074
rect 21870 27022 21922 27074
rect 16158 26910 16210 26962
rect 17278 26910 17330 26962
rect 20190 26910 20242 26962
rect 20526 26910 20578 26962
rect 20750 26910 20802 26962
rect 21310 26910 21362 26962
rect 16046 26798 16098 26850
rect 19742 26798 19794 26850
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 17838 26462 17890 26514
rect 17950 26462 18002 26514
rect 4286 26238 4338 26290
rect 15150 26238 15202 26290
rect 17726 26238 17778 26290
rect 18062 26238 18114 26290
rect 18286 26238 18338 26290
rect 21870 26238 21922 26290
rect 12238 26126 12290 26178
rect 14366 26126 14418 26178
rect 15598 26126 15650 26178
rect 19630 26126 19682 26178
rect 22542 26126 22594 26178
rect 24670 26126 24722 26178
rect 25342 26126 25394 26178
rect 1934 26014 1986 26066
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 14366 25678 14418 25730
rect 15822 25566 15874 25618
rect 17950 25566 18002 25618
rect 18510 25566 18562 25618
rect 15150 25454 15202 25506
rect 18622 25454 18674 25506
rect 18846 25454 18898 25506
rect 18958 25454 19010 25506
rect 19406 25454 19458 25506
rect 14702 25342 14754 25394
rect 18398 25342 18450 25394
rect 14478 25230 14530 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 15486 24894 15538 24946
rect 15598 24894 15650 24946
rect 23662 24894 23714 24946
rect 15262 24782 15314 24834
rect 26798 24782 26850 24834
rect 27694 24782 27746 24834
rect 4286 24670 4338 24722
rect 14926 24670 14978 24722
rect 15710 24670 15762 24722
rect 15934 24670 15986 24722
rect 19406 24670 19458 24722
rect 22654 24670 22706 24722
rect 23102 24670 23154 24722
rect 23438 24670 23490 24722
rect 26462 24670 26514 24722
rect 27022 24670 27074 24722
rect 27358 24670 27410 24722
rect 37886 24670 37938 24722
rect 12014 24558 12066 24610
rect 14142 24558 14194 24610
rect 16382 24558 16434 24610
rect 18174 24558 18226 24610
rect 20078 24558 20130 24610
rect 22206 24558 22258 24610
rect 23550 24558 23602 24610
rect 1934 24446 1986 24498
rect 27134 24446 27186 24498
rect 40014 24446 40066 24498
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 28030 24110 28082 24162
rect 1934 23998 1986 24050
rect 14814 23998 14866 24050
rect 19854 23998 19906 24050
rect 21422 23998 21474 24050
rect 22990 23998 23042 24050
rect 26686 23998 26738 24050
rect 27134 23998 27186 24050
rect 40014 23998 40066 24050
rect 4286 23886 4338 23938
rect 14142 23886 14194 23938
rect 14926 23886 14978 23938
rect 19966 23886 20018 23938
rect 20190 23886 20242 23938
rect 20414 23886 20466 23938
rect 21534 23886 21586 23938
rect 22654 23886 22706 23938
rect 23774 23886 23826 23938
rect 37662 23886 37714 23938
rect 14366 23774 14418 23826
rect 14478 23774 14530 23826
rect 15262 23774 15314 23826
rect 19742 23774 19794 23826
rect 20638 23774 20690 23826
rect 21310 23774 21362 23826
rect 21758 23774 21810 23826
rect 22206 23774 22258 23826
rect 23214 23774 23266 23826
rect 23326 23774 23378 23826
rect 23438 23774 23490 23826
rect 24558 23774 24610 23826
rect 27022 23774 27074 23826
rect 27358 23774 27410 23826
rect 27582 23774 27634 23826
rect 27918 23774 27970 23826
rect 28030 23774 28082 23826
rect 15374 23662 15426 23714
rect 15598 23662 15650 23714
rect 18062 23662 18114 23714
rect 18398 23662 18450 23714
rect 18734 23662 18786 23714
rect 19070 23662 19122 23714
rect 22318 23662 22370 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 12238 23326 12290 23378
rect 17726 23326 17778 23378
rect 18398 23326 18450 23378
rect 21982 23326 22034 23378
rect 22094 23326 22146 23378
rect 22878 23326 22930 23378
rect 25454 23326 25506 23378
rect 26350 23326 26402 23378
rect 15374 23214 15426 23266
rect 18622 23214 18674 23266
rect 20638 23214 20690 23266
rect 23550 23214 23602 23266
rect 24334 23214 24386 23266
rect 26462 23214 26514 23266
rect 27582 23214 27634 23266
rect 4286 23102 4338 23154
rect 12462 23102 12514 23154
rect 15262 23102 15314 23154
rect 15598 23102 15650 23154
rect 17614 23102 17666 23154
rect 17838 23102 17890 23154
rect 18286 23102 18338 23154
rect 18958 23102 19010 23154
rect 19406 23102 19458 23154
rect 19854 23102 19906 23154
rect 20862 23102 20914 23154
rect 22206 23102 22258 23154
rect 22654 23102 22706 23154
rect 22878 23102 22930 23154
rect 23102 23102 23154 23154
rect 23326 23102 23378 23154
rect 23774 23102 23826 23154
rect 24110 23102 24162 23154
rect 26126 23102 26178 23154
rect 26798 23102 26850 23154
rect 37662 23102 37714 23154
rect 13022 22990 13074 23042
rect 25230 22990 25282 23042
rect 25454 22990 25506 23042
rect 29710 22990 29762 23042
rect 1934 22878 1986 22930
rect 24446 22878 24498 22930
rect 40014 22878 40066 22930
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 17278 22542 17330 22594
rect 19630 22542 19682 22594
rect 20414 22542 20466 22594
rect 1934 22430 1986 22482
rect 9886 22430 9938 22482
rect 21870 22430 21922 22482
rect 28590 22430 28642 22482
rect 29262 22430 29314 22482
rect 4286 22318 4338 22370
rect 12798 22318 12850 22370
rect 13694 22318 13746 22370
rect 14478 22318 14530 22370
rect 15150 22318 15202 22370
rect 15598 22318 15650 22370
rect 15822 22318 15874 22370
rect 17838 22318 17890 22370
rect 19070 22318 19122 22370
rect 19294 22318 19346 22370
rect 20078 22318 20130 22370
rect 21310 22318 21362 22370
rect 23438 22318 23490 22370
rect 25790 22318 25842 22370
rect 12014 22206 12066 22258
rect 13470 22206 13522 22258
rect 14926 22206 14978 22258
rect 15038 22206 15090 22258
rect 15262 22206 15314 22258
rect 15934 22206 15986 22258
rect 17166 22206 17218 22258
rect 17278 22206 17330 22258
rect 18734 22206 18786 22258
rect 19518 22206 19570 22258
rect 19854 22206 19906 22258
rect 21422 22206 21474 22258
rect 25118 22206 25170 22258
rect 26462 22206 26514 22258
rect 16046 22094 16098 22146
rect 16158 22094 16210 22146
rect 16830 22094 16882 22146
rect 18062 22094 18114 22146
rect 18398 22094 18450 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 15038 21758 15090 21810
rect 17950 21758 18002 21810
rect 25342 21758 25394 21810
rect 25566 21758 25618 21810
rect 26462 21758 26514 21810
rect 26910 21758 26962 21810
rect 27358 21758 27410 21810
rect 14142 21646 14194 21698
rect 14478 21646 14530 21698
rect 14702 21646 14754 21698
rect 15822 21646 15874 21698
rect 16270 21646 16322 21698
rect 25230 21646 25282 21698
rect 4286 21534 4338 21586
rect 13470 21534 13522 21586
rect 15262 21534 15314 21586
rect 15598 21534 15650 21586
rect 16494 21534 16546 21586
rect 17726 21534 17778 21586
rect 18958 21534 19010 21586
rect 19294 21534 19346 21586
rect 26014 21534 26066 21586
rect 26238 21534 26290 21586
rect 26574 21534 26626 21586
rect 27022 21534 27074 21586
rect 27134 21534 27186 21586
rect 1934 21422 1986 21474
rect 10670 21422 10722 21474
rect 12798 21422 12850 21474
rect 14254 21422 14306 21474
rect 18510 21422 18562 21474
rect 22878 21422 22930 21474
rect 15262 21310 15314 21362
rect 16158 21310 16210 21362
rect 18062 21310 18114 21362
rect 26014 21310 26066 21362
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 22206 20974 22258 21026
rect 26798 20862 26850 20914
rect 40014 20862 40066 20914
rect 13918 20750 13970 20802
rect 14478 20750 14530 20802
rect 15038 20750 15090 20802
rect 20078 20750 20130 20802
rect 21870 20750 21922 20802
rect 22878 20750 22930 20802
rect 37662 20750 37714 20802
rect 14814 20638 14866 20690
rect 17838 20638 17890 20690
rect 21646 20638 21698 20690
rect 22094 20638 22146 20690
rect 13582 20526 13634 20578
rect 13806 20526 13858 20578
rect 14142 20526 14194 20578
rect 14366 20526 14418 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 20190 20190 20242 20242
rect 23550 20190 23602 20242
rect 26350 20190 26402 20242
rect 15822 20078 15874 20130
rect 17950 20078 18002 20130
rect 18734 20078 18786 20130
rect 19854 20078 19906 20130
rect 20526 20078 20578 20130
rect 22430 20078 22482 20130
rect 24222 20078 24274 20130
rect 25566 20078 25618 20130
rect 16046 19966 16098 20018
rect 16382 19966 16434 20018
rect 18286 19966 18338 20018
rect 18622 19966 18674 20018
rect 19630 19966 19682 20018
rect 21534 19966 21586 20018
rect 22094 19966 22146 20018
rect 22654 19966 22706 20018
rect 22990 19966 23042 20018
rect 23214 19966 23266 20018
rect 23886 19966 23938 20018
rect 25790 19966 25842 20018
rect 26798 19966 26850 20018
rect 13806 19854 13858 19906
rect 19294 19854 19346 19906
rect 27470 19854 27522 19906
rect 29598 19854 29650 19906
rect 15710 19742 15762 19794
rect 22766 19742 22818 19794
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 18734 19406 18786 19458
rect 23550 19406 23602 19458
rect 19070 19294 19122 19346
rect 19518 19294 19570 19346
rect 21310 19294 21362 19346
rect 23102 19294 23154 19346
rect 26798 19294 26850 19346
rect 14030 19182 14082 19234
rect 14702 19182 14754 19234
rect 15150 19182 15202 19234
rect 17614 19182 17666 19234
rect 18622 19182 18674 19234
rect 19406 19182 19458 19234
rect 21758 19182 21810 19234
rect 22542 19182 22594 19234
rect 22878 19182 22930 19234
rect 25678 19182 25730 19234
rect 26574 19182 26626 19234
rect 27022 19182 27074 19234
rect 27134 19182 27186 19234
rect 27806 19182 27858 19234
rect 16606 19070 16658 19122
rect 17278 19070 17330 19122
rect 22206 19070 22258 19122
rect 23214 19070 23266 19122
rect 23662 19070 23714 19122
rect 25342 19070 25394 19122
rect 27582 19070 27634 19122
rect 28142 19070 28194 19122
rect 14478 18958 14530 19010
rect 14590 18958 14642 19010
rect 16942 18958 16994 19010
rect 25454 18958 25506 19010
rect 25902 18958 25954 19010
rect 26238 18958 26290 19010
rect 27918 18958 27970 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 15486 18622 15538 18674
rect 17950 18622 18002 18674
rect 21422 18622 21474 18674
rect 23326 18622 23378 18674
rect 25454 18622 25506 18674
rect 26238 18622 26290 18674
rect 14590 18510 14642 18562
rect 16158 18510 16210 18562
rect 20862 18510 20914 18562
rect 25230 18510 25282 18562
rect 27358 18510 27410 18562
rect 4286 18398 4338 18450
rect 11454 18398 11506 18450
rect 12126 18398 12178 18450
rect 14926 18398 14978 18450
rect 15150 18398 15202 18450
rect 15710 18398 15762 18450
rect 16494 18398 16546 18450
rect 17726 18398 17778 18450
rect 18286 18398 18338 18450
rect 18510 18398 18562 18450
rect 19742 18398 19794 18450
rect 20414 18398 20466 18450
rect 21422 18398 21474 18450
rect 21982 18398 22034 18450
rect 22094 18398 22146 18450
rect 22430 18398 22482 18450
rect 23998 18398 24050 18450
rect 24670 18398 24722 18450
rect 25790 18398 25842 18450
rect 26574 18398 26626 18450
rect 37662 18398 37714 18450
rect 14254 18286 14306 18338
rect 14702 18286 14754 18338
rect 19406 18286 19458 18338
rect 23774 18286 23826 18338
rect 29486 18286 29538 18338
rect 1934 18174 1986 18226
rect 18846 18174 18898 18226
rect 19966 18174 20018 18226
rect 22654 18174 22706 18226
rect 22878 18174 22930 18226
rect 25566 18174 25618 18226
rect 40014 18174 40066 18226
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 15262 17726 15314 17778
rect 17390 17726 17442 17778
rect 20414 17726 20466 17778
rect 22206 17726 22258 17778
rect 14478 17614 14530 17666
rect 18734 17614 18786 17666
rect 20638 17614 20690 17666
rect 21758 17614 21810 17666
rect 23214 17614 23266 17666
rect 23998 17614 24050 17666
rect 27918 17614 27970 17666
rect 19742 17502 19794 17554
rect 23438 17502 23490 17554
rect 27582 17502 27634 17554
rect 27694 17502 27746 17554
rect 17838 17390 17890 17442
rect 19070 17390 19122 17442
rect 20078 17390 20130 17442
rect 23774 17390 23826 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 14478 17054 14530 17106
rect 18734 17054 18786 17106
rect 21086 17054 21138 17106
rect 21422 17054 21474 17106
rect 27358 17054 27410 17106
rect 13246 16942 13298 16994
rect 27246 16942 27298 16994
rect 14030 16830 14082 16882
rect 19070 16830 19122 16882
rect 27134 16830 27186 16882
rect 27694 16830 27746 16882
rect 37886 16830 37938 16882
rect 11118 16718 11170 16770
rect 39902 16718 39954 16770
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 27694 16270 27746 16322
rect 19966 16158 20018 16210
rect 40014 16158 40066 16210
rect 18510 16046 18562 16098
rect 18734 16046 18786 16098
rect 19070 16046 19122 16098
rect 19294 16046 19346 16098
rect 19518 16046 19570 16098
rect 20190 16046 20242 16098
rect 24110 16046 24162 16098
rect 26126 16046 26178 16098
rect 26574 16046 26626 16098
rect 27022 16046 27074 16098
rect 27582 16046 27634 16098
rect 37662 16046 37714 16098
rect 18286 15934 18338 15986
rect 24446 15934 24498 15986
rect 25902 15934 25954 15986
rect 26686 15934 26738 15986
rect 18622 15822 18674 15874
rect 19182 15822 19234 15874
rect 20526 15822 20578 15874
rect 26350 15822 26402 15874
rect 26910 15822 26962 15874
rect 27694 15822 27746 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 15598 15486 15650 15538
rect 22878 15486 22930 15538
rect 23102 15486 23154 15538
rect 25230 15486 25282 15538
rect 26238 15486 26290 15538
rect 16382 15374 16434 15426
rect 27358 15374 27410 15426
rect 15822 15262 15874 15314
rect 16158 15262 16210 15314
rect 23438 15262 23490 15314
rect 25342 15262 25394 15314
rect 25454 15262 25506 15314
rect 25790 15262 25842 15314
rect 26574 15262 26626 15314
rect 37662 15262 37714 15314
rect 15150 15150 15202 15202
rect 15262 15150 15314 15202
rect 22990 15150 23042 15202
rect 29486 15150 29538 15202
rect 40014 15150 40066 15202
rect 15934 15038 15986 15090
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 14590 14590 14642 14642
rect 16718 14590 16770 14642
rect 18622 14590 18674 14642
rect 20750 14590 20802 14642
rect 22878 14590 22930 14642
rect 25006 14590 25058 14642
rect 26126 14590 26178 14642
rect 28254 14590 28306 14642
rect 13918 14478 13970 14530
rect 17838 14478 17890 14530
rect 22094 14478 22146 14530
rect 25342 14478 25394 14530
rect 29262 14478 29314 14530
rect 17502 14254 17554 14306
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 16718 13918 16770 13970
rect 14254 13806 14306 13858
rect 27918 13806 27970 13858
rect 13582 13694 13634 13746
rect 19406 13694 19458 13746
rect 20302 13694 20354 13746
rect 23550 13694 23602 13746
rect 25342 13694 25394 13746
rect 27694 13694 27746 13746
rect 16382 13582 16434 13634
rect 16830 13582 16882 13634
rect 17502 13582 17554 13634
rect 19182 13582 19234 13634
rect 20974 13582 21026 13634
rect 23102 13582 23154 13634
rect 19742 13470 19794 13522
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 17166 13022 17218 13074
rect 15822 12910 15874 12962
rect 16606 12910 16658 12962
rect 20190 12910 20242 12962
rect 16158 12798 16210 12850
rect 20414 12798 20466 12850
rect 15934 12686 15986 12738
rect 16046 12686 16098 12738
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 17390 4286 17442 4338
rect 18510 4174 18562 4226
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 26126 3614 26178 3666
rect 17054 3502 17106 3554
rect 25230 3502 25282 3554
rect 18062 3278 18114 3330
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
<< metal2 >>
rect 17472 41200 17584 42000
rect 18144 41200 18256 42000
rect 18816 41200 18928 42000
rect 22176 41200 22288 42000
rect 22848 41200 22960 42000
rect 24864 41200 24976 42000
rect 26880 41200 26992 42000
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 17500 38276 17556 41200
rect 17500 38210 17556 38220
rect 17836 38050 17892 38062
rect 17836 37998 17838 38050
rect 17890 37998 17892 38050
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 1708 36372 1764 36382
rect 1708 36278 1764 36316
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 4172 28308 4228 28318
rect 1932 26066 1988 26078
rect 1932 26014 1934 26066
rect 1986 26014 1988 26066
rect 1932 25620 1988 26014
rect 1932 25554 1988 25564
rect 1932 24500 1988 24510
rect 1932 24406 1988 24444
rect 1932 24050 1988 24062
rect 1932 23998 1934 24050
rect 1986 23998 1988 24050
rect 1932 23604 1988 23998
rect 1932 23538 1988 23548
rect 1932 22932 1988 22942
rect 1932 22838 1988 22876
rect 1932 22484 1988 22494
rect 1932 22390 1988 22428
rect 4172 22148 4228 28252
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 16492 27076 16548 27086
rect 16380 27074 16548 27076
rect 16380 27022 16494 27074
rect 16546 27022 16548 27074
rect 16380 27020 16548 27022
rect 16156 26962 16212 26974
rect 16156 26910 16158 26962
rect 16210 26910 16212 26962
rect 16044 26850 16100 26862
rect 16044 26798 16046 26850
rect 16098 26798 16100 26850
rect 4284 26292 4340 26302
rect 4284 26198 4340 26236
rect 12236 26292 12292 26302
rect 12236 26178 12292 26236
rect 15148 26290 15204 26302
rect 15148 26238 15150 26290
rect 15202 26238 15204 26290
rect 12236 26126 12238 26178
rect 12290 26126 12292 26178
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 12236 25732 12292 26126
rect 12236 25666 12292 25676
rect 14364 26178 14420 26190
rect 14364 26126 14366 26178
rect 14418 26126 14420 26178
rect 14364 25730 14420 26126
rect 14364 25678 14366 25730
rect 14418 25678 14420 25730
rect 14364 25666 14420 25678
rect 15148 26180 15204 26238
rect 15596 26180 15652 26190
rect 15148 26178 15652 26180
rect 15148 26126 15598 26178
rect 15650 26126 15652 26178
rect 15148 26124 15652 26126
rect 15148 25506 15204 26124
rect 15596 26114 15652 26124
rect 15148 25454 15150 25506
rect 15202 25454 15204 25506
rect 14700 25396 14756 25406
rect 14700 25302 14756 25340
rect 14476 25282 14532 25294
rect 14476 25230 14478 25282
rect 14530 25230 14532 25282
rect 14476 24948 14532 25230
rect 14476 24882 14532 24892
rect 4284 24724 4340 24734
rect 4284 24630 4340 24668
rect 12012 24724 12068 24734
rect 12012 24610 12068 24668
rect 14812 24724 14868 24734
rect 12012 24558 12014 24610
rect 12066 24558 12068 24610
rect 12012 24546 12068 24558
rect 14140 24610 14196 24622
rect 14140 24558 14142 24610
rect 14194 24558 14196 24610
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 4284 23940 4340 23950
rect 4284 23846 4340 23884
rect 12236 23940 12292 23950
rect 12236 23378 12292 23884
rect 14140 23938 14196 24558
rect 14812 24388 14868 24668
rect 14924 24724 14980 24734
rect 15148 24724 15204 25454
rect 15260 25732 15316 25742
rect 15260 24834 15316 25676
rect 15820 25620 15876 25630
rect 16044 25620 16100 26798
rect 16156 26516 16212 26910
rect 16156 26450 16212 26460
rect 15820 25618 16100 25620
rect 15820 25566 15822 25618
rect 15874 25566 16100 25618
rect 15820 25564 16100 25566
rect 15820 25554 15876 25564
rect 15484 25508 15540 25518
rect 15484 24946 15540 25452
rect 15484 24894 15486 24946
rect 15538 24894 15540 24946
rect 15484 24882 15540 24894
rect 15596 24948 15652 24958
rect 15596 24854 15652 24892
rect 15260 24782 15262 24834
rect 15314 24782 15316 24834
rect 15260 24770 15316 24782
rect 14924 24722 15204 24724
rect 14924 24670 14926 24722
rect 14978 24670 15204 24722
rect 14924 24668 15204 24670
rect 15708 24722 15764 24734
rect 15708 24670 15710 24722
rect 15762 24670 15764 24722
rect 14924 24612 14980 24668
rect 14924 24546 14980 24556
rect 14812 24332 14980 24388
rect 14812 24052 14868 24062
rect 14140 23886 14142 23938
rect 14194 23886 14196 23938
rect 14140 23874 14196 23886
rect 14364 24050 14868 24052
rect 14364 23998 14814 24050
rect 14866 23998 14868 24050
rect 14364 23996 14868 23998
rect 14364 23826 14420 23996
rect 14812 23986 14868 23996
rect 14924 23938 14980 24332
rect 15708 23940 15764 24670
rect 14924 23886 14926 23938
rect 14978 23886 14980 23938
rect 14924 23874 14980 23886
rect 15484 23884 15764 23940
rect 15932 24722 15988 24734
rect 15932 24670 15934 24722
rect 15986 24670 15988 24722
rect 14364 23774 14366 23826
rect 14418 23774 14420 23826
rect 14364 23762 14420 23774
rect 14476 23826 14532 23838
rect 15260 23828 15316 23838
rect 14476 23774 14478 23826
rect 14530 23774 14532 23826
rect 12236 23326 12238 23378
rect 12290 23326 12292 23378
rect 12236 23314 12292 23326
rect 14476 23380 14532 23774
rect 14476 23314 14532 23324
rect 15148 23826 15316 23828
rect 15148 23774 15262 23826
rect 15314 23774 15316 23826
rect 15148 23772 15316 23774
rect 4284 23154 4340 23166
rect 4284 23102 4286 23154
rect 4338 23102 4340 23154
rect 4284 23044 4340 23102
rect 4284 22978 4340 22988
rect 12460 23154 12516 23166
rect 12460 23102 12462 23154
rect 12514 23102 12516 23154
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 9884 22482 9940 22494
rect 9884 22430 9886 22482
rect 9938 22430 9940 22482
rect 4284 22372 4340 22382
rect 4284 22278 4340 22316
rect 9884 22372 9940 22430
rect 9884 22306 9940 22316
rect 12460 22372 12516 23102
rect 13020 23042 13076 23054
rect 13020 22990 13022 23042
rect 13074 22990 13076 23042
rect 12460 22306 12516 22316
rect 12796 22372 12852 22382
rect 13020 22372 13076 22990
rect 12796 22370 13076 22372
rect 12796 22318 12798 22370
rect 12850 22318 13076 22370
rect 12796 22316 13076 22318
rect 13468 23044 13524 23054
rect 12012 22260 12068 22270
rect 12012 22166 12068 22204
rect 4172 22082 4228 22092
rect 12796 21812 12852 22316
rect 13468 22258 13524 22988
rect 14140 22820 14196 22830
rect 13692 22372 13748 22382
rect 13692 22278 13748 22316
rect 13468 22206 13470 22258
rect 13522 22206 13524 22258
rect 13468 22194 13524 22206
rect 12796 21746 12852 21756
rect 13468 21812 13524 21822
rect 4284 21588 4340 21598
rect 4284 21494 4340 21532
rect 13468 21586 13524 21756
rect 14140 21700 14196 22764
rect 14924 22596 14980 22606
rect 15148 22596 15204 23772
rect 15260 23762 15316 23772
rect 15372 23716 15428 23726
rect 15484 23716 15540 23884
rect 15372 23714 15540 23716
rect 15372 23662 15374 23714
rect 15426 23662 15540 23714
rect 15372 23660 15540 23662
rect 15596 23716 15652 23726
rect 15372 23492 15428 23660
rect 15596 23622 15652 23660
rect 15372 23426 15428 23436
rect 15372 23266 15428 23278
rect 15372 23214 15374 23266
rect 15426 23214 15428 23266
rect 14980 22540 15204 22596
rect 15260 23154 15316 23166
rect 15260 23102 15262 23154
rect 15314 23102 15316 23154
rect 15260 22596 15316 23102
rect 15372 23044 15428 23214
rect 15596 23156 15652 23166
rect 15596 23154 15876 23156
rect 15596 23102 15598 23154
rect 15650 23102 15876 23154
rect 15596 23100 15876 23102
rect 15596 23090 15652 23100
rect 15372 22978 15428 22988
rect 15260 22540 15764 22596
rect 14476 22372 14532 22382
rect 14476 22278 14532 22316
rect 14924 22258 14980 22540
rect 15148 22428 15652 22484
rect 14924 22206 14926 22258
rect 14978 22206 14980 22258
rect 14924 22194 14980 22206
rect 15036 22372 15092 22382
rect 15036 22258 15092 22316
rect 15148 22370 15204 22428
rect 15148 22318 15150 22370
rect 15202 22318 15204 22370
rect 15148 22306 15204 22318
rect 15596 22370 15652 22428
rect 15596 22318 15598 22370
rect 15650 22318 15652 22370
rect 15596 22306 15652 22318
rect 15036 22206 15038 22258
rect 15090 22206 15092 22258
rect 15036 22194 15092 22206
rect 15260 22260 15316 22270
rect 15260 22258 15540 22260
rect 15260 22206 15262 22258
rect 15314 22206 15540 22258
rect 15260 22204 15540 22206
rect 15260 22194 15316 22204
rect 14588 22036 14644 22046
rect 13468 21534 13470 21586
rect 13522 21534 13524 21586
rect 1932 21476 1988 21486
rect 1932 21382 1988 21420
rect 10668 21474 10724 21486
rect 10668 21422 10670 21474
rect 10722 21422 10724 21474
rect 10668 21364 10724 21422
rect 12796 21476 12852 21486
rect 12796 21382 12852 21420
rect 10668 21298 10724 21308
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 12124 20132 12180 20142
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 4284 18452 4340 18462
rect 4284 18358 4340 18396
rect 11452 18452 11508 18462
rect 11452 18358 11508 18396
rect 12124 18450 12180 20076
rect 13468 19908 13524 21534
rect 13916 21698 14196 21700
rect 13916 21646 14142 21698
rect 14194 21646 14196 21698
rect 13916 21644 14196 21646
rect 13916 20802 13972 21644
rect 14140 21634 14196 21644
rect 14476 21924 14532 21934
rect 14476 21698 14532 21868
rect 14476 21646 14478 21698
rect 14530 21646 14532 21698
rect 14476 21634 14532 21646
rect 14252 21476 14308 21486
rect 14252 21382 14308 21420
rect 13916 20750 13918 20802
rect 13970 20750 13972 20802
rect 13916 20738 13972 20750
rect 14476 20804 14532 20814
rect 14588 20804 14644 21980
rect 15036 21812 15092 21822
rect 14700 21810 15092 21812
rect 14700 21758 15038 21810
rect 15090 21758 15092 21810
rect 14700 21756 15092 21758
rect 14700 21698 14756 21756
rect 15036 21746 15092 21756
rect 14700 21646 14702 21698
rect 14754 21646 14756 21698
rect 14700 21634 14756 21646
rect 15260 21588 15316 21598
rect 15260 21586 15428 21588
rect 15260 21534 15262 21586
rect 15314 21534 15428 21586
rect 15260 21532 15428 21534
rect 15260 21522 15316 21532
rect 15260 21364 15316 21374
rect 15260 21270 15316 21308
rect 14476 20802 14644 20804
rect 14476 20750 14478 20802
rect 14530 20750 14644 20802
rect 14476 20748 14644 20750
rect 14476 20738 14532 20748
rect 14588 20692 14644 20748
rect 15036 20802 15092 20814
rect 15036 20750 15038 20802
rect 15090 20750 15092 20802
rect 14812 20692 14868 20702
rect 14588 20690 14868 20692
rect 14588 20638 14814 20690
rect 14866 20638 14868 20690
rect 14588 20636 14868 20638
rect 14812 20626 14868 20636
rect 13580 20578 13636 20590
rect 13580 20526 13582 20578
rect 13634 20526 13636 20578
rect 13580 20132 13636 20526
rect 13804 20578 13860 20590
rect 14140 20580 14196 20590
rect 13804 20526 13806 20578
rect 13858 20526 13860 20578
rect 13804 20468 13860 20526
rect 14028 20578 14196 20580
rect 14028 20526 14142 20578
rect 14194 20526 14196 20578
rect 14028 20524 14196 20526
rect 14028 20468 14084 20524
rect 14140 20514 14196 20524
rect 14364 20578 14420 20590
rect 14364 20526 14366 20578
rect 14418 20526 14420 20578
rect 13804 20412 14084 20468
rect 14364 20356 14420 20526
rect 14364 20300 14532 20356
rect 13580 20066 13636 20076
rect 14476 20132 14532 20300
rect 14476 20066 14532 20076
rect 13804 19908 13860 19918
rect 13468 19906 13860 19908
rect 13468 19854 13806 19906
rect 13858 19854 13860 19906
rect 13468 19852 13860 19854
rect 13804 18564 13860 19852
rect 14924 19796 14980 19806
rect 14700 19572 14756 19582
rect 13804 18498 13860 18508
rect 14028 19234 14084 19246
rect 14028 19182 14030 19234
rect 14082 19182 14084 19234
rect 12124 18398 12126 18450
rect 12178 18398 12180 18450
rect 12124 18386 12180 18398
rect 13244 18340 13300 18350
rect 1932 18228 1988 18238
rect 1932 18134 1988 18172
rect 11116 18116 11172 18126
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 11116 16770 11172 18060
rect 13244 16994 13300 18284
rect 14028 18116 14084 19182
rect 14700 19234 14756 19516
rect 14700 19182 14702 19234
rect 14754 19182 14756 19234
rect 14700 19170 14756 19182
rect 14476 19012 14532 19022
rect 14364 19010 14532 19012
rect 14364 18958 14478 19010
rect 14530 18958 14532 19010
rect 14364 18956 14532 18958
rect 14364 18452 14420 18956
rect 14476 18946 14532 18956
rect 14588 19010 14644 19022
rect 14588 18958 14590 19010
rect 14642 18958 14644 19010
rect 14364 18386 14420 18396
rect 14476 18564 14532 18574
rect 14252 18338 14308 18350
rect 14252 18286 14254 18338
rect 14306 18286 14308 18338
rect 14252 18228 14308 18286
rect 14252 18162 14308 18172
rect 14028 18050 14084 18060
rect 14476 17666 14532 18508
rect 14588 18562 14644 18958
rect 14588 18510 14590 18562
rect 14642 18510 14644 18562
rect 14588 18498 14644 18510
rect 14924 18450 14980 19740
rect 15036 19348 15092 20750
rect 15036 19282 15092 19292
rect 15148 19236 15204 19246
rect 15148 18676 15204 19180
rect 15148 18610 15204 18620
rect 15260 19124 15316 19134
rect 14924 18398 14926 18450
rect 14978 18398 14980 18450
rect 14924 18386 14980 18398
rect 15148 18452 15204 18462
rect 15148 18358 15204 18396
rect 14700 18340 14756 18350
rect 14700 18246 14756 18284
rect 15260 17778 15316 19068
rect 15372 18004 15428 21532
rect 15484 19572 15540 22204
rect 15708 21700 15764 22540
rect 15820 22370 15876 23100
rect 15932 23044 15988 24670
rect 16380 24612 16436 27020
rect 16492 27010 16548 27020
rect 17276 26962 17332 26974
rect 17276 26910 17278 26962
rect 17330 26910 17332 26962
rect 17276 25620 17332 26910
rect 17836 26514 17892 37998
rect 18172 37492 18228 41200
rect 18620 38276 18676 38286
rect 18620 38182 18676 38220
rect 18396 37492 18452 37502
rect 18172 37490 18452 37492
rect 18172 37438 18398 37490
rect 18450 37438 18452 37490
rect 18172 37436 18452 37438
rect 18396 37426 18452 37436
rect 18844 37492 18900 41200
rect 22204 38276 22260 41200
rect 22428 38276 22484 38286
rect 22204 38274 22484 38276
rect 22204 38222 22430 38274
rect 22482 38222 22484 38274
rect 22204 38220 22484 38222
rect 22428 38210 22484 38220
rect 22876 38276 22932 41200
rect 22876 38210 22932 38220
rect 21532 38050 21588 38062
rect 21532 37998 21534 38050
rect 21586 37998 21588 38050
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 18844 37426 18900 37436
rect 20076 37492 20132 37502
rect 20076 37398 20132 37436
rect 19404 37266 19460 37278
rect 19404 37214 19406 37266
rect 19458 37214 19460 37266
rect 19404 27188 19460 37214
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 20524 28644 20580 28654
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 19740 27972 19796 27982
rect 19740 27878 19796 27916
rect 19516 27858 19572 27870
rect 19516 27806 19518 27858
rect 19570 27806 19572 27858
rect 19516 27412 19572 27806
rect 20188 27860 20244 27870
rect 20188 27766 20244 27804
rect 20412 27524 20468 27534
rect 19516 27346 19572 27356
rect 20300 27468 20412 27524
rect 19852 27188 19908 27198
rect 19404 27186 19908 27188
rect 19404 27134 19406 27186
rect 19458 27134 19854 27186
rect 19906 27134 19908 27186
rect 19404 27132 19908 27134
rect 19404 27122 19460 27132
rect 19852 27122 19908 27132
rect 20300 27186 20356 27468
rect 20412 27458 20468 27468
rect 20300 27134 20302 27186
rect 20354 27134 20356 27186
rect 20300 27122 20356 27134
rect 20188 26962 20244 26974
rect 20188 26910 20190 26962
rect 20242 26910 20244 26962
rect 19740 26852 19796 26862
rect 19516 26850 19796 26852
rect 19516 26798 19742 26850
rect 19794 26798 19796 26850
rect 19516 26796 19796 26798
rect 17836 26462 17838 26514
rect 17890 26462 17892 26514
rect 17276 25554 17332 25564
rect 17724 26290 17780 26302
rect 17724 26238 17726 26290
rect 17778 26238 17780 26290
rect 17724 25508 17780 26238
rect 17836 25620 17892 26462
rect 17948 26516 18004 26526
rect 17948 26422 18004 26460
rect 18060 26290 18116 26302
rect 18060 26238 18062 26290
rect 18114 26238 18116 26290
rect 17948 25620 18004 25630
rect 17836 25618 18004 25620
rect 17836 25566 17950 25618
rect 18002 25566 18004 25618
rect 17836 25564 18004 25566
rect 17948 25554 18004 25564
rect 17724 25442 17780 25452
rect 18060 24836 18116 26238
rect 18284 26292 18340 26302
rect 18284 26290 18452 26292
rect 18284 26238 18286 26290
rect 18338 26238 18452 26290
rect 18284 26236 18452 26238
rect 18284 26226 18340 26236
rect 17724 24780 18116 24836
rect 18396 25394 18452 26236
rect 18508 25620 18564 25630
rect 18508 25526 18564 25564
rect 18620 25508 18676 25518
rect 18620 25506 18788 25508
rect 18620 25454 18622 25506
rect 18674 25454 18788 25506
rect 18620 25452 18788 25454
rect 18620 25442 18676 25452
rect 18396 25342 18398 25394
rect 18450 25342 18452 25394
rect 16380 24518 16436 24556
rect 16940 24612 16996 24622
rect 16156 23604 16212 23614
rect 15932 22978 15988 22988
rect 16044 23492 16100 23502
rect 15820 22318 15822 22370
rect 15874 22318 15876 22370
rect 15820 22306 15876 22318
rect 15932 22260 15988 22270
rect 15932 22166 15988 22204
rect 16044 22146 16100 23436
rect 16044 22094 16046 22146
rect 16098 22094 16100 22146
rect 16044 22036 16100 22094
rect 16044 21970 16100 21980
rect 16156 22146 16212 23548
rect 16156 22094 16158 22146
rect 16210 22094 16212 22146
rect 16156 21924 16212 22094
rect 16156 21858 16212 21868
rect 16380 23044 16436 23054
rect 15820 21700 15876 21710
rect 16268 21700 16324 21710
rect 15708 21698 16324 21700
rect 15708 21646 15822 21698
rect 15874 21646 16270 21698
rect 16322 21646 16324 21698
rect 15708 21644 16324 21646
rect 15820 21634 15876 21644
rect 16268 21634 16324 21644
rect 15596 21586 15652 21598
rect 15596 21534 15598 21586
rect 15650 21534 15652 21586
rect 15596 20020 15652 21534
rect 16156 21362 16212 21374
rect 16156 21310 16158 21362
rect 16210 21310 16212 21362
rect 16156 21252 16212 21310
rect 16156 21186 16212 21196
rect 15596 19954 15652 19964
rect 15820 20132 15876 20142
rect 15708 19796 15764 19806
rect 15708 19702 15764 19740
rect 15484 19506 15540 19516
rect 15484 19348 15540 19358
rect 15484 19012 15540 19292
rect 15820 19124 15876 20076
rect 16044 20018 16100 20030
rect 16044 19966 16046 20018
rect 16098 19966 16100 20018
rect 16044 19908 16100 19966
rect 16380 20018 16436 22988
rect 16604 22372 16660 22382
rect 16380 19966 16382 20018
rect 16434 19966 16436 20018
rect 16380 19954 16436 19966
rect 16492 21586 16548 21598
rect 16492 21534 16494 21586
rect 16546 21534 16548 21586
rect 16044 19842 16100 19852
rect 16492 19796 16548 21534
rect 16492 19730 16548 19740
rect 16604 21252 16660 22316
rect 16828 22148 16884 22158
rect 16828 21588 16884 22092
rect 16828 21522 16884 21532
rect 15820 19058 15876 19068
rect 16380 19348 16436 19358
rect 15484 18674 15540 18956
rect 15484 18622 15486 18674
rect 15538 18622 15540 18674
rect 15484 18610 15540 18622
rect 16156 18562 16212 18574
rect 16156 18510 16158 18562
rect 16210 18510 16212 18562
rect 15708 18450 15764 18462
rect 15708 18398 15710 18450
rect 15762 18398 15764 18450
rect 15708 18228 15764 18398
rect 15708 18162 15764 18172
rect 16156 18452 16212 18510
rect 15372 17938 15428 17948
rect 15260 17726 15262 17778
rect 15314 17726 15316 17778
rect 15260 17714 15316 17726
rect 14476 17614 14478 17666
rect 14530 17614 14532 17666
rect 14476 17108 14532 17614
rect 13244 16942 13246 16994
rect 13298 16942 13300 16994
rect 13244 16930 13300 16942
rect 14028 17106 14532 17108
rect 14028 17054 14478 17106
rect 14530 17054 14532 17106
rect 14028 17052 14532 17054
rect 11116 16718 11118 16770
rect 11170 16718 11172 16770
rect 11116 16706 11172 16718
rect 14028 16882 14084 17052
rect 14476 17042 14532 17052
rect 14028 16830 14030 16882
rect 14082 16830 14084 16882
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 13916 14532 13972 14542
rect 14028 14532 14084 16830
rect 16156 16772 16212 18396
rect 15932 16716 16212 16772
rect 14588 15540 14644 15550
rect 13580 14530 14084 14532
rect 13580 14478 13918 14530
rect 13970 14478 14084 14530
rect 13580 14476 14084 14478
rect 14252 15204 14308 15214
rect 13580 13746 13636 14476
rect 13916 14466 13972 14476
rect 14252 13858 14308 15148
rect 14588 14642 14644 15484
rect 15596 15540 15652 15578
rect 15596 15474 15652 15484
rect 15708 15428 15764 15438
rect 15148 15204 15204 15242
rect 15148 15138 15204 15148
rect 15260 15202 15316 15214
rect 15260 15150 15262 15202
rect 15314 15150 15316 15202
rect 14588 14590 14590 14642
rect 14642 14590 14644 14642
rect 14588 14578 14644 14590
rect 14252 13806 14254 13858
rect 14306 13806 14308 13858
rect 14252 13794 14308 13806
rect 13580 13694 13582 13746
rect 13634 13694 13636 13746
rect 13580 13682 13636 13694
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 15260 12628 15316 15150
rect 15708 12852 15764 15372
rect 15820 15316 15876 15326
rect 15932 15316 15988 16716
rect 16380 15428 16436 19292
rect 16604 19122 16660 21196
rect 16940 19236 16996 24556
rect 17724 23378 17780 24780
rect 18172 24612 18228 24622
rect 18172 24518 18228 24556
rect 17724 23326 17726 23378
rect 17778 23326 17780 23378
rect 17724 23314 17780 23326
rect 18060 23714 18116 23726
rect 18060 23662 18062 23714
rect 18114 23662 18116 23714
rect 17276 23156 17332 23166
rect 17276 22820 17332 23100
rect 17164 22596 17220 22606
rect 17164 22258 17220 22540
rect 17276 22594 17332 22764
rect 17612 23154 17668 23166
rect 17612 23102 17614 23154
rect 17666 23102 17668 23154
rect 17612 22708 17668 23102
rect 17612 22642 17668 22652
rect 17836 23154 17892 23166
rect 17836 23102 17838 23154
rect 17890 23102 17892 23154
rect 17276 22542 17278 22594
rect 17330 22542 17332 22594
rect 17276 22530 17332 22542
rect 17836 22596 17892 23102
rect 17836 22530 17892 22540
rect 17836 22372 17892 22382
rect 18060 22372 18116 23662
rect 18396 23716 18452 25342
rect 18396 23622 18452 23660
rect 18732 23940 18788 25452
rect 18844 25506 18900 25518
rect 18844 25454 18846 25506
rect 18898 25454 18900 25506
rect 18844 24164 18900 25454
rect 18844 24098 18900 24108
rect 18956 25508 19012 25518
rect 18956 23940 19012 25452
rect 19404 25508 19460 25518
rect 19516 25508 19572 26796
rect 19740 26786 19796 26796
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 19404 25506 19572 25508
rect 19404 25454 19406 25506
rect 19458 25454 19572 25506
rect 19404 25452 19572 25454
rect 19628 26178 19684 26190
rect 19628 26126 19630 26178
rect 19682 26126 19684 26178
rect 19404 25442 19460 25452
rect 19404 24724 19460 24734
rect 19404 24630 19460 24668
rect 19628 24612 19684 26126
rect 20188 25508 20244 26910
rect 20524 26962 20580 28588
rect 20860 27972 20916 27982
rect 20860 27878 20916 27916
rect 20524 26910 20526 26962
rect 20578 26910 20580 26962
rect 20524 26898 20580 26910
rect 20748 26962 20804 26974
rect 20748 26910 20750 26962
rect 20802 26910 20804 26962
rect 20188 25442 20244 25452
rect 20748 25284 20804 26910
rect 21308 26964 21364 26974
rect 21308 26870 21364 26908
rect 20748 25218 20804 25228
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 20076 24612 20132 24622
rect 19628 24546 19684 24556
rect 19852 24610 20132 24612
rect 19852 24558 20078 24610
rect 20130 24558 20132 24610
rect 19852 24556 20132 24558
rect 18732 23714 18788 23884
rect 18732 23662 18734 23714
rect 18786 23662 18788 23714
rect 18732 23604 18788 23662
rect 18732 23538 18788 23548
rect 18844 23884 19012 23940
rect 19628 24052 19684 24062
rect 18396 23380 18452 23390
rect 18396 23286 18452 23324
rect 18732 23380 18788 23390
rect 18620 23268 18676 23278
rect 18620 23174 18676 23212
rect 18284 23154 18340 23166
rect 18284 23102 18286 23154
rect 18338 23102 18340 23154
rect 17164 22206 17166 22258
rect 17218 22206 17220 22258
rect 17164 19908 17220 22206
rect 17276 22370 18228 22372
rect 17276 22318 17838 22370
rect 17890 22318 18228 22370
rect 17276 22316 18228 22318
rect 17276 22258 17332 22316
rect 17836 22306 17892 22316
rect 17276 22206 17278 22258
rect 17330 22206 17332 22258
rect 17276 22194 17332 22206
rect 17948 22148 18004 22158
rect 17948 21810 18004 22092
rect 18060 22146 18116 22158
rect 18060 22094 18062 22146
rect 18114 22094 18116 22146
rect 18060 22036 18116 22094
rect 18060 21970 18116 21980
rect 17948 21758 17950 21810
rect 18002 21758 18004 21810
rect 17948 21746 18004 21758
rect 17724 21588 17780 21598
rect 17612 21586 17780 21588
rect 17612 21534 17726 21586
rect 17778 21534 17780 21586
rect 17612 21532 17780 21534
rect 17612 20132 17668 21532
rect 17724 21522 17780 21532
rect 18060 21364 18116 21374
rect 18060 21270 18116 21308
rect 17612 20066 17668 20076
rect 17836 20690 17892 20702
rect 17836 20638 17838 20690
rect 17890 20638 17892 20690
rect 17164 19842 17220 19852
rect 16940 19170 16996 19180
rect 17612 19796 17668 19806
rect 17612 19234 17668 19740
rect 17612 19182 17614 19234
rect 17666 19182 17668 19234
rect 17612 19170 17668 19182
rect 17836 19236 17892 20638
rect 17948 20130 18004 20142
rect 17948 20078 17950 20130
rect 18002 20078 18004 20130
rect 17948 19908 18004 20078
rect 17948 19842 18004 19852
rect 16604 19070 16606 19122
rect 16658 19070 16660 19122
rect 16604 19058 16660 19070
rect 17276 19124 17332 19134
rect 17276 19030 17332 19068
rect 16940 19012 16996 19022
rect 16940 18918 16996 18956
rect 17724 18564 17780 18574
rect 16492 18450 16548 18462
rect 17724 18452 17780 18508
rect 16492 18398 16494 18450
rect 16546 18398 16548 18450
rect 16492 18004 16548 18398
rect 16492 17938 16548 17948
rect 17388 18450 17780 18452
rect 17388 18398 17726 18450
rect 17778 18398 17780 18450
rect 17388 18396 17780 18398
rect 17388 17778 17444 18396
rect 17724 18386 17780 18396
rect 17388 17726 17390 17778
rect 17442 17726 17444 17778
rect 17388 17714 17444 17726
rect 16380 15334 16436 15372
rect 17836 17442 17892 19180
rect 17948 18676 18004 18686
rect 18172 18676 18228 22316
rect 18284 21476 18340 23102
rect 18732 23044 18788 23324
rect 18620 22708 18676 22718
rect 18396 22148 18452 22158
rect 18396 22054 18452 22092
rect 18508 21476 18564 21486
rect 18284 21420 18508 21476
rect 18508 21382 18564 21420
rect 18620 20244 18676 22652
rect 18732 22258 18788 22988
rect 18732 22206 18734 22258
rect 18786 22206 18788 22258
rect 18732 22194 18788 22206
rect 18844 22148 18900 23884
rect 19292 23828 19348 23838
rect 19180 23772 19292 23828
rect 19068 23714 19124 23726
rect 19068 23662 19070 23714
rect 19122 23662 19124 23714
rect 19068 23492 19124 23662
rect 19068 23426 19124 23436
rect 18956 23154 19012 23166
rect 18956 23102 18958 23154
rect 19010 23102 19012 23154
rect 18956 22484 19012 23102
rect 19068 22484 19124 22494
rect 18956 22428 19068 22484
rect 19068 22370 19124 22428
rect 19068 22318 19070 22370
rect 19122 22318 19124 22370
rect 19068 22306 19124 22318
rect 18844 22092 19124 22148
rect 18508 20188 18676 20244
rect 18956 21586 19012 21598
rect 18956 21534 18958 21586
rect 19010 21534 19012 21586
rect 18956 21364 19012 21534
rect 18284 20018 18340 20030
rect 18284 19966 18286 20018
rect 18338 19966 18340 20018
rect 18284 19908 18340 19966
rect 18396 19908 18452 19918
rect 18284 19852 18396 19908
rect 18396 19842 18452 19852
rect 17948 18674 18228 18676
rect 17948 18622 17950 18674
rect 18002 18622 18228 18674
rect 17948 18620 18228 18622
rect 17948 18610 18004 18620
rect 18172 18452 18228 18620
rect 18396 19012 18452 19022
rect 18284 18452 18340 18462
rect 18172 18450 18340 18452
rect 18172 18398 18286 18450
rect 18338 18398 18340 18450
rect 18172 18396 18340 18398
rect 18396 18452 18452 18956
rect 18508 18676 18564 20188
rect 18732 20132 18788 20142
rect 18732 20038 18788 20076
rect 18620 20020 18676 20030
rect 18620 19460 18676 19964
rect 18732 19460 18788 19470
rect 18620 19458 18788 19460
rect 18620 19406 18734 19458
rect 18786 19406 18788 19458
rect 18620 19404 18788 19406
rect 18620 19236 18676 19246
rect 18620 19142 18676 19180
rect 18508 18620 18676 18676
rect 18508 18452 18564 18462
rect 18396 18450 18564 18452
rect 18396 18398 18510 18450
rect 18562 18398 18564 18450
rect 18396 18396 18564 18398
rect 18284 18386 18340 18396
rect 18508 18386 18564 18396
rect 17836 17390 17838 17442
rect 17890 17390 17892 17442
rect 15820 15314 15988 15316
rect 15820 15262 15822 15314
rect 15874 15262 15988 15314
rect 15820 15260 15988 15262
rect 16156 15316 16212 15326
rect 16156 15314 16324 15316
rect 16156 15262 16158 15314
rect 16210 15262 16324 15314
rect 16156 15260 16324 15262
rect 15820 12962 15876 15260
rect 16156 15250 16212 15260
rect 15932 15092 15988 15102
rect 15932 14998 15988 15036
rect 16268 14420 16324 15260
rect 16716 14644 16772 14654
rect 16716 14642 16884 14644
rect 16716 14590 16718 14642
rect 16770 14590 16884 14642
rect 16716 14588 16884 14590
rect 16716 14578 16772 14588
rect 16268 14364 16772 14420
rect 16716 13970 16772 14364
rect 16716 13918 16718 13970
rect 16770 13918 16772 13970
rect 16716 13906 16772 13918
rect 16380 13634 16436 13646
rect 16380 13582 16382 13634
rect 16434 13582 16436 13634
rect 16380 13188 16436 13582
rect 16828 13634 16884 14588
rect 17836 14530 17892 17390
rect 18620 17108 18676 18620
rect 18732 17666 18788 19404
rect 18956 19236 19012 21308
rect 19068 19346 19124 22092
rect 19068 19294 19070 19346
rect 19122 19294 19124 19346
rect 19068 19282 19124 19294
rect 19180 19348 19236 23772
rect 19292 23762 19348 23772
rect 19404 23492 19460 23502
rect 19404 23154 19460 23436
rect 19628 23380 19684 23996
rect 19852 24050 19908 24556
rect 20076 24546 20132 24556
rect 21532 24612 21588 37998
rect 21980 38052 22036 38062
rect 21980 28756 22036 37996
rect 24556 38052 24612 38062
rect 24556 37958 24612 37996
rect 24892 37492 24948 41200
rect 26908 38610 26964 41200
rect 26908 38558 26910 38610
rect 26962 38558 26964 38610
rect 26908 38546 26964 38558
rect 27468 38610 27524 38622
rect 27468 38558 27470 38610
rect 27522 38558 27524 38610
rect 25564 38276 25620 38286
rect 25564 38182 25620 38220
rect 27468 37938 27524 38558
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 27468 37886 27470 37938
rect 27522 37886 27524 37938
rect 27468 37874 27524 37886
rect 24892 37426 24948 37436
rect 26236 37492 26292 37502
rect 26236 37398 26292 37436
rect 25228 37266 25284 37278
rect 25228 37214 25230 37266
rect 25282 37214 25284 37266
rect 21980 28754 23044 28756
rect 21980 28702 21982 28754
rect 22034 28702 23044 28754
rect 21980 28700 23044 28702
rect 21980 28690 22036 28700
rect 21868 28644 21924 28654
rect 21868 28550 21924 28588
rect 21756 27860 21812 27870
rect 21644 27524 21700 27534
rect 21644 27298 21700 27468
rect 21644 27246 21646 27298
rect 21698 27246 21700 27298
rect 21644 27234 21700 27246
rect 21756 26908 21812 27804
rect 22988 27746 23044 28700
rect 23548 27860 23604 27870
rect 23548 27766 23604 27804
rect 22988 27694 22990 27746
rect 23042 27694 23044 27746
rect 22988 27682 23044 27694
rect 21868 27076 21924 27114
rect 21868 27010 21924 27020
rect 22652 27076 22708 27086
rect 22708 27020 22820 27076
rect 22652 27010 22708 27020
rect 21756 26852 21924 26908
rect 21868 26290 21924 26852
rect 21868 26238 21870 26290
rect 21922 26238 21924 26290
rect 21868 24724 21924 26238
rect 22540 26178 22596 26190
rect 22540 26126 22542 26178
rect 22594 26126 22596 26178
rect 21868 24658 21924 24668
rect 21980 25284 22036 25294
rect 21588 24556 21812 24612
rect 21532 24546 21588 24556
rect 21532 24276 21588 24286
rect 21420 24052 21476 24062
rect 19852 23998 19854 24050
rect 19906 23998 19908 24050
rect 19852 23986 19908 23998
rect 20412 24050 21476 24052
rect 20412 23998 21422 24050
rect 21474 23998 21476 24050
rect 20412 23996 21476 23998
rect 19964 23938 20020 23950
rect 19964 23886 19966 23938
rect 20018 23886 20020 23938
rect 19740 23828 19796 23838
rect 19740 23734 19796 23772
rect 19964 23716 20020 23886
rect 20188 23940 20244 23950
rect 20188 23846 20244 23884
rect 20412 23938 20468 23996
rect 21420 23986 21476 23996
rect 21532 24052 21588 24220
rect 20412 23886 20414 23938
rect 20466 23886 20468 23938
rect 20412 23874 20468 23886
rect 21532 23938 21588 23996
rect 21532 23886 21534 23938
rect 21586 23886 21588 23938
rect 21532 23874 21588 23886
rect 20636 23828 20692 23838
rect 20524 23826 20692 23828
rect 20524 23774 20638 23826
rect 20690 23774 20692 23826
rect 20524 23772 20692 23774
rect 19964 23660 20244 23716
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 19628 23324 19796 23380
rect 19404 23102 19406 23154
rect 19458 23102 19460 23154
rect 19292 22596 19348 22606
rect 19292 22370 19348 22540
rect 19292 22318 19294 22370
rect 19346 22318 19348 22370
rect 19292 22306 19348 22318
rect 19292 22148 19348 22158
rect 19404 22148 19460 23102
rect 19348 22092 19460 22148
rect 19516 23268 19572 23278
rect 19516 22258 19572 23212
rect 19628 22596 19684 22606
rect 19628 22502 19684 22540
rect 19740 22372 19796 23324
rect 19852 23156 19908 23166
rect 19852 23062 19908 23100
rect 20188 23156 20244 23660
rect 20188 23090 20244 23100
rect 20188 22708 20244 22718
rect 19516 22206 19518 22258
rect 19570 22206 19572 22258
rect 19292 22082 19348 22092
rect 19516 22036 19572 22206
rect 19516 21970 19572 21980
rect 19628 22316 19796 22372
rect 20076 22372 20132 22382
rect 20188 22372 20244 22652
rect 20412 22596 20468 22606
rect 20524 22596 20580 23772
rect 20636 23762 20692 23772
rect 21308 23826 21364 23838
rect 21308 23774 21310 23826
rect 21362 23774 21364 23826
rect 21308 23380 21364 23774
rect 21756 23826 21812 24556
rect 21980 24500 22036 25228
rect 22204 24612 22260 24622
rect 22204 24518 22260 24556
rect 21756 23774 21758 23826
rect 21810 23774 21812 23826
rect 21756 23762 21812 23774
rect 21868 24444 22036 24500
rect 20636 23268 20692 23278
rect 20636 23266 20804 23268
rect 20636 23214 20638 23266
rect 20690 23214 20804 23266
rect 20636 23212 20804 23214
rect 20636 23202 20692 23212
rect 20412 22594 20580 22596
rect 20412 22542 20414 22594
rect 20466 22542 20580 22594
rect 20412 22540 20580 22542
rect 20748 23156 20804 23212
rect 20412 22530 20468 22540
rect 20076 22370 20244 22372
rect 20076 22318 20078 22370
rect 20130 22318 20244 22370
rect 20076 22316 20244 22318
rect 19292 21588 19348 21598
rect 19292 21494 19348 21532
rect 19628 21364 19684 22316
rect 20076 22306 20132 22316
rect 19852 22260 19908 22270
rect 19852 22166 19908 22204
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 19180 19282 19236 19292
rect 19292 21308 19684 21364
rect 19292 19906 19348 21308
rect 20076 20804 20132 20814
rect 20076 20710 20132 20748
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 20188 20242 20244 22316
rect 20188 20190 20190 20242
rect 20242 20190 20244 20242
rect 20188 20178 20244 20190
rect 20524 22372 20580 22382
rect 19292 19854 19294 19906
rect 19346 19854 19348 19906
rect 18956 19170 19012 19180
rect 18844 18228 18900 18238
rect 18844 18226 19236 18228
rect 18844 18174 18846 18226
rect 18898 18174 19236 18226
rect 18844 18172 19236 18174
rect 18844 18162 18900 18172
rect 18732 17614 18734 17666
rect 18786 17614 18788 17666
rect 18732 17602 18788 17614
rect 19068 17444 19124 17454
rect 18844 17442 19124 17444
rect 18844 17390 19070 17442
rect 19122 17390 19124 17442
rect 18844 17388 19124 17390
rect 18732 17108 18788 17118
rect 18620 17106 18788 17108
rect 18620 17054 18734 17106
rect 18786 17054 18788 17106
rect 18620 17052 18788 17054
rect 18284 16100 18340 16110
rect 18284 15986 18340 16044
rect 18508 16100 18564 16110
rect 18620 16100 18676 17052
rect 18732 17042 18788 17052
rect 18508 16098 18676 16100
rect 18508 16046 18510 16098
rect 18562 16046 18676 16098
rect 18508 16044 18676 16046
rect 18732 16100 18788 16110
rect 18844 16100 18900 17388
rect 19068 17378 19124 17388
rect 19068 16884 19124 16894
rect 19068 16790 19124 16828
rect 18732 16098 18900 16100
rect 18732 16046 18734 16098
rect 18786 16046 18900 16098
rect 18732 16044 18900 16046
rect 18508 16034 18564 16044
rect 18732 16034 18788 16044
rect 18284 15934 18286 15986
rect 18338 15934 18340 15986
rect 18284 15922 18340 15934
rect 18844 15988 18900 16044
rect 19068 16100 19124 16110
rect 19180 16100 19236 18172
rect 19124 16044 19236 16100
rect 19292 16098 19348 19854
rect 19404 20132 19460 20142
rect 19404 19234 19460 20076
rect 19852 20132 19908 20142
rect 19852 20038 19908 20076
rect 20524 20130 20580 22316
rect 20524 20078 20526 20130
rect 20578 20078 20580 20130
rect 19628 20018 19684 20030
rect 19628 19966 19630 20018
rect 19682 19966 19684 20018
rect 19404 19182 19406 19234
rect 19458 19182 19460 19234
rect 19404 19170 19460 19182
rect 19516 19346 19572 19358
rect 19516 19294 19518 19346
rect 19570 19294 19572 19346
rect 19516 18676 19572 19294
rect 19404 18338 19460 18350
rect 19404 18286 19406 18338
rect 19458 18286 19460 18338
rect 19404 16884 19460 18286
rect 19404 16818 19460 16828
rect 19292 16046 19294 16098
rect 19346 16046 19348 16098
rect 19068 16006 19124 16044
rect 19292 16034 19348 16046
rect 19516 16098 19572 18620
rect 19628 19236 19684 19966
rect 19628 17556 19684 19180
rect 20188 19908 20244 19918
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 19740 18452 19796 18462
rect 20188 18452 20244 19852
rect 20524 19908 20580 20078
rect 20524 19842 20580 19852
rect 19740 18450 20356 18452
rect 19740 18398 19742 18450
rect 19794 18398 20356 18450
rect 19740 18396 20356 18398
rect 19740 18386 19796 18396
rect 19964 18226 20020 18238
rect 19964 18174 19966 18226
rect 20018 18174 20020 18226
rect 19964 18116 20020 18174
rect 20076 18116 20132 18126
rect 19964 18060 20076 18116
rect 20076 18050 20132 18060
rect 20300 17780 20356 18396
rect 20412 18450 20468 18462
rect 20412 18398 20414 18450
rect 20466 18398 20468 18450
rect 20412 18228 20468 18398
rect 20412 18116 20468 18172
rect 20748 18116 20804 23100
rect 20860 23154 20916 23166
rect 20860 23102 20862 23154
rect 20914 23102 20916 23154
rect 20860 21476 20916 23102
rect 21308 22708 21364 23324
rect 21308 22642 21364 22652
rect 21868 22482 21924 24444
rect 22092 24164 22148 24174
rect 21980 23380 22036 23390
rect 21980 23286 22036 23324
rect 22092 23378 22148 24108
rect 22204 23826 22260 23838
rect 22204 23774 22206 23826
rect 22258 23774 22260 23826
rect 22204 23548 22260 23774
rect 22316 23714 22372 23726
rect 22316 23662 22318 23714
rect 22370 23662 22372 23714
rect 22316 23548 22372 23662
rect 22540 23604 22596 26126
rect 22652 24724 22708 24734
rect 22652 24630 22708 24668
rect 22652 24164 22708 24174
rect 22652 23938 22708 24108
rect 22652 23886 22654 23938
rect 22706 23886 22708 23938
rect 22652 23874 22708 23886
rect 22316 23492 22484 23548
rect 22540 23538 22596 23548
rect 22204 23482 22260 23492
rect 22428 23426 22484 23436
rect 22764 23492 22820 27020
rect 25228 26908 25284 37214
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 24668 26852 25284 26908
rect 24668 26178 24724 26852
rect 24668 26126 24670 26178
rect 24722 26126 24724 26178
rect 23660 25956 23716 25966
rect 23660 24946 23716 25900
rect 24668 25956 24724 26126
rect 24668 25890 24724 25900
rect 25340 26178 25396 26190
rect 25340 26126 25342 26178
rect 25394 26126 25396 26178
rect 23660 24894 23662 24946
rect 23714 24894 23716 24946
rect 23660 24882 23716 24894
rect 23100 24722 23156 24734
rect 23100 24670 23102 24722
rect 23154 24670 23156 24722
rect 22988 24052 23044 24062
rect 22988 23958 23044 23996
rect 22988 23604 23044 23614
rect 22764 23426 22820 23436
rect 22876 23492 23044 23548
rect 22092 23326 22094 23378
rect 22146 23326 22148 23378
rect 22092 23314 22148 23326
rect 22876 23378 22932 23492
rect 23100 23380 23156 24670
rect 23436 24722 23492 24734
rect 23436 24670 23438 24722
rect 23490 24670 23492 24722
rect 23436 24276 23492 24670
rect 23772 24724 23828 24734
rect 23436 24210 23492 24220
rect 23548 24610 23604 24622
rect 23548 24558 23550 24610
rect 23602 24558 23604 24610
rect 23212 23826 23268 23838
rect 23212 23774 23214 23826
rect 23266 23774 23268 23826
rect 23212 23716 23268 23774
rect 23324 23828 23380 23838
rect 23324 23734 23380 23772
rect 23436 23826 23492 23838
rect 23436 23774 23438 23826
rect 23490 23774 23492 23826
rect 23212 23650 23268 23660
rect 22876 23326 22878 23378
rect 22930 23326 22932 23378
rect 22876 23314 22932 23326
rect 22988 23324 23156 23380
rect 22428 23268 22484 23278
rect 22204 23156 22260 23166
rect 22428 23156 22484 23212
rect 22204 23154 22484 23156
rect 22204 23102 22206 23154
rect 22258 23102 22484 23154
rect 22204 23100 22484 23102
rect 22652 23156 22708 23166
rect 22876 23156 22932 23166
rect 22652 23154 22820 23156
rect 22652 23102 22654 23154
rect 22706 23102 22820 23154
rect 22652 23100 22820 23102
rect 22204 23090 22260 23100
rect 22652 23090 22708 23100
rect 21868 22430 21870 22482
rect 21922 22430 21924 22482
rect 21868 22418 21924 22430
rect 21308 22372 21364 22382
rect 21308 22278 21364 22316
rect 21980 22372 22036 22382
rect 20860 20692 20916 21420
rect 20860 20626 20916 20636
rect 21420 22260 21476 22270
rect 21308 20132 21364 20142
rect 21308 19346 21364 20076
rect 21420 20020 21476 22204
rect 21868 20804 21924 20814
rect 21980 20804 22036 22316
rect 22204 22260 22260 22270
rect 21868 20802 22036 20804
rect 21868 20750 21870 20802
rect 21922 20750 22036 20802
rect 21868 20748 22036 20750
rect 21868 20738 21924 20748
rect 21644 20692 21700 20702
rect 21644 20598 21700 20636
rect 21532 20020 21588 20030
rect 21420 20018 21588 20020
rect 21420 19966 21534 20018
rect 21586 19966 21588 20018
rect 21420 19964 21588 19966
rect 21420 19796 21476 19964
rect 21532 19954 21588 19964
rect 21980 19796 22036 20748
rect 22092 21252 22148 21262
rect 22092 20690 22148 21196
rect 22204 21026 22260 22204
rect 22204 20974 22206 21026
rect 22258 20974 22260 21026
rect 22204 20962 22260 20974
rect 22092 20638 22094 20690
rect 22146 20638 22148 20690
rect 22092 20626 22148 20638
rect 22428 20130 22484 20142
rect 22428 20078 22430 20130
rect 22482 20078 22484 20130
rect 22092 20020 22148 20030
rect 22428 20020 22484 20078
rect 22092 20018 22484 20020
rect 22092 19966 22094 20018
rect 22146 19966 22484 20018
rect 22092 19964 22484 19966
rect 22092 19954 22148 19964
rect 21980 19740 22148 19796
rect 21420 19730 21476 19740
rect 21308 19294 21310 19346
rect 21362 19294 21364 19346
rect 21308 19282 21364 19294
rect 21756 19234 21812 19246
rect 21756 19182 21758 19234
rect 21810 19182 21812 19234
rect 21420 18676 21476 18714
rect 21420 18610 21476 18620
rect 20860 18564 20916 18574
rect 20860 18470 20916 18508
rect 20412 18060 20692 18116
rect 20412 17780 20468 17790
rect 20300 17778 20468 17780
rect 20300 17726 20414 17778
rect 20466 17726 20468 17778
rect 20300 17724 20468 17726
rect 20412 17714 20468 17724
rect 20636 17666 20692 18060
rect 20748 18050 20804 18060
rect 21420 18450 21476 18462
rect 21420 18398 21422 18450
rect 21474 18398 21476 18450
rect 21420 18340 21476 18398
rect 20636 17614 20638 17666
rect 20690 17614 20692 17666
rect 20636 17602 20692 17614
rect 19740 17556 19796 17566
rect 19628 17554 19796 17556
rect 19628 17502 19742 17554
rect 19794 17502 19796 17554
rect 19628 17500 19796 17502
rect 19740 17490 19796 17500
rect 20076 17444 20132 17482
rect 20076 17378 20132 17388
rect 21084 17444 21140 17454
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 21084 17108 21140 17388
rect 20748 17106 21140 17108
rect 20748 17054 21086 17106
rect 21138 17054 21140 17106
rect 20748 17052 21140 17054
rect 19964 16884 20020 16894
rect 19964 16210 20020 16828
rect 19964 16158 19966 16210
rect 20018 16158 20020 16210
rect 19964 16146 20020 16158
rect 19516 16046 19518 16098
rect 19570 16046 19572 16098
rect 18844 15922 18900 15932
rect 18620 15874 18676 15886
rect 18620 15822 18622 15874
rect 18674 15822 18676 15874
rect 18620 15540 18676 15822
rect 17836 14478 17838 14530
rect 17890 14478 17892 14530
rect 16828 13582 16830 13634
rect 16882 13582 16884 13634
rect 15820 12910 15822 12962
rect 15874 12910 15876 12962
rect 15820 12898 15876 12910
rect 15932 13132 16436 13188
rect 16604 13524 16660 13534
rect 15932 12964 15988 13132
rect 15932 12908 16100 12964
rect 15708 12786 15764 12796
rect 15932 12738 15988 12750
rect 15932 12686 15934 12738
rect 15986 12686 15988 12738
rect 15932 12628 15988 12686
rect 15260 12572 15988 12628
rect 16044 12738 16100 12908
rect 16604 12962 16660 13468
rect 16604 12910 16606 12962
rect 16658 12910 16660 12962
rect 16604 12898 16660 12910
rect 16156 12852 16212 12862
rect 16156 12758 16212 12796
rect 16044 12686 16046 12738
rect 16098 12686 16100 12738
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 16044 11620 16100 12686
rect 16044 11554 16100 11564
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 16828 8428 16884 13582
rect 17500 14308 17556 14318
rect 17836 14308 17892 14478
rect 18508 15484 18676 15540
rect 19180 15874 19236 15886
rect 19180 15822 19182 15874
rect 19234 15822 19236 15874
rect 18508 14420 18564 15484
rect 19180 15092 19236 15822
rect 19516 15204 19572 16046
rect 20188 16100 20244 16110
rect 20188 16006 20244 16044
rect 20524 15874 20580 15886
rect 20524 15822 20526 15874
rect 20578 15822 20580 15874
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 19516 15138 19572 15148
rect 20524 15540 20580 15822
rect 18620 15036 19236 15092
rect 18620 14642 18676 15036
rect 20524 14868 20580 15484
rect 18620 14590 18622 14642
rect 18674 14590 18676 14642
rect 18620 14578 18676 14590
rect 20188 14812 20580 14868
rect 18508 14364 19460 14420
rect 17500 14306 17892 14308
rect 17500 14254 17502 14306
rect 17554 14254 17892 14306
rect 17500 14252 17892 14254
rect 17500 13634 17556 14252
rect 19404 13746 19460 14364
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 19404 13694 19406 13746
rect 19458 13694 19460 13746
rect 19404 13682 19460 13694
rect 17500 13582 17502 13634
rect 17554 13582 17556 13634
rect 17164 13076 17220 13086
rect 17500 13076 17556 13582
rect 19180 13634 19236 13646
rect 19180 13582 19182 13634
rect 19234 13582 19236 13634
rect 19180 13524 19236 13582
rect 19180 13458 19236 13468
rect 19740 13524 19796 13534
rect 20188 13524 20244 14812
rect 20748 14642 20804 17052
rect 21084 17042 21140 17052
rect 21420 17106 21476 18284
rect 21756 18452 21812 19182
rect 22092 18788 22148 19740
rect 22428 19460 22484 19964
rect 22428 19394 22484 19404
rect 22540 20132 22596 20142
rect 22204 19348 22260 19358
rect 22204 19122 22260 19292
rect 22540 19234 22596 20076
rect 22540 19182 22542 19234
rect 22594 19182 22596 19234
rect 22540 19170 22596 19182
rect 22652 20018 22708 20030
rect 22652 19966 22654 20018
rect 22706 19966 22708 20018
rect 22204 19070 22206 19122
rect 22258 19070 22260 19122
rect 22204 19058 22260 19070
rect 22428 19124 22484 19134
rect 22092 18732 22260 18788
rect 21980 18452 22036 18462
rect 21756 18450 22036 18452
rect 21756 18398 21982 18450
rect 22034 18398 22036 18450
rect 21756 18396 22036 18398
rect 21756 17666 21812 18396
rect 21980 18386 22036 18396
rect 22092 18452 22148 18462
rect 22092 18358 22148 18396
rect 22204 18004 22260 18732
rect 22428 18564 22484 19068
rect 22652 19012 22708 19966
rect 22764 19796 22820 23100
rect 22876 23062 22932 23100
rect 22876 22708 22932 22718
rect 22988 22708 23044 23324
rect 22932 22652 23044 22708
rect 23100 23154 23156 23166
rect 23100 23102 23102 23154
rect 23154 23102 23156 23154
rect 23100 23044 23156 23102
rect 22876 22642 22932 22652
rect 23100 22260 23156 22988
rect 23324 23154 23380 23166
rect 23324 23102 23326 23154
rect 23378 23102 23380 23154
rect 23324 22932 23380 23102
rect 23436 23044 23492 23774
rect 23548 23266 23604 24558
rect 23772 23938 23828 24668
rect 25340 24724 25396 26126
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 27580 24948 27636 24958
rect 26796 24834 26852 24846
rect 26796 24782 26798 24834
rect 26850 24782 26852 24834
rect 25340 24658 25396 24668
rect 26460 24724 26516 24734
rect 26516 24668 26628 24724
rect 26460 24630 26516 24668
rect 23772 23886 23774 23938
rect 23826 23886 23828 23938
rect 23772 23874 23828 23886
rect 24556 23828 24612 23838
rect 24556 23734 24612 23772
rect 25452 23716 25508 23726
rect 25452 23378 25508 23660
rect 25452 23326 25454 23378
rect 25506 23326 25508 23378
rect 25452 23314 25508 23326
rect 26348 23604 26404 23614
rect 26348 23378 26404 23548
rect 26348 23326 26350 23378
rect 26402 23326 26404 23378
rect 26348 23314 26404 23326
rect 23548 23214 23550 23266
rect 23602 23214 23604 23266
rect 23548 23202 23604 23214
rect 24332 23268 24388 23278
rect 24332 23174 24388 23212
rect 26460 23268 26516 23278
rect 26460 23174 26516 23212
rect 23772 23154 23828 23166
rect 23772 23102 23774 23154
rect 23826 23102 23828 23154
rect 23772 23044 23828 23102
rect 23436 22988 23828 23044
rect 23324 22866 23380 22876
rect 23772 22484 23828 22988
rect 23436 22372 23492 22382
rect 23436 22278 23492 22316
rect 23100 22194 23156 22204
rect 22876 21474 22932 21486
rect 22876 21422 22878 21474
rect 22930 21422 22932 21474
rect 22876 20804 22932 21422
rect 22876 20710 22932 20748
rect 23548 20244 23604 20254
rect 23772 20244 23828 22428
rect 24108 23154 24164 23166
rect 24108 23102 24110 23154
rect 24162 23102 24164 23154
rect 24108 21252 24164 23102
rect 25116 23156 25172 23166
rect 24444 22932 24500 22942
rect 24444 22148 24500 22876
rect 25116 22260 25172 23100
rect 26124 23156 26180 23166
rect 26572 23156 26628 24668
rect 26796 24276 26852 24782
rect 27580 24836 27636 24892
rect 27692 24836 27748 24846
rect 27580 24834 27748 24836
rect 27580 24782 27694 24834
rect 27746 24782 27748 24834
rect 27580 24780 27748 24782
rect 27692 24770 27748 24780
rect 26796 24210 26852 24220
rect 27020 24722 27076 24734
rect 27020 24670 27022 24722
rect 27074 24670 27076 24722
rect 26684 24052 26740 24062
rect 26684 23958 26740 23996
rect 27020 23826 27076 24670
rect 27356 24724 27412 24734
rect 27356 24722 27636 24724
rect 27356 24670 27358 24722
rect 27410 24670 27636 24722
rect 27356 24668 27636 24670
rect 27356 24658 27412 24668
rect 27132 24500 27188 24510
rect 27132 24498 27524 24500
rect 27132 24446 27134 24498
rect 27186 24446 27524 24498
rect 27132 24444 27524 24446
rect 27132 24434 27188 24444
rect 27132 24052 27188 24062
rect 27132 23958 27188 23996
rect 27020 23774 27022 23826
rect 27074 23774 27076 23826
rect 26908 23268 26964 23278
rect 26796 23156 26852 23166
rect 26572 23154 26852 23156
rect 26572 23102 26798 23154
rect 26850 23102 26852 23154
rect 26572 23100 26852 23102
rect 26124 23062 26180 23100
rect 25228 23044 25284 23054
rect 25228 22950 25284 22988
rect 25452 23042 25508 23054
rect 25452 22990 25454 23042
rect 25506 22990 25508 23042
rect 24444 22082 24500 22092
rect 25004 22258 25172 22260
rect 25004 22206 25118 22258
rect 25170 22206 25172 22258
rect 25004 22204 25172 22206
rect 24108 21186 24164 21196
rect 23548 20242 23828 20244
rect 23548 20190 23550 20242
rect 23602 20190 23828 20242
rect 23548 20188 23828 20190
rect 23548 20178 23604 20188
rect 24220 20132 24276 20142
rect 24220 20038 24276 20076
rect 25004 20132 25060 22204
rect 25116 22194 25172 22204
rect 25340 21812 25396 21822
rect 25340 21718 25396 21756
rect 25228 21698 25284 21710
rect 25228 21646 25230 21698
rect 25282 21646 25284 21698
rect 25228 21588 25284 21646
rect 25340 21588 25396 21598
rect 25228 21532 25340 21588
rect 25340 21522 25396 21532
rect 25452 20356 25508 22990
rect 25676 23044 25732 23054
rect 25564 21812 25620 21822
rect 25676 21812 25732 22988
rect 26236 22596 26292 22606
rect 25788 22484 25844 22494
rect 25788 22370 25844 22428
rect 25788 22318 25790 22370
rect 25842 22318 25844 22370
rect 25788 22306 25844 22318
rect 25564 21810 25732 21812
rect 25564 21758 25566 21810
rect 25618 21758 25732 21810
rect 25564 21756 25732 21758
rect 25900 21812 25956 21822
rect 25564 21746 25620 21756
rect 25452 20300 25732 20356
rect 25004 20066 25060 20076
rect 25564 20130 25620 20142
rect 25564 20078 25566 20130
rect 25618 20078 25620 20130
rect 22988 20020 23044 20030
rect 23212 20020 23268 20030
rect 22988 20018 23268 20020
rect 22988 19966 22990 20018
rect 23042 19966 23214 20018
rect 23266 19966 23268 20018
rect 22988 19964 23268 19966
rect 22988 19954 23044 19964
rect 22764 19702 22820 19740
rect 23100 19346 23156 19964
rect 23212 19954 23268 19964
rect 23884 20018 23940 20030
rect 23884 19966 23886 20018
rect 23938 19966 23940 20018
rect 23548 19460 23604 19470
rect 23548 19366 23604 19404
rect 23100 19294 23102 19346
rect 23154 19294 23156 19346
rect 23100 19282 23156 19294
rect 22652 18946 22708 18956
rect 22876 19234 22932 19246
rect 22876 19182 22878 19234
rect 22930 19182 22932 19234
rect 22428 18450 22484 18508
rect 22428 18398 22430 18450
rect 22482 18398 22484 18450
rect 22428 18386 22484 18398
rect 22876 18452 22932 19182
rect 22876 18386 22932 18396
rect 23212 19122 23268 19134
rect 23212 19070 23214 19122
rect 23266 19070 23268 19122
rect 23212 18340 23268 19070
rect 23660 19124 23716 19134
rect 23660 19030 23716 19068
rect 23324 18676 23380 18686
rect 23324 18582 23380 18620
rect 23212 18274 23268 18284
rect 23436 18452 23492 18462
rect 22652 18228 22708 18238
rect 22652 18134 22708 18172
rect 22876 18226 22932 18238
rect 22876 18174 22878 18226
rect 22930 18174 22932 18226
rect 22204 17778 22260 17948
rect 22204 17726 22206 17778
rect 22258 17726 22260 17778
rect 22204 17714 22260 17726
rect 21756 17614 21758 17666
rect 21810 17614 21812 17666
rect 21756 17602 21812 17614
rect 22876 17668 22932 18174
rect 23212 17668 23268 17678
rect 22876 17666 23268 17668
rect 22876 17614 23214 17666
rect 23266 17614 23268 17666
rect 22876 17612 23268 17614
rect 21420 17054 21422 17106
rect 21474 17054 21476 17106
rect 21420 17042 21476 17054
rect 22876 16772 22932 16782
rect 22876 15538 22932 16716
rect 22876 15486 22878 15538
rect 22930 15486 22932 15538
rect 22876 15474 22932 15486
rect 23100 15540 23156 15550
rect 23100 15446 23156 15484
rect 22988 15202 23044 15214
rect 22988 15150 22990 15202
rect 23042 15150 23044 15202
rect 20748 14590 20750 14642
rect 20802 14590 20804 14642
rect 20748 14578 20804 14590
rect 22876 14644 22932 14654
rect 22988 14644 23044 15150
rect 22876 14642 23044 14644
rect 22876 14590 22878 14642
rect 22930 14590 23044 14642
rect 22876 14588 23044 14590
rect 22876 14578 22932 14588
rect 22092 14530 22148 14542
rect 22092 14478 22094 14530
rect 22146 14478 22148 14530
rect 20300 13748 20356 13758
rect 20300 13654 20356 13692
rect 22092 13748 22148 14478
rect 22092 13682 22148 13692
rect 20972 13636 21028 13646
rect 19740 13522 20132 13524
rect 19740 13470 19742 13522
rect 19794 13470 20132 13522
rect 19740 13468 20132 13470
rect 19740 13458 19796 13468
rect 17164 13074 17556 13076
rect 17164 13022 17166 13074
rect 17218 13022 17556 13074
rect 17164 13020 17556 13022
rect 17164 13010 17220 13020
rect 20076 12964 20132 13468
rect 20188 13458 20244 13468
rect 20412 13634 21028 13636
rect 20412 13582 20974 13634
rect 21026 13582 21028 13634
rect 20412 13580 21028 13582
rect 20188 12964 20244 12974
rect 20076 12962 20244 12964
rect 20076 12910 20190 12962
rect 20242 12910 20244 12962
rect 20076 12908 20244 12910
rect 20188 12898 20244 12908
rect 20412 12850 20468 13580
rect 20972 13570 21028 13580
rect 23100 13636 23156 13646
rect 23212 13636 23268 17612
rect 23436 17554 23492 18396
rect 23772 18340 23828 18350
rect 23884 18340 23940 19966
rect 25564 19572 25620 20078
rect 25564 19506 25620 19516
rect 25676 19460 25732 20300
rect 25788 20132 25844 20142
rect 25788 20018 25844 20076
rect 25788 19966 25790 20018
rect 25842 19966 25844 20018
rect 25788 19954 25844 19966
rect 25676 19404 25844 19460
rect 25116 19236 25172 19246
rect 25116 18676 25172 19180
rect 25676 19236 25732 19246
rect 25676 19142 25732 19180
rect 25228 19124 25284 19134
rect 25228 18788 25284 19068
rect 25340 19124 25396 19134
rect 25340 19030 25396 19068
rect 25452 19012 25508 19022
rect 25676 19012 25732 19022
rect 25452 19010 25676 19012
rect 25452 18958 25454 19010
rect 25506 18958 25676 19010
rect 25452 18956 25676 18958
rect 25452 18946 25508 18956
rect 25676 18946 25732 18956
rect 25228 18732 25508 18788
rect 25116 18620 25284 18676
rect 24668 18564 24724 18574
rect 23828 18284 23940 18340
rect 23996 18452 24052 18462
rect 23772 18246 23828 18284
rect 23996 17666 24052 18396
rect 24668 18450 24724 18508
rect 25228 18562 25284 18620
rect 25452 18674 25508 18732
rect 25788 18676 25844 19404
rect 25452 18622 25454 18674
rect 25506 18622 25508 18674
rect 25452 18610 25508 18622
rect 25564 18620 25844 18676
rect 25900 19010 25956 21756
rect 26012 21588 26068 21626
rect 26068 21532 26180 21588
rect 26012 21522 26068 21532
rect 25900 18958 25902 19010
rect 25954 18958 25956 19010
rect 25900 18676 25956 18958
rect 25228 18510 25230 18562
rect 25282 18510 25284 18562
rect 25228 18498 25284 18510
rect 25564 18452 25620 18620
rect 25900 18610 25956 18620
rect 26012 21362 26068 21374
rect 26012 21310 26014 21362
rect 26066 21310 26068 21362
rect 24668 18398 24670 18450
rect 24722 18398 24724 18450
rect 24668 18386 24724 18398
rect 25452 18396 25620 18452
rect 25788 18452 25844 18462
rect 26012 18452 26068 21310
rect 26124 18564 26180 21532
rect 26236 21586 26292 22540
rect 26796 22484 26852 23100
rect 26460 22258 26516 22270
rect 26460 22206 26462 22258
rect 26514 22206 26516 22258
rect 26460 21810 26516 22206
rect 26460 21758 26462 21810
rect 26514 21758 26516 21810
rect 26460 21746 26516 21758
rect 26236 21534 26238 21586
rect 26290 21534 26292 21586
rect 26236 21522 26292 21534
rect 26572 21588 26628 21598
rect 26572 21494 26628 21532
rect 26796 20914 26852 22428
rect 26796 20862 26798 20914
rect 26850 20862 26852 20914
rect 26348 20244 26404 20254
rect 26796 20244 26852 20862
rect 26348 20242 26852 20244
rect 26348 20190 26350 20242
rect 26402 20190 26852 20242
rect 26348 20188 26852 20190
rect 26236 19012 26292 19022
rect 26236 18918 26292 18956
rect 26236 18676 26292 18686
rect 26348 18676 26404 20188
rect 26796 20018 26852 20188
rect 26796 19966 26798 20018
rect 26850 19966 26852 20018
rect 26796 19954 26852 19966
rect 26908 21810 26964 23212
rect 27020 23044 27076 23774
rect 27356 23828 27412 23838
rect 27356 23734 27412 23772
rect 27468 23268 27524 24444
rect 27580 24276 27636 24668
rect 37884 24722 37940 24734
rect 37884 24670 37886 24722
rect 37938 24670 37940 24722
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 27580 24220 28084 24276
rect 35196 24266 35460 24276
rect 28028 24162 28084 24220
rect 28028 24110 28030 24162
rect 28082 24110 28084 24162
rect 28028 24098 28084 24110
rect 28028 23940 28084 23950
rect 27580 23826 27636 23838
rect 27580 23774 27582 23826
rect 27634 23774 27636 23826
rect 27580 23604 27636 23774
rect 27580 23538 27636 23548
rect 27916 23826 27972 23838
rect 27916 23774 27918 23826
rect 27970 23774 27972 23826
rect 27580 23268 27636 23278
rect 27468 23266 27636 23268
rect 27468 23214 27582 23266
rect 27634 23214 27636 23266
rect 27468 23212 27636 23214
rect 27580 23202 27636 23212
rect 27916 23268 27972 23774
rect 28028 23826 28084 23884
rect 28028 23774 28030 23826
rect 28082 23774 28084 23826
rect 28028 23762 28084 23774
rect 29708 23940 29764 23950
rect 27916 23202 27972 23212
rect 27020 22978 27076 22988
rect 29708 23042 29764 23884
rect 37660 23940 37716 23950
rect 37660 23846 37716 23884
rect 37884 23828 37940 24670
rect 40012 24498 40068 24510
rect 40012 24446 40014 24498
rect 40066 24446 40068 24498
rect 40012 24276 40068 24446
rect 40012 24210 40068 24220
rect 37884 23762 37940 23772
rect 40012 24050 40068 24062
rect 40012 23998 40014 24050
rect 40066 23998 40068 24050
rect 40012 23604 40068 23998
rect 40012 23538 40068 23548
rect 29708 22990 29710 23042
rect 29762 22990 29764 23042
rect 29708 22978 29764 22990
rect 37660 23154 37716 23166
rect 37660 23102 37662 23154
rect 37714 23102 37716 23154
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 26908 21758 26910 21810
rect 26962 21758 26964 21810
rect 26796 19348 26852 19358
rect 26796 19254 26852 19292
rect 26572 19236 26628 19246
rect 26572 19142 26628 19180
rect 26684 19012 26740 19022
rect 26236 18674 26628 18676
rect 26236 18622 26238 18674
rect 26290 18622 26628 18674
rect 26236 18620 26628 18622
rect 26236 18610 26292 18620
rect 26124 18498 26180 18508
rect 25844 18396 26068 18452
rect 23996 17614 23998 17666
rect 24050 17614 24052 17666
rect 23996 17602 24052 17614
rect 23436 17502 23438 17554
rect 23490 17502 23492 17554
rect 23436 17490 23492 17502
rect 23772 17442 23828 17454
rect 23772 17390 23774 17442
rect 23826 17390 23828 17442
rect 23772 16884 23828 17390
rect 23772 16100 23828 16828
rect 25452 16772 25508 18396
rect 25788 18358 25844 18396
rect 25564 18228 25620 18238
rect 25564 18226 26180 18228
rect 25564 18174 25566 18226
rect 25618 18174 26180 18226
rect 25564 18172 26180 18174
rect 25564 18162 25620 18172
rect 25452 16706 25508 16716
rect 24108 16100 24164 16110
rect 23772 16098 24164 16100
rect 23772 16046 24110 16098
rect 24162 16046 24164 16098
rect 23772 16044 24164 16046
rect 24108 16034 24164 16044
rect 24444 16100 24500 16110
rect 24444 15986 24500 16044
rect 25788 16100 25844 16110
rect 24444 15934 24446 15986
rect 24498 15934 24500 15986
rect 24444 15922 24500 15934
rect 25228 15988 25284 15998
rect 25228 15538 25284 15932
rect 25228 15486 25230 15538
rect 25282 15486 25284 15538
rect 25228 15474 25284 15486
rect 23436 15316 23492 15326
rect 23436 15222 23492 15260
rect 25340 15316 25396 15326
rect 25340 15222 25396 15260
rect 25452 15314 25508 15326
rect 25452 15262 25454 15314
rect 25506 15262 25508 15314
rect 25452 14756 25508 15262
rect 25788 15314 25844 16044
rect 26124 16098 26180 18172
rect 26124 16046 26126 16098
rect 26178 16046 26180 16098
rect 26124 16034 26180 16046
rect 25900 15988 25956 15998
rect 25900 15894 25956 15932
rect 26348 15876 26404 15886
rect 25788 15262 25790 15314
rect 25842 15262 25844 15314
rect 25788 15250 25844 15262
rect 26124 15874 26404 15876
rect 26124 15822 26350 15874
rect 26402 15822 26404 15874
rect 26124 15820 26404 15822
rect 25228 14700 25508 14756
rect 25004 14644 25060 14654
rect 25228 14644 25284 14700
rect 25004 14642 25284 14644
rect 25004 14590 25006 14642
rect 25058 14590 25284 14642
rect 25004 14588 25284 14590
rect 25004 14578 25060 14588
rect 23548 13748 23604 13758
rect 23548 13654 23604 13692
rect 23100 13634 23268 13636
rect 23100 13582 23102 13634
rect 23154 13582 23268 13634
rect 23100 13580 23268 13582
rect 23100 13570 23156 13580
rect 20412 12798 20414 12850
rect 20466 12798 20468 12850
rect 20412 12786 20468 12798
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 17388 11620 17444 11630
rect 16828 8372 17108 8428
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 16156 4228 16212 4238
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 16156 800 16212 4172
rect 17052 3554 17108 8372
rect 17388 4338 17444 11564
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 17388 4286 17390 4338
rect 17442 4286 17444 4338
rect 17388 4274 17444 4286
rect 18508 4228 18564 4238
rect 18508 4134 18564 4172
rect 17052 3502 17054 3554
rect 17106 3502 17108 3554
rect 17052 3490 17108 3502
rect 24892 3668 24948 3678
rect 16828 3444 16884 3454
rect 16828 800 16884 3388
rect 18060 3444 18116 3454
rect 18060 3330 18116 3388
rect 18060 3278 18062 3330
rect 18114 3278 18116 3330
rect 18060 3266 18116 3278
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 24892 800 24948 3612
rect 25228 3554 25284 14588
rect 26124 14642 26180 15820
rect 26348 15810 26404 15820
rect 26460 15652 26516 18620
rect 26572 18450 26628 18620
rect 26684 18564 26740 18956
rect 26908 18676 26964 21758
rect 27356 22596 27412 22606
rect 27356 21810 27412 22540
rect 28588 22596 28644 22606
rect 28588 22482 28644 22540
rect 37660 22596 37716 23102
rect 40012 22932 40068 22942
rect 40012 22838 40068 22876
rect 37660 22530 37716 22540
rect 28588 22430 28590 22482
rect 28642 22430 28644 22482
rect 28588 22418 28644 22430
rect 29260 22484 29316 22494
rect 29260 22390 29316 22428
rect 27356 21758 27358 21810
rect 27410 21758 27412 21810
rect 27356 21746 27412 21758
rect 27804 22148 27860 22158
rect 27020 21588 27076 21598
rect 27020 21494 27076 21532
rect 27132 21586 27188 21598
rect 27132 21534 27134 21586
rect 27186 21534 27188 21586
rect 27132 20804 27188 21534
rect 27132 20738 27188 20748
rect 27468 19906 27524 19918
rect 27468 19854 27470 19906
rect 27522 19854 27524 19906
rect 27020 19796 27076 19806
rect 27020 19234 27076 19740
rect 27468 19348 27524 19854
rect 27468 19282 27524 19292
rect 27020 19182 27022 19234
rect 27074 19182 27076 19234
rect 27020 19170 27076 19182
rect 27132 19234 27188 19246
rect 27132 19182 27134 19234
rect 27186 19182 27188 19234
rect 27132 19124 27188 19182
rect 27804 19234 27860 22092
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 40012 20914 40068 20926
rect 40012 20862 40014 20914
rect 40066 20862 40068 20914
rect 37660 20802 37716 20814
rect 37660 20750 37662 20802
rect 37714 20750 37716 20802
rect 27804 19182 27806 19234
rect 27858 19182 27860 19234
rect 27804 19170 27860 19182
rect 29596 19908 29652 19918
rect 27580 19124 27636 19134
rect 28140 19124 28196 19134
rect 27132 19122 27636 19124
rect 27132 19070 27582 19122
rect 27634 19070 27636 19122
rect 27132 19068 27636 19070
rect 27132 19012 27188 19068
rect 27580 19058 27636 19068
rect 28028 19122 28196 19124
rect 28028 19070 28142 19122
rect 28194 19070 28196 19122
rect 28028 19068 28196 19070
rect 27916 19012 27972 19022
rect 27132 18946 27188 18956
rect 27692 19010 27972 19012
rect 27692 18958 27918 19010
rect 27970 18958 27972 19010
rect 27692 18956 27972 18958
rect 26908 18610 26964 18620
rect 27244 18676 27300 18686
rect 27692 18676 27748 18956
rect 27916 18946 27972 18956
rect 26684 18498 26740 18508
rect 26572 18398 26574 18450
rect 26626 18398 26628 18450
rect 26572 18386 26628 18398
rect 27244 16994 27300 18620
rect 27356 18620 27748 18676
rect 27356 18562 27412 18620
rect 27356 18510 27358 18562
rect 27410 18510 27412 18562
rect 27356 18498 27412 18510
rect 27692 18340 27748 18350
rect 27580 17554 27636 17566
rect 27580 17502 27582 17554
rect 27634 17502 27636 17554
rect 27244 16942 27246 16994
rect 27298 16942 27300 16994
rect 27244 16930 27300 16942
rect 27356 17106 27412 17118
rect 27356 17054 27358 17106
rect 27410 17054 27412 17106
rect 27132 16882 27188 16894
rect 27132 16830 27134 16882
rect 27186 16830 27188 16882
rect 26572 16098 26628 16110
rect 26572 16046 26574 16098
rect 26626 16046 26628 16098
rect 26572 15988 26628 16046
rect 27020 16100 27076 16110
rect 27020 16006 27076 16044
rect 26684 15988 26740 15998
rect 26572 15986 26740 15988
rect 26572 15934 26686 15986
rect 26738 15934 26740 15986
rect 26572 15932 26740 15934
rect 26684 15922 26740 15932
rect 27132 15988 27188 16830
rect 27132 15922 27188 15932
rect 26908 15874 26964 15886
rect 26908 15822 26910 15874
rect 26962 15822 26964 15874
rect 26908 15764 26964 15822
rect 26908 15698 26964 15708
rect 26124 14590 26126 14642
rect 26178 14590 26180 14642
rect 26124 14578 26180 14590
rect 26236 15596 26516 15652
rect 26236 15538 26292 15596
rect 26236 15486 26238 15538
rect 26290 15486 26292 15538
rect 25340 14532 25396 14542
rect 25340 13748 25396 14476
rect 26236 14532 26292 15486
rect 26460 15316 26516 15596
rect 27356 15426 27412 17054
rect 27580 16100 27636 17502
rect 27692 17554 27748 18284
rect 27916 17668 27972 17678
rect 28028 17668 28084 19068
rect 28140 19058 28196 19068
rect 29596 19124 29652 19852
rect 37660 19908 37716 20750
rect 40012 20244 40068 20862
rect 40012 20178 40068 20188
rect 37660 19842 37716 19852
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 29596 19058 29652 19068
rect 37660 18452 37716 18462
rect 37660 18358 37716 18396
rect 29484 18340 29540 18350
rect 29484 18246 29540 18284
rect 40012 18228 40068 18238
rect 40012 18134 40068 18172
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 27916 17666 28084 17668
rect 27916 17614 27918 17666
rect 27970 17614 28084 17666
rect 27916 17612 28084 17614
rect 27916 17602 27972 17612
rect 27692 17502 27694 17554
rect 27746 17502 27748 17554
rect 27692 17490 27748 17502
rect 27692 16882 27748 16894
rect 27692 16830 27694 16882
rect 27746 16830 27748 16882
rect 27692 16322 27748 16830
rect 37884 16882 37940 16894
rect 37884 16830 37886 16882
rect 37938 16830 37940 16882
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 27692 16270 27694 16322
rect 27746 16270 27748 16322
rect 27692 16258 27748 16270
rect 27580 16006 27636 16044
rect 37660 16098 37716 16110
rect 37660 16046 37662 16098
rect 37714 16046 37716 16098
rect 27356 15374 27358 15426
rect 27410 15374 27412 15426
rect 27356 15362 27412 15374
rect 27692 15874 27748 15886
rect 27692 15822 27694 15874
rect 27746 15822 27748 15874
rect 26572 15316 26628 15326
rect 26460 15314 26628 15316
rect 26460 15262 26574 15314
rect 26626 15262 26628 15314
rect 26460 15260 26628 15262
rect 26572 15250 26628 15260
rect 27692 15204 27748 15822
rect 27692 15138 27748 15148
rect 28252 15764 28308 15774
rect 28252 14644 28308 15708
rect 37660 15764 37716 16046
rect 37660 15698 37716 15708
rect 37660 15314 37716 15326
rect 37660 15262 37662 15314
rect 37714 15262 37716 15314
rect 29484 15204 29540 15214
rect 29484 15110 29540 15148
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 26236 14466 26292 14476
rect 27692 14642 28308 14644
rect 27692 14590 28254 14642
rect 28306 14590 28308 14642
rect 27692 14588 28308 14590
rect 25340 13654 25396 13692
rect 27692 13746 27748 14588
rect 28252 14578 28308 14588
rect 29260 14532 29316 14542
rect 29260 14438 29316 14476
rect 27916 13860 27972 13870
rect 27916 13766 27972 13804
rect 37660 13860 37716 15262
rect 37884 15204 37940 16830
rect 39900 16770 39956 16782
rect 39900 16718 39902 16770
rect 39954 16718 39956 16770
rect 39900 16212 39956 16718
rect 39900 16146 39956 16156
rect 40012 16210 40068 16222
rect 40012 16158 40014 16210
rect 40066 16158 40068 16210
rect 40012 15540 40068 16158
rect 40012 15474 40068 15484
rect 37884 15138 37940 15148
rect 40012 15202 40068 15214
rect 40012 15150 40014 15202
rect 40066 15150 40068 15202
rect 40012 14868 40068 15150
rect 40012 14802 40068 14812
rect 37660 13794 37716 13804
rect 27692 13694 27694 13746
rect 27746 13694 27748 13746
rect 27692 13682 27748 13694
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 26124 3668 26180 3678
rect 26124 3574 26180 3612
rect 25228 3502 25230 3554
rect 25282 3502 25284 3554
rect 25228 3490 25284 3502
rect 16128 0 16240 800
rect 16800 0 16912 800
rect 24864 0 24976 800
<< via2 >>
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 17500 38220 17556 38276
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 1708 36370 1764 36372
rect 1708 36318 1710 36370
rect 1710 36318 1762 36370
rect 1762 36318 1764 36370
rect 1708 36316 1764 36318
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 4172 28252 4228 28308
rect 1932 25564 1988 25620
rect 1932 24498 1988 24500
rect 1932 24446 1934 24498
rect 1934 24446 1986 24498
rect 1986 24446 1988 24498
rect 1932 24444 1988 24446
rect 1932 23548 1988 23604
rect 1932 22930 1988 22932
rect 1932 22878 1934 22930
rect 1934 22878 1986 22930
rect 1986 22878 1988 22930
rect 1932 22876 1988 22878
rect 1932 22482 1988 22484
rect 1932 22430 1934 22482
rect 1934 22430 1986 22482
rect 1986 22430 1988 22482
rect 1932 22428 1988 22430
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 4284 26290 4340 26292
rect 4284 26238 4286 26290
rect 4286 26238 4338 26290
rect 4338 26238 4340 26290
rect 4284 26236 4340 26238
rect 12236 26236 12292 26292
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 12236 25676 12292 25732
rect 14700 25394 14756 25396
rect 14700 25342 14702 25394
rect 14702 25342 14754 25394
rect 14754 25342 14756 25394
rect 14700 25340 14756 25342
rect 14476 24892 14532 24948
rect 4284 24722 4340 24724
rect 4284 24670 4286 24722
rect 4286 24670 4338 24722
rect 4338 24670 4340 24722
rect 4284 24668 4340 24670
rect 12012 24668 12068 24724
rect 14812 24668 14868 24724
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 4284 23938 4340 23940
rect 4284 23886 4286 23938
rect 4286 23886 4338 23938
rect 4338 23886 4340 23938
rect 4284 23884 4340 23886
rect 12236 23884 12292 23940
rect 15260 25676 15316 25732
rect 16156 26460 16212 26516
rect 15484 25452 15540 25508
rect 15596 24946 15652 24948
rect 15596 24894 15598 24946
rect 15598 24894 15650 24946
rect 15650 24894 15652 24946
rect 15596 24892 15652 24894
rect 14924 24556 14980 24612
rect 14476 23324 14532 23380
rect 4284 22988 4340 23044
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 4284 22370 4340 22372
rect 4284 22318 4286 22370
rect 4286 22318 4338 22370
rect 4338 22318 4340 22370
rect 4284 22316 4340 22318
rect 9884 22316 9940 22372
rect 12460 22316 12516 22372
rect 13468 22988 13524 23044
rect 12012 22258 12068 22260
rect 12012 22206 12014 22258
rect 12014 22206 12066 22258
rect 12066 22206 12068 22258
rect 12012 22204 12068 22206
rect 4172 22092 4228 22148
rect 14140 22764 14196 22820
rect 13692 22370 13748 22372
rect 13692 22318 13694 22370
rect 13694 22318 13746 22370
rect 13746 22318 13748 22370
rect 13692 22316 13748 22318
rect 12796 21756 12852 21812
rect 13468 21756 13524 21812
rect 4284 21586 4340 21588
rect 4284 21534 4286 21586
rect 4286 21534 4338 21586
rect 4338 21534 4340 21586
rect 4284 21532 4340 21534
rect 15596 23714 15652 23716
rect 15596 23662 15598 23714
rect 15598 23662 15650 23714
rect 15650 23662 15652 23714
rect 15596 23660 15652 23662
rect 15372 23436 15428 23492
rect 14924 22540 14980 22596
rect 15372 22988 15428 23044
rect 14476 22370 14532 22372
rect 14476 22318 14478 22370
rect 14478 22318 14530 22370
rect 14530 22318 14532 22370
rect 14476 22316 14532 22318
rect 15036 22316 15092 22372
rect 14588 21980 14644 22036
rect 1932 21474 1988 21476
rect 1932 21422 1934 21474
rect 1934 21422 1986 21474
rect 1986 21422 1988 21474
rect 1932 21420 1988 21422
rect 12796 21474 12852 21476
rect 12796 21422 12798 21474
rect 12798 21422 12850 21474
rect 12850 21422 12852 21474
rect 12796 21420 12852 21422
rect 10668 21308 10724 21364
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 12124 20076 12180 20132
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 4284 18450 4340 18452
rect 4284 18398 4286 18450
rect 4286 18398 4338 18450
rect 4338 18398 4340 18450
rect 4284 18396 4340 18398
rect 11452 18450 11508 18452
rect 11452 18398 11454 18450
rect 11454 18398 11506 18450
rect 11506 18398 11508 18450
rect 11452 18396 11508 18398
rect 14476 21868 14532 21924
rect 14252 21474 14308 21476
rect 14252 21422 14254 21474
rect 14254 21422 14306 21474
rect 14306 21422 14308 21474
rect 14252 21420 14308 21422
rect 15260 21362 15316 21364
rect 15260 21310 15262 21362
rect 15262 21310 15314 21362
rect 15314 21310 15316 21362
rect 15260 21308 15316 21310
rect 13580 20076 13636 20132
rect 14476 20076 14532 20132
rect 14924 19740 14980 19796
rect 14700 19516 14756 19572
rect 13804 18508 13860 18564
rect 13244 18284 13300 18340
rect 1932 18226 1988 18228
rect 1932 18174 1934 18226
rect 1934 18174 1986 18226
rect 1986 18174 1988 18226
rect 1932 18172 1988 18174
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 11116 18060 11172 18116
rect 14364 18396 14420 18452
rect 14476 18508 14532 18564
rect 14252 18172 14308 18228
rect 14028 18060 14084 18116
rect 15036 19292 15092 19348
rect 15148 19234 15204 19236
rect 15148 19182 15150 19234
rect 15150 19182 15202 19234
rect 15202 19182 15204 19234
rect 15148 19180 15204 19182
rect 15148 18620 15204 18676
rect 15260 19068 15316 19124
rect 15148 18450 15204 18452
rect 15148 18398 15150 18450
rect 15150 18398 15202 18450
rect 15202 18398 15204 18450
rect 15148 18396 15204 18398
rect 14700 18338 14756 18340
rect 14700 18286 14702 18338
rect 14702 18286 14754 18338
rect 14754 18286 14756 18338
rect 14700 18284 14756 18286
rect 18620 38274 18676 38276
rect 18620 38222 18622 38274
rect 18622 38222 18674 38274
rect 18674 38222 18676 38274
rect 18620 38220 18676 38222
rect 22876 38220 22932 38276
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 18844 37436 18900 37492
rect 20076 37490 20132 37492
rect 20076 37438 20078 37490
rect 20078 37438 20130 37490
rect 20130 37438 20132 37490
rect 20076 37436 20132 37438
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 20524 28588 20580 28644
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 19740 27970 19796 27972
rect 19740 27918 19742 27970
rect 19742 27918 19794 27970
rect 19794 27918 19796 27970
rect 19740 27916 19796 27918
rect 20188 27858 20244 27860
rect 20188 27806 20190 27858
rect 20190 27806 20242 27858
rect 20242 27806 20244 27858
rect 20188 27804 20244 27806
rect 19516 27356 19572 27412
rect 20412 27468 20468 27524
rect 17276 25564 17332 25620
rect 17948 26514 18004 26516
rect 17948 26462 17950 26514
rect 17950 26462 18002 26514
rect 18002 26462 18004 26514
rect 17948 26460 18004 26462
rect 17724 25452 17780 25508
rect 18508 25618 18564 25620
rect 18508 25566 18510 25618
rect 18510 25566 18562 25618
rect 18562 25566 18564 25618
rect 18508 25564 18564 25566
rect 16380 24610 16436 24612
rect 16380 24558 16382 24610
rect 16382 24558 16434 24610
rect 16434 24558 16436 24610
rect 16380 24556 16436 24558
rect 16940 24556 16996 24612
rect 16156 23548 16212 23604
rect 15932 22988 15988 23044
rect 16044 23436 16100 23492
rect 15932 22258 15988 22260
rect 15932 22206 15934 22258
rect 15934 22206 15986 22258
rect 15986 22206 15988 22258
rect 15932 22204 15988 22206
rect 16044 21980 16100 22036
rect 16156 21868 16212 21924
rect 16380 22988 16436 23044
rect 16156 21196 16212 21252
rect 15596 19964 15652 20020
rect 15820 20130 15876 20132
rect 15820 20078 15822 20130
rect 15822 20078 15874 20130
rect 15874 20078 15876 20130
rect 15820 20076 15876 20078
rect 15708 19794 15764 19796
rect 15708 19742 15710 19794
rect 15710 19742 15762 19794
rect 15762 19742 15764 19794
rect 15708 19740 15764 19742
rect 15484 19516 15540 19572
rect 15484 19292 15540 19348
rect 16604 22316 16660 22372
rect 16044 19852 16100 19908
rect 16492 19740 16548 19796
rect 16828 22146 16884 22148
rect 16828 22094 16830 22146
rect 16830 22094 16882 22146
rect 16882 22094 16884 22146
rect 16828 22092 16884 22094
rect 16828 21532 16884 21588
rect 16604 21196 16660 21252
rect 15820 19068 15876 19124
rect 16380 19292 16436 19348
rect 15484 18956 15540 19012
rect 15708 18172 15764 18228
rect 16156 18396 16212 18452
rect 15372 17948 15428 18004
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 14588 15484 14644 15540
rect 14252 15148 14308 15204
rect 15596 15538 15652 15540
rect 15596 15486 15598 15538
rect 15598 15486 15650 15538
rect 15650 15486 15652 15538
rect 15596 15484 15652 15486
rect 15708 15372 15764 15428
rect 15148 15202 15204 15204
rect 15148 15150 15150 15202
rect 15150 15150 15202 15202
rect 15202 15150 15204 15202
rect 15148 15148 15204 15150
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 18172 24610 18228 24612
rect 18172 24558 18174 24610
rect 18174 24558 18226 24610
rect 18226 24558 18228 24610
rect 18172 24556 18228 24558
rect 17276 23100 17332 23156
rect 17276 22764 17332 22820
rect 17164 22540 17220 22596
rect 17612 22652 17668 22708
rect 17836 22540 17892 22596
rect 18396 23714 18452 23716
rect 18396 23662 18398 23714
rect 18398 23662 18450 23714
rect 18450 23662 18452 23714
rect 18396 23660 18452 23662
rect 18844 24108 18900 24164
rect 18956 25506 19012 25508
rect 18956 25454 18958 25506
rect 18958 25454 19010 25506
rect 19010 25454 19012 25506
rect 18956 25452 19012 25454
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 19404 24722 19460 24724
rect 19404 24670 19406 24722
rect 19406 24670 19458 24722
rect 19458 24670 19460 24722
rect 19404 24668 19460 24670
rect 20860 27970 20916 27972
rect 20860 27918 20862 27970
rect 20862 27918 20914 27970
rect 20914 27918 20916 27970
rect 20860 27916 20916 27918
rect 20188 25452 20244 25508
rect 21308 26962 21364 26964
rect 21308 26910 21310 26962
rect 21310 26910 21362 26962
rect 21362 26910 21364 26962
rect 21308 26908 21364 26910
rect 20748 25228 20804 25284
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 19628 24556 19684 24612
rect 18732 23884 18788 23940
rect 18732 23548 18788 23604
rect 19628 23996 19684 24052
rect 18396 23378 18452 23380
rect 18396 23326 18398 23378
rect 18398 23326 18450 23378
rect 18450 23326 18452 23378
rect 18396 23324 18452 23326
rect 18732 23324 18788 23380
rect 18620 23266 18676 23268
rect 18620 23214 18622 23266
rect 18622 23214 18674 23266
rect 18674 23214 18676 23266
rect 18620 23212 18676 23214
rect 17948 22092 18004 22148
rect 18060 21980 18116 22036
rect 18060 21362 18116 21364
rect 18060 21310 18062 21362
rect 18062 21310 18114 21362
rect 18114 21310 18116 21362
rect 18060 21308 18116 21310
rect 17612 20076 17668 20132
rect 17164 19852 17220 19908
rect 16940 19180 16996 19236
rect 17612 19740 17668 19796
rect 17948 19852 18004 19908
rect 17836 19180 17892 19236
rect 17276 19122 17332 19124
rect 17276 19070 17278 19122
rect 17278 19070 17330 19122
rect 17330 19070 17332 19122
rect 17276 19068 17332 19070
rect 16940 19010 16996 19012
rect 16940 18958 16942 19010
rect 16942 18958 16994 19010
rect 16994 18958 16996 19010
rect 16940 18956 16996 18958
rect 17724 18508 17780 18564
rect 16492 17948 16548 18004
rect 16380 15426 16436 15428
rect 16380 15374 16382 15426
rect 16382 15374 16434 15426
rect 16434 15374 16436 15426
rect 16380 15372 16436 15374
rect 18732 22988 18788 23044
rect 18620 22652 18676 22708
rect 18396 22146 18452 22148
rect 18396 22094 18398 22146
rect 18398 22094 18450 22146
rect 18450 22094 18452 22146
rect 18396 22092 18452 22094
rect 18508 21474 18564 21476
rect 18508 21422 18510 21474
rect 18510 21422 18562 21474
rect 18562 21422 18564 21474
rect 18508 21420 18564 21422
rect 19292 23772 19348 23828
rect 19068 23436 19124 23492
rect 19068 22428 19124 22484
rect 18956 21308 19012 21364
rect 18396 19852 18452 19908
rect 18396 18956 18452 19012
rect 18732 20130 18788 20132
rect 18732 20078 18734 20130
rect 18734 20078 18786 20130
rect 18786 20078 18788 20130
rect 18732 20076 18788 20078
rect 18620 20018 18676 20020
rect 18620 19966 18622 20018
rect 18622 19966 18674 20018
rect 18674 19966 18676 20018
rect 18620 19964 18676 19966
rect 18620 19234 18676 19236
rect 18620 19182 18622 19234
rect 18622 19182 18674 19234
rect 18674 19182 18676 19234
rect 18620 19180 18676 19182
rect 15932 15090 15988 15092
rect 15932 15038 15934 15090
rect 15934 15038 15986 15090
rect 15986 15038 15988 15090
rect 15932 15036 15988 15038
rect 19404 23436 19460 23492
rect 21980 37996 22036 38052
rect 24556 38050 24612 38052
rect 24556 37998 24558 38050
rect 24558 37998 24610 38050
rect 24610 37998 24612 38050
rect 24556 37996 24612 37998
rect 25564 38274 25620 38276
rect 25564 38222 25566 38274
rect 25566 38222 25618 38274
rect 25618 38222 25620 38274
rect 25564 38220 25620 38222
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 24892 37436 24948 37492
rect 26236 37490 26292 37492
rect 26236 37438 26238 37490
rect 26238 37438 26290 37490
rect 26290 37438 26292 37490
rect 26236 37436 26292 37438
rect 21868 28642 21924 28644
rect 21868 28590 21870 28642
rect 21870 28590 21922 28642
rect 21922 28590 21924 28642
rect 21868 28588 21924 28590
rect 21756 27804 21812 27860
rect 21644 27468 21700 27524
rect 23548 27858 23604 27860
rect 23548 27806 23550 27858
rect 23550 27806 23602 27858
rect 23602 27806 23604 27858
rect 23548 27804 23604 27806
rect 21868 27074 21924 27076
rect 21868 27022 21870 27074
rect 21870 27022 21922 27074
rect 21922 27022 21924 27074
rect 21868 27020 21924 27022
rect 22652 27020 22708 27076
rect 21868 24668 21924 24724
rect 21980 25228 22036 25284
rect 21532 24556 21588 24612
rect 21532 24220 21588 24276
rect 19740 23826 19796 23828
rect 19740 23774 19742 23826
rect 19742 23774 19794 23826
rect 19794 23774 19796 23826
rect 19740 23772 19796 23774
rect 20188 23938 20244 23940
rect 20188 23886 20190 23938
rect 20190 23886 20242 23938
rect 20242 23886 20244 23938
rect 20188 23884 20244 23886
rect 21532 23996 21588 24052
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 19292 22540 19348 22596
rect 19292 22092 19348 22148
rect 19516 23212 19572 23268
rect 19628 22594 19684 22596
rect 19628 22542 19630 22594
rect 19630 22542 19682 22594
rect 19682 22542 19684 22594
rect 19628 22540 19684 22542
rect 19852 23154 19908 23156
rect 19852 23102 19854 23154
rect 19854 23102 19906 23154
rect 19906 23102 19908 23154
rect 19852 23100 19908 23102
rect 20188 23100 20244 23156
rect 20188 22652 20244 22708
rect 19516 21980 19572 22036
rect 22204 24610 22260 24612
rect 22204 24558 22206 24610
rect 22206 24558 22258 24610
rect 22258 24558 22260 24610
rect 22204 24556 22260 24558
rect 21308 23324 21364 23380
rect 20748 23100 20804 23156
rect 19292 21586 19348 21588
rect 19292 21534 19294 21586
rect 19294 21534 19346 21586
rect 19346 21534 19348 21586
rect 19292 21532 19348 21534
rect 19852 22258 19908 22260
rect 19852 22206 19854 22258
rect 19854 22206 19906 22258
rect 19906 22206 19908 22258
rect 19852 22204 19908 22206
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 19180 19292 19236 19348
rect 20076 20802 20132 20804
rect 20076 20750 20078 20802
rect 20078 20750 20130 20802
rect 20130 20750 20132 20802
rect 20076 20748 20132 20750
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 20524 22316 20580 22372
rect 18956 19180 19012 19236
rect 18284 16044 18340 16100
rect 19068 16882 19124 16884
rect 19068 16830 19070 16882
rect 19070 16830 19122 16882
rect 19122 16830 19124 16882
rect 19068 16828 19124 16830
rect 19068 16098 19124 16100
rect 19068 16046 19070 16098
rect 19070 16046 19122 16098
rect 19122 16046 19124 16098
rect 19068 16044 19124 16046
rect 19404 20076 19460 20132
rect 19852 20130 19908 20132
rect 19852 20078 19854 20130
rect 19854 20078 19906 20130
rect 19906 20078 19908 20130
rect 19852 20076 19908 20078
rect 19516 18620 19572 18676
rect 19404 16828 19460 16884
rect 19628 19180 19684 19236
rect 20188 19852 20244 19908
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 20524 19852 20580 19908
rect 20076 18060 20132 18116
rect 20412 18172 20468 18228
rect 21308 22652 21364 22708
rect 22092 24108 22148 24164
rect 21980 23378 22036 23380
rect 21980 23326 21982 23378
rect 21982 23326 22034 23378
rect 22034 23326 22036 23378
rect 21980 23324 22036 23326
rect 22204 23492 22260 23548
rect 22652 24722 22708 24724
rect 22652 24670 22654 24722
rect 22654 24670 22706 24722
rect 22706 24670 22708 24722
rect 22652 24668 22708 24670
rect 22652 24108 22708 24164
rect 22540 23548 22596 23604
rect 22428 23436 22484 23492
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 23660 25900 23716 25956
rect 24668 25900 24724 25956
rect 22988 24050 23044 24052
rect 22988 23998 22990 24050
rect 22990 23998 23042 24050
rect 23042 23998 23044 24050
rect 22988 23996 23044 23998
rect 22988 23548 23044 23604
rect 22764 23436 22820 23492
rect 23772 24668 23828 24724
rect 23436 24220 23492 24276
rect 23324 23826 23380 23828
rect 23324 23774 23326 23826
rect 23326 23774 23378 23826
rect 23378 23774 23380 23826
rect 23324 23772 23380 23774
rect 23212 23660 23268 23716
rect 22428 23212 22484 23268
rect 21308 22370 21364 22372
rect 21308 22318 21310 22370
rect 21310 22318 21362 22370
rect 21362 22318 21364 22370
rect 21308 22316 21364 22318
rect 21980 22316 22036 22372
rect 20860 21420 20916 21476
rect 20860 20636 20916 20692
rect 21420 22258 21476 22260
rect 21420 22206 21422 22258
rect 21422 22206 21474 22258
rect 21474 22206 21476 22258
rect 21420 22204 21476 22206
rect 21308 20076 21364 20132
rect 22204 22204 22260 22260
rect 21644 20690 21700 20692
rect 21644 20638 21646 20690
rect 21646 20638 21698 20690
rect 21698 20638 21700 20690
rect 21644 20636 21700 20638
rect 21420 19740 21476 19796
rect 22092 21196 22148 21252
rect 21420 18674 21476 18676
rect 21420 18622 21422 18674
rect 21422 18622 21474 18674
rect 21474 18622 21476 18674
rect 21420 18620 21476 18622
rect 20860 18562 20916 18564
rect 20860 18510 20862 18562
rect 20862 18510 20914 18562
rect 20914 18510 20916 18562
rect 20860 18508 20916 18510
rect 20748 18060 20804 18116
rect 21420 18284 21476 18340
rect 20076 17442 20132 17444
rect 20076 17390 20078 17442
rect 20078 17390 20130 17442
rect 20130 17390 20132 17442
rect 20076 17388 20132 17390
rect 21084 17388 21140 17444
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 19964 16828 20020 16884
rect 18844 15932 18900 15988
rect 16604 13468 16660 13524
rect 15708 12796 15764 12852
rect 16156 12850 16212 12852
rect 16156 12798 16158 12850
rect 16158 12798 16210 12850
rect 16210 12798 16212 12850
rect 16156 12796 16212 12798
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 16044 11564 16100 11620
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 20188 16098 20244 16100
rect 20188 16046 20190 16098
rect 20190 16046 20242 16098
rect 20242 16046 20244 16098
rect 20188 16044 20244 16046
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 19516 15148 19572 15204
rect 20524 15484 20580 15540
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 19180 13468 19236 13524
rect 22428 19404 22484 19460
rect 22540 20076 22596 20132
rect 22204 19292 22260 19348
rect 22428 19068 22484 19124
rect 22092 18450 22148 18452
rect 22092 18398 22094 18450
rect 22094 18398 22146 18450
rect 22146 18398 22148 18450
rect 22092 18396 22148 18398
rect 22876 23154 22932 23156
rect 22876 23102 22878 23154
rect 22878 23102 22930 23154
rect 22930 23102 22932 23154
rect 22876 23100 22932 23102
rect 22876 22652 22932 22708
rect 23100 22988 23156 23044
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 27580 24892 27636 24948
rect 25340 24668 25396 24724
rect 26460 24722 26516 24724
rect 26460 24670 26462 24722
rect 26462 24670 26514 24722
rect 26514 24670 26516 24722
rect 26460 24668 26516 24670
rect 24556 23826 24612 23828
rect 24556 23774 24558 23826
rect 24558 23774 24610 23826
rect 24610 23774 24612 23826
rect 24556 23772 24612 23774
rect 25452 23660 25508 23716
rect 26348 23548 26404 23604
rect 24332 23266 24388 23268
rect 24332 23214 24334 23266
rect 24334 23214 24386 23266
rect 24386 23214 24388 23266
rect 24332 23212 24388 23214
rect 26460 23266 26516 23268
rect 26460 23214 26462 23266
rect 26462 23214 26514 23266
rect 26514 23214 26516 23266
rect 26460 23212 26516 23214
rect 23324 22876 23380 22932
rect 23772 22428 23828 22484
rect 23436 22370 23492 22372
rect 23436 22318 23438 22370
rect 23438 22318 23490 22370
rect 23490 22318 23492 22370
rect 23436 22316 23492 22318
rect 23100 22204 23156 22260
rect 22876 20802 22932 20804
rect 22876 20750 22878 20802
rect 22878 20750 22930 20802
rect 22930 20750 22932 20802
rect 22876 20748 22932 20750
rect 25116 23100 25172 23156
rect 24444 22930 24500 22932
rect 24444 22878 24446 22930
rect 24446 22878 24498 22930
rect 24498 22878 24500 22930
rect 24444 22876 24500 22878
rect 26124 23154 26180 23156
rect 26124 23102 26126 23154
rect 26126 23102 26178 23154
rect 26178 23102 26180 23154
rect 26124 23100 26180 23102
rect 26796 24220 26852 24276
rect 26684 24050 26740 24052
rect 26684 23998 26686 24050
rect 26686 23998 26738 24050
rect 26738 23998 26740 24050
rect 26684 23996 26740 23998
rect 27132 24050 27188 24052
rect 27132 23998 27134 24050
rect 27134 23998 27186 24050
rect 27186 23998 27188 24050
rect 27132 23996 27188 23998
rect 26908 23212 26964 23268
rect 25228 23042 25284 23044
rect 25228 22990 25230 23042
rect 25230 22990 25282 23042
rect 25282 22990 25284 23042
rect 25228 22988 25284 22990
rect 24444 22092 24500 22148
rect 24108 21196 24164 21252
rect 24220 20130 24276 20132
rect 24220 20078 24222 20130
rect 24222 20078 24274 20130
rect 24274 20078 24276 20130
rect 24220 20076 24276 20078
rect 25340 21810 25396 21812
rect 25340 21758 25342 21810
rect 25342 21758 25394 21810
rect 25394 21758 25396 21810
rect 25340 21756 25396 21758
rect 25340 21532 25396 21588
rect 25676 22988 25732 23044
rect 26236 22540 26292 22596
rect 25788 22428 25844 22484
rect 25900 21756 25956 21812
rect 25004 20076 25060 20132
rect 22764 19794 22820 19796
rect 22764 19742 22766 19794
rect 22766 19742 22818 19794
rect 22818 19742 22820 19794
rect 22764 19740 22820 19742
rect 23548 19458 23604 19460
rect 23548 19406 23550 19458
rect 23550 19406 23602 19458
rect 23602 19406 23604 19458
rect 23548 19404 23604 19406
rect 22652 18956 22708 19012
rect 22428 18508 22484 18564
rect 22876 18396 22932 18452
rect 23660 19122 23716 19124
rect 23660 19070 23662 19122
rect 23662 19070 23714 19122
rect 23714 19070 23716 19122
rect 23660 19068 23716 19070
rect 23324 18674 23380 18676
rect 23324 18622 23326 18674
rect 23326 18622 23378 18674
rect 23378 18622 23380 18674
rect 23324 18620 23380 18622
rect 23212 18284 23268 18340
rect 23436 18396 23492 18452
rect 22652 18226 22708 18228
rect 22652 18174 22654 18226
rect 22654 18174 22706 18226
rect 22706 18174 22708 18226
rect 22652 18172 22708 18174
rect 22204 17948 22260 18004
rect 22876 16716 22932 16772
rect 23100 15538 23156 15540
rect 23100 15486 23102 15538
rect 23102 15486 23154 15538
rect 23154 15486 23156 15538
rect 23100 15484 23156 15486
rect 20300 13746 20356 13748
rect 20300 13694 20302 13746
rect 20302 13694 20354 13746
rect 20354 13694 20356 13746
rect 20300 13692 20356 13694
rect 22092 13692 22148 13748
rect 20188 13468 20244 13524
rect 25564 19516 25620 19572
rect 25788 20076 25844 20132
rect 25116 19180 25172 19236
rect 25676 19234 25732 19236
rect 25676 19182 25678 19234
rect 25678 19182 25730 19234
rect 25730 19182 25732 19234
rect 25676 19180 25732 19182
rect 25228 19068 25284 19124
rect 25340 19122 25396 19124
rect 25340 19070 25342 19122
rect 25342 19070 25394 19122
rect 25394 19070 25396 19122
rect 25340 19068 25396 19070
rect 25676 18956 25732 19012
rect 24668 18508 24724 18564
rect 23772 18338 23828 18340
rect 23772 18286 23774 18338
rect 23774 18286 23826 18338
rect 23826 18286 23828 18338
rect 23772 18284 23828 18286
rect 23996 18450 24052 18452
rect 23996 18398 23998 18450
rect 23998 18398 24050 18450
rect 24050 18398 24052 18450
rect 23996 18396 24052 18398
rect 26012 21586 26068 21588
rect 26012 21534 26014 21586
rect 26014 21534 26066 21586
rect 26066 21534 26068 21586
rect 26012 21532 26068 21534
rect 25900 18620 25956 18676
rect 26796 22428 26852 22484
rect 26572 21586 26628 21588
rect 26572 21534 26574 21586
rect 26574 21534 26626 21586
rect 26626 21534 26628 21586
rect 26572 21532 26628 21534
rect 26236 19010 26292 19012
rect 26236 18958 26238 19010
rect 26238 18958 26290 19010
rect 26290 18958 26292 19010
rect 26236 18956 26292 18958
rect 27356 23826 27412 23828
rect 27356 23774 27358 23826
rect 27358 23774 27410 23826
rect 27410 23774 27412 23826
rect 27356 23772 27412 23774
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 28028 23884 28084 23940
rect 27580 23548 27636 23604
rect 29708 23884 29764 23940
rect 27916 23212 27972 23268
rect 27020 22988 27076 23044
rect 37660 23938 37716 23940
rect 37660 23886 37662 23938
rect 37662 23886 37714 23938
rect 37714 23886 37716 23938
rect 37660 23884 37716 23886
rect 40012 24220 40068 24276
rect 37884 23772 37940 23828
rect 40012 23548 40068 23604
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 26796 19346 26852 19348
rect 26796 19294 26798 19346
rect 26798 19294 26850 19346
rect 26850 19294 26852 19346
rect 26796 19292 26852 19294
rect 26572 19234 26628 19236
rect 26572 19182 26574 19234
rect 26574 19182 26626 19234
rect 26626 19182 26628 19234
rect 26572 19180 26628 19182
rect 26684 18956 26740 19012
rect 26124 18508 26180 18564
rect 25788 18450 25844 18452
rect 25788 18398 25790 18450
rect 25790 18398 25842 18450
rect 25842 18398 25844 18450
rect 25788 18396 25844 18398
rect 23772 16828 23828 16884
rect 25452 16716 25508 16772
rect 24444 16044 24500 16100
rect 25788 16044 25844 16100
rect 25228 15932 25284 15988
rect 23436 15314 23492 15316
rect 23436 15262 23438 15314
rect 23438 15262 23490 15314
rect 23490 15262 23492 15314
rect 23436 15260 23492 15262
rect 25340 15314 25396 15316
rect 25340 15262 25342 15314
rect 25342 15262 25394 15314
rect 25394 15262 25396 15314
rect 25340 15260 25396 15262
rect 25900 15986 25956 15988
rect 25900 15934 25902 15986
rect 25902 15934 25954 15986
rect 25954 15934 25956 15986
rect 25900 15932 25956 15934
rect 23548 13746 23604 13748
rect 23548 13694 23550 13746
rect 23550 13694 23602 13746
rect 23602 13694 23604 13746
rect 23548 13692 23604 13694
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 17388 11564 17444 11620
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 16156 4172 16212 4228
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 18508 4226 18564 4228
rect 18508 4174 18510 4226
rect 18510 4174 18562 4226
rect 18562 4174 18564 4226
rect 18508 4172 18564 4174
rect 24892 3612 24948 3668
rect 16828 3388 16884 3444
rect 18060 3388 18116 3444
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 27356 22540 27412 22596
rect 28588 22540 28644 22596
rect 40012 22930 40068 22932
rect 40012 22878 40014 22930
rect 40014 22878 40066 22930
rect 40066 22878 40068 22930
rect 40012 22876 40068 22878
rect 37660 22540 37716 22596
rect 29260 22482 29316 22484
rect 29260 22430 29262 22482
rect 29262 22430 29314 22482
rect 29314 22430 29316 22482
rect 29260 22428 29316 22430
rect 27804 22092 27860 22148
rect 27020 21586 27076 21588
rect 27020 21534 27022 21586
rect 27022 21534 27074 21586
rect 27074 21534 27076 21586
rect 27020 21532 27076 21534
rect 27132 20748 27188 20804
rect 27020 19740 27076 19796
rect 27468 19292 27524 19348
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 29596 19906 29652 19908
rect 29596 19854 29598 19906
rect 29598 19854 29650 19906
rect 29650 19854 29652 19906
rect 29596 19852 29652 19854
rect 27132 18956 27188 19012
rect 26908 18620 26964 18676
rect 27244 18620 27300 18676
rect 26684 18508 26740 18564
rect 27692 18284 27748 18340
rect 27020 16098 27076 16100
rect 27020 16046 27022 16098
rect 27022 16046 27074 16098
rect 27074 16046 27076 16098
rect 27020 16044 27076 16046
rect 27132 15932 27188 15988
rect 26908 15708 26964 15764
rect 25340 14530 25396 14532
rect 25340 14478 25342 14530
rect 25342 14478 25394 14530
rect 25394 14478 25396 14530
rect 25340 14476 25396 14478
rect 40012 20188 40068 20244
rect 37660 19852 37716 19908
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 29596 19068 29652 19124
rect 37660 18450 37716 18452
rect 37660 18398 37662 18450
rect 37662 18398 37714 18450
rect 37714 18398 37716 18450
rect 37660 18396 37716 18398
rect 29484 18338 29540 18340
rect 29484 18286 29486 18338
rect 29486 18286 29538 18338
rect 29538 18286 29540 18338
rect 29484 18284 29540 18286
rect 40012 18226 40068 18228
rect 40012 18174 40014 18226
rect 40014 18174 40066 18226
rect 40066 18174 40068 18226
rect 40012 18172 40068 18174
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 27580 16098 27636 16100
rect 27580 16046 27582 16098
rect 27582 16046 27634 16098
rect 27634 16046 27636 16098
rect 27580 16044 27636 16046
rect 27692 15148 27748 15204
rect 28252 15708 28308 15764
rect 37660 15708 37716 15764
rect 29484 15202 29540 15204
rect 29484 15150 29486 15202
rect 29486 15150 29538 15202
rect 29538 15150 29540 15202
rect 29484 15148 29540 15150
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 26236 14476 26292 14532
rect 25340 13746 25396 13748
rect 25340 13694 25342 13746
rect 25342 13694 25394 13746
rect 25394 13694 25396 13746
rect 25340 13692 25396 13694
rect 29260 14530 29316 14532
rect 29260 14478 29262 14530
rect 29262 14478 29314 14530
rect 29314 14478 29316 14530
rect 29260 14476 29316 14478
rect 27916 13858 27972 13860
rect 27916 13806 27918 13858
rect 27918 13806 27970 13858
rect 27970 13806 27972 13858
rect 27916 13804 27972 13806
rect 39900 16156 39956 16212
rect 40012 15484 40068 15540
rect 37884 15148 37940 15204
rect 40012 14812 40068 14868
rect 37660 13804 37716 13860
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 26124 3666 26180 3668
rect 26124 3614 26126 3666
rect 26126 3614 26178 3666
rect 26178 3614 26180 3666
rect 26124 3612 26180 3614
<< metal3 >>
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 17490 38220 17500 38276
rect 17556 38220 18620 38276
rect 18676 38220 18686 38276
rect 22866 38220 22876 38276
rect 22932 38220 25564 38276
rect 25620 38220 25630 38276
rect 21970 37996 21980 38052
rect 22036 37996 24556 38052
rect 24612 37996 24622 38052
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 18834 37436 18844 37492
rect 18900 37436 20076 37492
rect 20132 37436 20142 37492
rect 24882 37436 24892 37492
rect 24948 37436 26236 37492
rect 26292 37436 26302 37492
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 0 36372 800 36400
rect 0 36316 1708 36372
rect 1764 36316 1774 36372
rect 0 36288 800 36316
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 20514 28588 20524 28644
rect 20580 28588 21868 28644
rect 21924 28588 21934 28644
rect 0 28308 800 28336
rect 0 28252 4172 28308
rect 4228 28252 4238 28308
rect 0 28224 800 28252
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 19730 27916 19740 27972
rect 19796 27916 20860 27972
rect 20916 27916 20926 27972
rect 20178 27804 20188 27860
rect 20244 27804 21756 27860
rect 21812 27804 23548 27860
rect 23604 27804 23614 27860
rect 20402 27468 20412 27524
rect 20468 27468 21644 27524
rect 21700 27468 21710 27524
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 19506 27356 19516 27412
rect 19572 27356 21364 27412
rect 21308 26964 21364 27356
rect 21858 27020 21868 27076
rect 21924 27020 22652 27076
rect 22708 27020 22718 27076
rect 21298 26908 21308 26964
rect 21364 26908 21374 26964
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 16146 26460 16156 26516
rect 16212 26460 17948 26516
rect 18004 26460 18014 26516
rect 4274 26236 4284 26292
rect 4340 26236 12236 26292
rect 12292 26236 12302 26292
rect 23650 25900 23660 25956
rect 23716 25900 24668 25956
rect 24724 25900 24734 25956
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 12226 25676 12236 25732
rect 12292 25676 15260 25732
rect 15316 25676 15326 25732
rect 0 25620 800 25648
rect 0 25564 1932 25620
rect 1988 25564 1998 25620
rect 17266 25564 17276 25620
rect 17332 25564 18508 25620
rect 18564 25564 18574 25620
rect 0 25536 800 25564
rect 15474 25452 15484 25508
rect 15540 25452 17724 25508
rect 17780 25452 18956 25508
rect 19012 25452 20188 25508
rect 20244 25452 20254 25508
rect 14690 25340 14700 25396
rect 14756 25340 15148 25396
rect 15092 25284 15148 25340
rect 15092 25228 20748 25284
rect 20804 25228 21980 25284
rect 22036 25228 22046 25284
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 14466 24892 14476 24948
rect 14532 24892 15596 24948
rect 15652 24892 15662 24948
rect 26852 24892 27580 24948
rect 27636 24892 27646 24948
rect 26852 24724 26908 24892
rect 4274 24668 4284 24724
rect 4340 24668 12012 24724
rect 12068 24668 14812 24724
rect 14868 24668 14878 24724
rect 19394 24668 19404 24724
rect 19460 24668 21868 24724
rect 21924 24668 22652 24724
rect 22708 24668 23772 24724
rect 23828 24668 25340 24724
rect 25396 24668 26460 24724
rect 26516 24668 26908 24724
rect 14914 24556 14924 24612
rect 14980 24556 16380 24612
rect 16436 24556 16940 24612
rect 16996 24556 18172 24612
rect 18228 24556 19628 24612
rect 19684 24556 19694 24612
rect 21522 24556 21532 24612
rect 21588 24556 22204 24612
rect 22260 24556 22270 24612
rect 1922 24444 1932 24500
rect 1988 24444 1998 24500
rect 0 24276 800 24304
rect 1932 24276 1988 24444
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 41200 24276 42000 24304
rect 0 24220 1988 24276
rect 21522 24220 21532 24276
rect 21588 24220 23436 24276
rect 23492 24220 26796 24276
rect 26852 24220 26862 24276
rect 40002 24220 40012 24276
rect 40068 24220 42000 24276
rect 0 24192 800 24220
rect 41200 24192 42000 24220
rect 18834 24108 18844 24164
rect 18900 24108 22092 24164
rect 22148 24108 22652 24164
rect 22708 24108 22718 24164
rect 22988 24108 26908 24164
rect 22988 24052 23044 24108
rect 26852 24052 26908 24108
rect 19618 23996 19628 24052
rect 19684 23996 21532 24052
rect 21588 23996 21598 24052
rect 22978 23996 22988 24052
rect 23044 23996 23054 24052
rect 26674 23996 26684 24052
rect 26740 23996 26750 24052
rect 26852 23996 27132 24052
rect 27188 23996 27198 24052
rect 4274 23884 4284 23940
rect 4340 23884 12236 23940
rect 12292 23884 12302 23940
rect 18722 23884 18732 23940
rect 18788 23884 20188 23940
rect 20244 23884 20254 23940
rect 26684 23828 26740 23996
rect 28018 23884 28028 23940
rect 28084 23884 29708 23940
rect 29764 23884 37660 23940
rect 37716 23884 37726 23940
rect 15596 23772 19292 23828
rect 19348 23772 19740 23828
rect 19796 23772 19806 23828
rect 23314 23772 23324 23828
rect 23380 23772 24556 23828
rect 24612 23772 24622 23828
rect 26684 23772 27356 23828
rect 27412 23772 37884 23828
rect 37940 23772 37950 23828
rect 15596 23716 15652 23772
rect 15586 23660 15596 23716
rect 15652 23660 15662 23716
rect 18386 23660 18396 23716
rect 18452 23660 23212 23716
rect 23268 23660 25452 23716
rect 25508 23660 25518 23716
rect 0 23604 800 23632
rect 41200 23604 42000 23632
rect 0 23548 1932 23604
rect 1988 23548 1998 23604
rect 16146 23548 16156 23604
rect 16212 23548 18732 23604
rect 18788 23548 18798 23604
rect 22530 23548 22540 23604
rect 22596 23548 22988 23604
rect 23044 23548 23054 23604
rect 26338 23548 26348 23604
rect 26404 23548 27580 23604
rect 27636 23548 27646 23604
rect 40002 23548 40012 23604
rect 40068 23548 42000 23604
rect 0 23520 800 23548
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 22194 23492 22204 23548
rect 22260 23492 22270 23548
rect 41200 23520 42000 23548
rect 15362 23436 15372 23492
rect 15428 23436 16044 23492
rect 16100 23436 16110 23492
rect 19058 23436 19068 23492
rect 19124 23436 19404 23492
rect 19460 23436 19470 23492
rect 20188 23436 22260 23492
rect 22418 23436 22428 23492
rect 22484 23436 22522 23492
rect 22726 23436 22764 23492
rect 22820 23436 22830 23492
rect 20188 23380 20244 23436
rect 14466 23324 14476 23380
rect 14532 23324 18396 23380
rect 18452 23324 18462 23380
rect 18722 23324 18732 23380
rect 18788 23324 20244 23380
rect 21298 23324 21308 23380
rect 21364 23324 21980 23380
rect 22036 23324 22046 23380
rect 18610 23212 18620 23268
rect 18676 23212 19516 23268
rect 19572 23212 22428 23268
rect 22484 23212 24332 23268
rect 24388 23212 24398 23268
rect 26450 23212 26460 23268
rect 26516 23212 26908 23268
rect 26964 23212 27916 23268
rect 27972 23212 27982 23268
rect 17266 23100 17276 23156
rect 17332 23100 19852 23156
rect 19908 23100 19918 23156
rect 20178 23100 20188 23156
rect 20244 23100 20748 23156
rect 20804 23100 20814 23156
rect 22418 23100 22428 23156
rect 22484 23100 22876 23156
rect 22932 23100 22942 23156
rect 25106 23100 25116 23156
rect 25172 23100 26124 23156
rect 26180 23100 26190 23156
rect 4274 22988 4284 23044
rect 4340 22988 13468 23044
rect 13524 22988 13534 23044
rect 15362 22988 15372 23044
rect 15428 22988 15932 23044
rect 15988 22988 16380 23044
rect 16436 22988 18732 23044
rect 18788 22988 18798 23044
rect 23090 22988 23100 23044
rect 23156 22988 25228 23044
rect 25284 22988 25294 23044
rect 25666 22988 25676 23044
rect 25732 22988 27020 23044
rect 27076 22988 27086 23044
rect 0 22932 800 22960
rect 41200 22932 42000 22960
rect 0 22876 1932 22932
rect 1988 22876 1998 22932
rect 23314 22876 23324 22932
rect 23380 22876 24444 22932
rect 24500 22876 24510 22932
rect 40002 22876 40012 22932
rect 40068 22876 42000 22932
rect 0 22848 800 22876
rect 41200 22848 42000 22876
rect 14130 22764 14140 22820
rect 14196 22764 17276 22820
rect 17332 22764 17342 22820
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 15092 22652 17612 22708
rect 17668 22652 18620 22708
rect 18676 22652 18686 22708
rect 20178 22652 20188 22708
rect 20244 22652 21308 22708
rect 21364 22652 22876 22708
rect 22932 22652 22942 22708
rect 15092 22596 15148 22652
rect 14914 22540 14924 22596
rect 14980 22540 15148 22596
rect 17154 22540 17164 22596
rect 17220 22540 17836 22596
rect 17892 22540 19292 22596
rect 19348 22540 19358 22596
rect 19618 22540 19628 22596
rect 19684 22540 22764 22596
rect 22820 22540 26236 22596
rect 26292 22540 26302 22596
rect 27346 22540 27356 22596
rect 27412 22540 28588 22596
rect 28644 22540 37660 22596
rect 37716 22540 37726 22596
rect 1922 22428 1932 22484
rect 1988 22428 1998 22484
rect 19058 22428 19068 22484
rect 19124 22428 23772 22484
rect 23828 22428 23838 22484
rect 25778 22428 25788 22484
rect 25844 22428 26796 22484
rect 26852 22428 29260 22484
rect 29316 22428 29326 22484
rect 0 22260 800 22288
rect 1932 22260 1988 22428
rect 4274 22316 4284 22372
rect 4340 22316 9884 22372
rect 9940 22316 12460 22372
rect 12516 22316 13692 22372
rect 13748 22316 14476 22372
rect 14532 22316 14542 22372
rect 15026 22316 15036 22372
rect 15092 22316 16604 22372
rect 16660 22316 16670 22372
rect 20514 22316 20524 22372
rect 20580 22316 21308 22372
rect 21364 22316 21374 22372
rect 21970 22316 21980 22372
rect 22036 22316 23436 22372
rect 23492 22316 23502 22372
rect 0 22204 1988 22260
rect 12002 22204 12012 22260
rect 12068 22204 15932 22260
rect 15988 22204 15998 22260
rect 19842 22204 19852 22260
rect 19908 22204 21420 22260
rect 21476 22204 21486 22260
rect 22194 22204 22204 22260
rect 22260 22204 23100 22260
rect 23156 22204 23166 22260
rect 0 22176 800 22204
rect 4162 22092 4172 22148
rect 4228 22092 16828 22148
rect 16884 22092 16894 22148
rect 17938 22092 17948 22148
rect 18004 22092 18396 22148
rect 18452 22092 19292 22148
rect 19348 22092 19358 22148
rect 24434 22092 24444 22148
rect 24500 22092 27804 22148
rect 27860 22092 27870 22148
rect 14578 21980 14588 22036
rect 14644 21980 16044 22036
rect 16100 21980 16110 22036
rect 18050 21980 18060 22036
rect 18116 21980 19516 22036
rect 19572 21980 19582 22036
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 14466 21868 14476 21924
rect 14532 21868 16156 21924
rect 16212 21868 16222 21924
rect 12786 21756 12796 21812
rect 12852 21756 13468 21812
rect 13524 21756 13534 21812
rect 25330 21756 25340 21812
rect 25396 21756 25900 21812
rect 25956 21756 25966 21812
rect 0 21588 800 21616
rect 0 21532 1988 21588
rect 4274 21532 4284 21588
rect 4340 21532 8428 21588
rect 16818 21532 16828 21588
rect 16884 21532 19292 21588
rect 19348 21532 19358 21588
rect 25330 21532 25340 21588
rect 25396 21532 26012 21588
rect 26068 21532 26078 21588
rect 26562 21532 26572 21588
rect 26628 21532 27020 21588
rect 27076 21532 27086 21588
rect 0 21504 800 21532
rect 1932 21476 1988 21532
rect 1922 21420 1932 21476
rect 1988 21420 1998 21476
rect 8372 21364 8428 21532
rect 12786 21420 12796 21476
rect 12852 21420 14252 21476
rect 14308 21420 14318 21476
rect 18498 21420 18508 21476
rect 18564 21420 20860 21476
rect 20916 21420 20926 21476
rect 8372 21308 10668 21364
rect 10724 21308 15260 21364
rect 15316 21308 15326 21364
rect 18050 21308 18060 21364
rect 18116 21308 18956 21364
rect 19012 21308 19022 21364
rect 16146 21196 16156 21252
rect 16212 21196 16604 21252
rect 16660 21196 22092 21252
rect 22148 21196 24108 21252
rect 24164 21196 24174 21252
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 20066 20748 20076 20804
rect 20132 20748 22876 20804
rect 22932 20748 22942 20804
rect 26852 20748 27132 20804
rect 27188 20748 27198 20804
rect 26852 20692 26908 20748
rect 20850 20636 20860 20692
rect 20916 20636 21644 20692
rect 21700 20636 26908 20692
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 41200 20244 42000 20272
rect 40002 20188 40012 20244
rect 40068 20188 42000 20244
rect 41200 20160 42000 20188
rect 12114 20076 12124 20132
rect 12180 20076 13580 20132
rect 13636 20076 13646 20132
rect 14466 20076 14476 20132
rect 14532 20076 15820 20132
rect 15876 20076 15886 20132
rect 17602 20076 17612 20132
rect 17668 20076 18732 20132
rect 18788 20076 19404 20132
rect 19460 20076 19852 20132
rect 19908 20076 21308 20132
rect 21364 20076 21374 20132
rect 22530 20076 22540 20132
rect 22596 20076 24220 20132
rect 24276 20076 25004 20132
rect 25060 20076 25788 20132
rect 25844 20076 25854 20132
rect 15586 19964 15596 20020
rect 15652 19964 18620 20020
rect 18676 19964 18686 20020
rect 16034 19852 16044 19908
rect 16100 19852 17164 19908
rect 17220 19852 17948 19908
rect 18004 19852 18014 19908
rect 18386 19852 18396 19908
rect 18452 19852 20188 19908
rect 20244 19852 20524 19908
rect 20580 19852 20590 19908
rect 29586 19852 29596 19908
rect 29652 19852 37660 19908
rect 37716 19852 37726 19908
rect 14914 19740 14924 19796
rect 14980 19740 15708 19796
rect 15764 19740 15774 19796
rect 16482 19740 16492 19796
rect 16548 19740 17612 19796
rect 17668 19740 21420 19796
rect 21476 19740 21486 19796
rect 22754 19740 22764 19796
rect 22820 19740 27020 19796
rect 27076 19740 27086 19796
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 14690 19516 14700 19572
rect 14756 19516 15484 19572
rect 15540 19516 25564 19572
rect 25620 19516 25630 19572
rect 22418 19404 22428 19460
rect 22484 19404 23548 19460
rect 23604 19404 23614 19460
rect 15026 19292 15036 19348
rect 15092 19292 15484 19348
rect 15540 19292 15550 19348
rect 16370 19292 16380 19348
rect 16436 19292 19180 19348
rect 19236 19292 22204 19348
rect 22260 19292 22270 19348
rect 15138 19180 15148 19236
rect 15204 19180 16940 19236
rect 16996 19180 17836 19236
rect 17892 19180 17902 19236
rect 18610 19180 18620 19236
rect 18676 19180 18956 19236
rect 19012 19180 19628 19236
rect 19684 19180 19694 19236
rect 19852 19180 25116 19236
rect 25172 19180 25182 19236
rect 19852 19124 19908 19180
rect 25340 19124 25396 19516
rect 26786 19292 26796 19348
rect 26852 19292 27468 19348
rect 27524 19292 27534 19348
rect 25666 19180 25676 19236
rect 25732 19180 26572 19236
rect 26628 19180 26638 19236
rect 15250 19068 15260 19124
rect 15316 19068 15820 19124
rect 15876 19068 17276 19124
rect 17332 19068 19908 19124
rect 22418 19068 22428 19124
rect 22484 19068 23660 19124
rect 23716 19068 23726 19124
rect 25218 19068 25228 19124
rect 25284 19068 25340 19124
rect 25396 19068 25406 19124
rect 26012 19068 29596 19124
rect 29652 19068 29662 19124
rect 26012 19012 26068 19068
rect 15474 18956 15484 19012
rect 15540 18956 16940 19012
rect 16996 18956 18396 19012
rect 18452 18956 22652 19012
rect 22708 18956 22718 19012
rect 25666 18956 25676 19012
rect 25732 18956 26068 19012
rect 26226 18956 26236 19012
rect 26292 18956 26302 19012
rect 26674 18956 26684 19012
rect 26740 18956 27132 19012
rect 27188 18956 27198 19012
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 26236 18676 26292 18956
rect 15092 18564 15148 18676
rect 15204 18620 15214 18676
rect 19506 18620 19516 18676
rect 19572 18620 21420 18676
rect 21476 18620 21486 18676
rect 23314 18620 23324 18676
rect 23380 18620 25900 18676
rect 25956 18620 25966 18676
rect 26236 18620 26908 18676
rect 26964 18620 27244 18676
rect 27300 18620 27310 18676
rect 13794 18508 13804 18564
rect 13860 18508 14476 18564
rect 14532 18508 15148 18564
rect 17714 18508 17724 18564
rect 17780 18508 20860 18564
rect 20916 18508 22428 18564
rect 22484 18508 22494 18564
rect 24658 18508 24668 18564
rect 24724 18508 26124 18564
rect 26180 18508 26684 18564
rect 26740 18508 26750 18564
rect 13804 18452 13860 18508
rect 4274 18396 4284 18452
rect 4340 18396 8428 18452
rect 11442 18396 11452 18452
rect 11508 18396 13860 18452
rect 14354 18396 14364 18452
rect 14420 18396 15148 18452
rect 15204 18396 16156 18452
rect 16212 18396 16222 18452
rect 22082 18396 22092 18452
rect 22148 18396 22876 18452
rect 22932 18396 23436 18452
rect 23492 18396 23996 18452
rect 24052 18396 24062 18452
rect 25778 18396 25788 18452
rect 25844 18396 25854 18452
rect 31892 18396 37660 18452
rect 37716 18396 37726 18452
rect 0 18228 800 18256
rect 0 18172 1932 18228
rect 1988 18172 1998 18228
rect 0 18144 800 18172
rect 8372 18116 8428 18396
rect 13234 18284 13244 18340
rect 13300 18284 14700 18340
rect 14756 18284 14766 18340
rect 21410 18284 21420 18340
rect 21476 18284 23212 18340
rect 23268 18284 23772 18340
rect 23828 18284 23838 18340
rect 14242 18172 14252 18228
rect 14308 18172 15708 18228
rect 15764 18172 20412 18228
rect 20468 18172 22652 18228
rect 22708 18172 22718 18228
rect 25788 18116 25844 18396
rect 31892 18340 31948 18396
rect 27682 18284 27692 18340
rect 27748 18284 29484 18340
rect 29540 18284 31948 18340
rect 41200 18228 42000 18256
rect 40002 18172 40012 18228
rect 40068 18172 42000 18228
rect 41200 18144 42000 18172
rect 8372 18060 11116 18116
rect 11172 18060 14028 18116
rect 14084 18060 14094 18116
rect 20066 18060 20076 18116
rect 20132 18060 20748 18116
rect 20804 18060 25844 18116
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 15362 17948 15372 18004
rect 15428 17948 16492 18004
rect 16548 17948 22204 18004
rect 22260 17948 22270 18004
rect 20066 17388 20076 17444
rect 20132 17388 21084 17444
rect 21140 17388 21150 17444
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 19058 16828 19068 16884
rect 19124 16828 19404 16884
rect 19460 16828 19964 16884
rect 20020 16828 23772 16884
rect 23828 16828 23838 16884
rect 22866 16716 22876 16772
rect 22932 16716 25452 16772
rect 25508 16716 25518 16772
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 41200 16212 42000 16240
rect 39890 16156 39900 16212
rect 39956 16156 42000 16212
rect 41200 16128 42000 16156
rect 18274 16044 18284 16100
rect 18340 16044 19068 16100
rect 19124 16044 20188 16100
rect 20244 16044 20254 16100
rect 24434 16044 24444 16100
rect 24500 16044 25788 16100
rect 25844 16044 27020 16100
rect 27076 16044 27580 16100
rect 27636 16044 27646 16100
rect 18834 15932 18844 15988
rect 18900 15932 25228 15988
rect 25284 15932 25900 15988
rect 25956 15932 27132 15988
rect 27188 15932 27198 15988
rect 26898 15708 26908 15764
rect 26964 15708 28252 15764
rect 28308 15708 37660 15764
rect 37716 15708 37726 15764
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 41200 15540 42000 15568
rect 14578 15484 14588 15540
rect 14644 15484 15596 15540
rect 15652 15484 15662 15540
rect 20514 15484 20524 15540
rect 20580 15484 23100 15540
rect 23156 15484 23166 15540
rect 40002 15484 40012 15540
rect 40068 15484 42000 15540
rect 41200 15456 42000 15484
rect 15698 15372 15708 15428
rect 15764 15372 16380 15428
rect 16436 15372 16446 15428
rect 23426 15260 23436 15316
rect 23492 15260 25340 15316
rect 25396 15260 25406 15316
rect 14242 15148 14252 15204
rect 14308 15148 15148 15204
rect 15204 15148 15214 15204
rect 15932 15148 19516 15204
rect 19572 15148 19582 15204
rect 27682 15148 27692 15204
rect 27748 15148 29484 15204
rect 29540 15148 37884 15204
rect 37940 15148 37950 15204
rect 15932 15092 15988 15148
rect 15922 15036 15932 15092
rect 15988 15036 15998 15092
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 41200 14868 42000 14896
rect 40002 14812 40012 14868
rect 40068 14812 42000 14868
rect 41200 14784 42000 14812
rect 25330 14476 25340 14532
rect 25396 14476 26236 14532
rect 26292 14476 29260 14532
rect 29316 14476 29326 14532
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 27906 13804 27916 13860
rect 27972 13804 37660 13860
rect 37716 13804 37726 13860
rect 20290 13692 20300 13748
rect 20356 13692 22092 13748
rect 22148 13692 23548 13748
rect 23604 13692 25340 13748
rect 25396 13692 25406 13748
rect 16594 13468 16604 13524
rect 16660 13468 19180 13524
rect 19236 13468 20188 13524
rect 20244 13468 20254 13524
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 15698 12796 15708 12852
rect 15764 12796 16156 12852
rect 16212 12796 16222 12852
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 16034 11564 16044 11620
rect 16100 11564 17388 11620
rect 17444 11564 17454 11620
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 16146 4172 16156 4228
rect 16212 4172 18508 4228
rect 18564 4172 18574 4228
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 24882 3612 24892 3668
rect 24948 3612 26124 3668
rect 26180 3612 26190 3668
rect 16818 3388 16828 3444
rect 16884 3388 18060 3444
rect 18116 3388 18126 3444
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
<< via3 >>
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 22428 23436 22484 23492
rect 22764 23436 22820 23492
rect 22428 23100 22484 23156
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 22764 22540 22820 22596
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
<< metal4 >>
rect 4448 38444 4768 38476
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 37660 20128 38476
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19808 34524 20128 36036
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 19808 23548 20128 25060
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 35168 38444 35488 38476
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 19808 21980 20128 23492
rect 22428 23492 22484 23502
rect 22428 23156 22484 23436
rect 22428 23090 22484 23100
rect 22764 23492 22820 23502
rect 22764 22596 22820 23436
rect 22764 22530 22820 22540
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _108_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 22288 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _109_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 25760 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _110_
timestamp 1698175906
transform 1 0 22960 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _111_
timestamp 1698175906
transform -1 0 24304 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _112_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 23968 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _113_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 27440 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _114_
timestamp 1698175906
transform -1 0 20272 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _115_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18480 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _116_
timestamp 1698175906
transform 1 0 18592 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _117_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 27776 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _118_
timestamp 1698175906
transform 1 0 20944 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _119_
timestamp 1698175906
transform 1 0 23744 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _120_
timestamp 1698175906
transform -1 0 22736 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _121_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 20944 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _122_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19152 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _123_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 22288 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _124_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 22064 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _125_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18480 0 -1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _126_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 20944 0 -1 20384
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _127_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21168 0 1 23520
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _128_
timestamp 1698175906
transform -1 0 23856 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _129_
timestamp 1698175906
transform -1 0 22288 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _130_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19712 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _131_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 18256 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _132_
timestamp 1698175906
transform -1 0 19264 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _133_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 20832 0 1 23520
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _134_
timestamp 1698175906
transform 1 0 17472 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _135_
timestamp 1698175906
transform 1 0 17584 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _136_
timestamp 1698175906
transform -1 0 16016 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _137_
timestamp 1698175906
transform -1 0 17136 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _138_
timestamp 1698175906
transform -1 0 23408 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _139_
timestamp 1698175906
transform 1 0 23072 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _140_
timestamp 1698175906
transform 1 0 23744 0 -1 23520
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _141_
timestamp 1698175906
transform 1 0 27440 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _142_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 23520 0 -1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _143_
timestamp 1698175906
transform -1 0 28336 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _144_
timestamp 1698175906
transform -1 0 23072 0 -1 20384
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _145_
timestamp 1698175906
transform -1 0 26096 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _146_
timestamp 1698175906
transform 1 0 25200 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _147_
timestamp 1698175906
transform 1 0 26544 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _148_
timestamp 1698175906
transform -1 0 17808 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _149_
timestamp 1698175906
transform -1 0 15344 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _150_
timestamp 1698175906
transform -1 0 14672 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _151_
timestamp 1698175906
transform -1 0 18480 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _152_
timestamp 1698175906
transform 1 0 17024 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _153_
timestamp 1698175906
transform -1 0 14112 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _154_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18144 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _155_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 21728 0 -1 18816
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _156_
timestamp 1698175906
transform 1 0 18928 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _157_
timestamp 1698175906
transform 1 0 19824 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _158_
timestamp 1698175906
transform -1 0 19264 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _159_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 18928 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _160_
timestamp 1698175906
transform 1 0 19040 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _161_
timestamp 1698175906
transform 1 0 19936 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _162_
timestamp 1698175906
transform 1 0 18928 0 1 21952
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _163_
timestamp 1698175906
transform -1 0 19152 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _164_
timestamp 1698175906
transform 1 0 26768 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _165_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 26768 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _166_
timestamp 1698175906
transform -1 0 25872 0 -1 18816
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _167_
timestamp 1698175906
transform -1 0 27216 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _168_
timestamp 1698175906
transform -1 0 26656 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _169_
timestamp 1698175906
transform 1 0 17920 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _170_
timestamp 1698175906
transform 1 0 25088 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _171_
timestamp 1698175906
transform -1 0 26656 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _172_
timestamp 1698175906
transform 1 0 26880 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _173_
timestamp 1698175906
transform 1 0 21840 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _174_
timestamp 1698175906
transform -1 0 23632 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _175_
timestamp 1698175906
transform 1 0 18256 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _176_
timestamp 1698175906
transform 1 0 16016 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _177_
timestamp 1698175906
transform 1 0 15120 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _178_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 15456 0 1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _179_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 15456 0 1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _180_
timestamp 1698175906
transform -1 0 15792 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_2  _181_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18368 0 -1 23520
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _182_
timestamp 1698175906
transform -1 0 14672 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _183_
timestamp 1698175906
transform 1 0 21504 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _184_
timestamp 1698175906
transform -1 0 16016 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _185_
timestamp 1698175906
transform 1 0 14000 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _186_
timestamp 1698175906
transform 1 0 21504 0 1 20384
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _187_
timestamp 1698175906
transform 1 0 25088 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _188_
timestamp 1698175906
transform 1 0 25088 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _189_
timestamp 1698175906
transform 1 0 22736 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _190_
timestamp 1698175906
transform 1 0 22064 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _191_
timestamp 1698175906
transform 1 0 23072 0 -1 25088
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _192_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 23744 0 -1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _193_
timestamp 1698175906
transform 1 0 27776 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _194_
timestamp 1698175906
transform -1 0 27440 0 -1 25088
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _195_
timestamp 1698175906
transform -1 0 20048 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _196_
timestamp 1698175906
transform 1 0 15120 0 -1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _197_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 25312 0 1 21952
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _198_
timestamp 1698175906
transform -1 0 14896 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _199_
timestamp 1698175906
transform -1 0 17024 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _200_
timestamp 1698175906
transform -1 0 16688 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _201_
timestamp 1698175906
transform -1 0 16576 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _202_
timestamp 1698175906
transform -1 0 20048 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _203_
timestamp 1698175906
transform -1 0 19488 0 1 25088
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _204_
timestamp 1698175906
transform -1 0 22176 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _205_
timestamp 1698175906
transform 1 0 20048 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _206_
timestamp 1698175906
transform -1 0 22064 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _207_
timestamp 1698175906
transform 1 0 19264 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _208_
timestamp 1698175906
transform 1 0 17472 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _209_
timestamp 1698175906
transform -1 0 18480 0 -1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _210_
timestamp 1698175906
transform -1 0 16352 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _211_
timestamp 1698175906
transform 1 0 15680 0 1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _212_
timestamp 1698175906
transform -1 0 15456 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _213_
timestamp 1698175906
transform -1 0 16464 0 -1 20384
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _214_
timestamp 1698175906
transform -1 0 14896 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _215_
timestamp 1698175906
transform 1 0 14448 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _216_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 26432 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _217_
timestamp 1698175906
transform 1 0 19152 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _218_
timestamp 1698175906
transform 1 0 26432 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _219_
timestamp 1698175906
transform 1 0 26544 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _220_
timestamp 1698175906
transform 1 0 14336 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _221_
timestamp 1698175906
transform 1 0 11200 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _222_
timestamp 1698175906
transform 1 0 17696 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _223_
timestamp 1698175906
transform 1 0 20048 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _224_
timestamp 1698175906
transform 1 0 25536 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _225_
timestamp 1698175906
transform 1 0 25200 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _226_
timestamp 1698175906
transform 1 0 23632 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _227_
timestamp 1698175906
transform -1 0 12992 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _228_
timestamp 1698175906
transform -1 0 15120 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _229_
timestamp 1698175906
transform -1 0 13776 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _230_
timestamp 1698175906
transform 1 0 21952 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _231_
timestamp 1698175906
transform 1 0 21616 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _232_
timestamp 1698175906
transform 1 0 26656 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _233_
timestamp 1698175906
transform -1 0 15344 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _234_
timestamp 1698175906
transform 1 0 13664 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _235_
timestamp 1698175906
transform 1 0 16352 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _236_
timestamp 1698175906
transform 1 0 19936 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _237_
timestamp 1698175906
transform 1 0 14896 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _238_
timestamp 1698175906
transform 1 0 13328 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _239_
timestamp 1698175906
transform -1 0 14224 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _243_
timestamp 1698175906
transform -1 0 12768 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _244_
timestamp 1698175906
transform 1 0 27440 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _245_
timestamp 1698175906
transform -1 0 14000 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__216__CLK dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 26208 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__217__CLK
timestamp 1698175906
transform 1 0 22624 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__218__CLK
timestamp 1698175906
transform 1 0 26208 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__219__CLK
timestamp 1698175906
transform 1 0 26320 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__220__CLK
timestamp 1698175906
transform 1 0 17808 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__221__CLK
timestamp 1698175906
transform 1 0 15120 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__222__CLK
timestamp 1698175906
transform 1 0 17472 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__223__CLK
timestamp 1698175906
transform 1 0 23520 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__224__CLK
timestamp 1698175906
transform 1 0 29232 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__225__CLK
timestamp 1698175906
transform 1 0 29232 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__226__CLK
timestamp 1698175906
transform 1 0 27664 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__227__CLK
timestamp 1698175906
transform 1 0 12992 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__228__CLK
timestamp 1698175906
transform 1 0 16352 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__229__CLK
timestamp 1698175906
transform 1 0 13776 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__230__CLK
timestamp 1698175906
transform 1 0 25312 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__231__CLK
timestamp 1698175906
transform 1 0 25312 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__232__CLK
timestamp 1698175906
transform 1 0 26432 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__233__CLK
timestamp 1698175906
transform 1 0 15568 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__234__CLK
timestamp 1698175906
transform 1 0 17472 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__235__CLK
timestamp 1698175906
transform 1 0 19600 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__236__CLK
timestamp 1698175906
transform -1 0 23632 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__237__CLK
timestamp 1698175906
transform 1 0 18144 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__238__CLK
timestamp 1698175906
transform -1 0 17248 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__239__CLK
timestamp 1698175906
transform 1 0 14448 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1698175906
transform 1 0 16800 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19152 0 -1 21952
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1698175906
transform -1 0 20944 0 1 20384
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1698175906
transform 1 0 22736 0 1 20384
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1568 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698175906
transform 1 0 5376 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698175906
transform 1 0 9184 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698175906
transform 1 0 12992 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_138 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 16800 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_165 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19824 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_169
timestamp 1698175906
transform 1 0 20272 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_172
timestamp 1698175906
transform 1 0 20608 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_206
timestamp 1698175906
transform 1 0 24416 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_210
timestamp 1698175906
transform 1 0 24864 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_237
timestamp 1698175906
transform 1 0 27888 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_240
timestamp 1698175906
transform 1 0 28224 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_274
timestamp 1698175906
transform 1 0 32032 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_308
timestamp 1698175906
transform 1 0 35840 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_342
timestamp 1698175906
transform 1 0 39648 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_346 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 40096 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_348
timestamp 1698175906
transform 1 0 40320 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1568 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698175906
transform 1 0 8736 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698175906
transform 1 0 9408 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698175906
transform 1 0 16576 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_168
timestamp 1698175906
transform 1 0 20160 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_200 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 23744 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_208
timestamp 1698175906
transform 1 0 24640 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_212
timestamp 1698175906
transform 1 0 25088 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_276
timestamp 1698175906
transform 1 0 32256 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_282
timestamp 1698175906
transform 1 0 32928 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_346
timestamp 1698175906
transform 1 0 40096 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_348
timestamp 1698175906
transform 1 0 40320 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698175906
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698175906
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698175906
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698175906
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_107
timestamp 1698175906
transform 1 0 13328 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_171
timestamp 1698175906
transform 1 0 20496 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_177
timestamp 1698175906
transform 1 0 21168 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_241
timestamp 1698175906
transform 1 0 28336 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698175906
transform 1 0 29008 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698175906
transform 1 0 36176 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_317
timestamp 1698175906
transform 1 0 36848 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698175906
transform 1 0 1568 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698175906
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698175906
transform 1 0 9408 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698175906
transform 1 0 16576 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_142
timestamp 1698175906
transform 1 0 17248 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_206
timestamp 1698175906
transform 1 0 24416 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_212
timestamp 1698175906
transform 1 0 25088 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_276
timestamp 1698175906
transform 1 0 32256 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_282
timestamp 1698175906
transform 1 0 32928 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_346
timestamp 1698175906
transform 1 0 40096 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_348
timestamp 1698175906
transform 1 0 40320 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698175906
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698175906
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698175906
transform 1 0 5488 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698175906
transform 1 0 12656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_107
timestamp 1698175906
transform 1 0 13328 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698175906
transform 1 0 20496 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_177
timestamp 1698175906
transform 1 0 21168 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_241
timestamp 1698175906
transform 1 0 28336 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698175906
transform 1 0 29008 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698175906
transform 1 0 36176 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_317
timestamp 1698175906
transform 1 0 36848 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698175906
transform 1 0 1568 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698175906
transform 1 0 8736 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698175906
transform 1 0 9408 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698175906
transform 1 0 16576 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_142
timestamp 1698175906
transform 1 0 17248 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_206
timestamp 1698175906
transform 1 0 24416 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_212
timestamp 1698175906
transform 1 0 25088 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698175906
transform 1 0 32256 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_282
timestamp 1698175906
transform 1 0 32928 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_346
timestamp 1698175906
transform 1 0 40096 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_348
timestamp 1698175906
transform 1 0 40320 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698175906
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698175906
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698175906
transform 1 0 5488 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698175906
transform 1 0 12656 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_107
timestamp 1698175906
transform 1 0 13328 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_171
timestamp 1698175906
transform 1 0 20496 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_177
timestamp 1698175906
transform 1 0 21168 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_241
timestamp 1698175906
transform 1 0 28336 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_247
timestamp 1698175906
transform 1 0 29008 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_311
timestamp 1698175906
transform 1 0 36176 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_317
timestamp 1698175906
transform 1 0 36848 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698175906
transform 1 0 1568 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698175906
transform 1 0 8736 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_72
timestamp 1698175906
transform 1 0 9408 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698175906
transform 1 0 16576 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_142
timestamp 1698175906
transform 1 0 17248 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_206
timestamp 1698175906
transform 1 0 24416 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_212
timestamp 1698175906
transform 1 0 25088 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_276
timestamp 1698175906
transform 1 0 32256 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_282
timestamp 1698175906
transform 1 0 32928 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_346
timestamp 1698175906
transform 1 0 40096 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_348
timestamp 1698175906
transform 1 0 40320 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698175906
transform 1 0 1568 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698175906
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_37
timestamp 1698175906
transform 1 0 5488 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_101
timestamp 1698175906
transform 1 0 12656 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_107
timestamp 1698175906
transform 1 0 13328 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_171
timestamp 1698175906
transform 1 0 20496 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_177
timestamp 1698175906
transform 1 0 21168 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_241
timestamp 1698175906
transform 1 0 28336 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_247
timestamp 1698175906
transform 1 0 29008 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_311
timestamp 1698175906
transform 1 0 36176 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_317
timestamp 1698175906
transform 1 0 36848 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698175906
transform 1 0 1568 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698175906
transform 1 0 8736 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_72
timestamp 1698175906
transform 1 0 9408 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_136
timestamp 1698175906
transform 1 0 16576 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_142
timestamp 1698175906
transform 1 0 17248 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_206
timestamp 1698175906
transform 1 0 24416 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_212
timestamp 1698175906
transform 1 0 25088 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_276
timestamp 1698175906
transform 1 0 32256 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_282
timestamp 1698175906
transform 1 0 32928 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_346
timestamp 1698175906
transform 1 0 40096 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_348
timestamp 1698175906
transform 1 0 40320 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698175906
transform 1 0 1568 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698175906
transform 1 0 5152 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_37
timestamp 1698175906
transform 1 0 5488 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698175906
transform 1 0 12656 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_107
timestamp 1698175906
transform 1 0 13328 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_171
timestamp 1698175906
transform 1 0 20496 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_177
timestamp 1698175906
transform 1 0 21168 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_241
timestamp 1698175906
transform 1 0 28336 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_247
timestamp 1698175906
transform 1 0 29008 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_311
timestamp 1698175906
transform 1 0 36176 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_317
timestamp 1698175906
transform 1 0 36848 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2
timestamp 1698175906
transform 1 0 1568 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698175906
transform 1 0 8736 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_72
timestamp 1698175906
transform 1 0 9408 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698175906
transform 1 0 16576 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_142
timestamp 1698175906
transform 1 0 17248 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_206
timestamp 1698175906
transform 1 0 24416 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_212
timestamp 1698175906
transform 1 0 25088 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_276
timestamp 1698175906
transform 1 0 32256 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_282
timestamp 1698175906
transform 1 0 32928 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_346
timestamp 1698175906
transform 1 0 40096 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_348
timestamp 1698175906
transform 1 0 40320 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698175906
transform 1 0 1568 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698175906
transform 1 0 5152 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_37
timestamp 1698175906
transform 1 0 5488 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698175906
transform 1 0 12656 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_107 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 13328 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_123
timestamp 1698175906
transform 1 0 15120 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_127
timestamp 1698175906
transform 1 0 15568 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_138
timestamp 1698175906
transform 1 0 16800 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_142
timestamp 1698175906
transform 1 0 17248 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_158
timestamp 1698175906
transform 1 0 19040 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_172
timestamp 1698175906
transform 1 0 20608 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_174
timestamp 1698175906
transform 1 0 20832 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_177
timestamp 1698175906
transform 1 0 21168 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_241
timestamp 1698175906
transform 1 0 28336 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_247
timestamp 1698175906
transform 1 0 29008 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_311
timestamp 1698175906
transform 1 0 36176 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_317
timestamp 1698175906
transform 1 0 36848 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_2
timestamp 1698175906
transform 1 0 1568 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_66
timestamp 1698175906
transform 1 0 8736 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_72
timestamp 1698175906
transform 1 0 9408 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_104
timestamp 1698175906
transform 1 0 12992 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_106
timestamp 1698175906
transform 1 0 13216 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_142
timestamp 1698175906
transform 1 0 17248 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_146
timestamp 1698175906
transform 1 0 17696 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_154
timestamp 1698175906
transform 1 0 18592 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_166
timestamp 1698175906
transform 1 0 19936 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_196
timestamp 1698175906
transform 1 0 23296 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_200
timestamp 1698175906
transform 1 0 23744 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_208
timestamp 1698175906
transform 1 0 24640 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_212
timestamp 1698175906
transform 1 0 25088 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_216
timestamp 1698175906
transform 1 0 25536 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_232
timestamp 1698175906
transform 1 0 27328 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_239
timestamp 1698175906
transform 1 0 28112 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_271
timestamp 1698175906
transform 1 0 31696 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_279
timestamp 1698175906
transform 1 0 32592 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_282
timestamp 1698175906
transform 1 0 32928 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_346
timestamp 1698175906
transform 1 0 40096 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_348
timestamp 1698175906
transform 1 0 40320 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698175906
transform 1 0 1568 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698175906
transform 1 0 5152 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_37
timestamp 1698175906
transform 1 0 5488 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_101
timestamp 1698175906
transform 1 0 12656 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_107
timestamp 1698175906
transform 1 0 13328 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_109
timestamp 1698175906
transform 1 0 13552 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_139
timestamp 1698175906
transform 1 0 16912 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_143
timestamp 1698175906
transform 1 0 17360 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_177
timestamp 1698175906
transform 1 0 21168 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_181
timestamp 1698175906
transform 1 0 21616 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_183
timestamp 1698175906
transform 1 0 21840 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_242
timestamp 1698175906
transform 1 0 28448 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_244
timestamp 1698175906
transform 1 0 28672 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_247
timestamp 1698175906
transform 1 0 29008 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_251
timestamp 1698175906
transform 1 0 29456 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_317
timestamp 1698175906
transform 1 0 36848 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_2
timestamp 1698175906
transform 1 0 1568 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_66
timestamp 1698175906
transform 1 0 8736 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_72
timestamp 1698175906
transform 1 0 9408 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_104
timestamp 1698175906
transform 1 0 12992 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_120
timestamp 1698175906
transform 1 0 14784 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_136
timestamp 1698175906
transform 1 0 16576 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_142
timestamp 1698175906
transform 1 0 17248 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_174
timestamp 1698175906
transform 1 0 20832 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_190
timestamp 1698175906
transform 1 0 22624 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_199
timestamp 1698175906
transform 1 0 23632 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_207
timestamp 1698175906
transform 1 0 24528 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_209
timestamp 1698175906
transform 1 0 24752 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_220
timestamp 1698175906
transform 1 0 25984 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_253
timestamp 1698175906
transform 1 0 29680 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_269
timestamp 1698175906
transform 1 0 31472 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_277
timestamp 1698175906
transform 1 0 32368 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_279
timestamp 1698175906
transform 1 0 32592 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_282
timestamp 1698175906
transform 1 0 32928 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_314
timestamp 1698175906
transform 1 0 36512 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_322
timestamp 1698175906
transform 1 0 37408 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_2
timestamp 1698175906
transform 1 0 1568 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698175906
transform 1 0 5152 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_37
timestamp 1698175906
transform 1 0 5488 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_101
timestamp 1698175906
transform 1 0 12656 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_107
timestamp 1698175906
transform 1 0 13328 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_139
timestamp 1698175906
transform 1 0 16912 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_147
timestamp 1698175906
transform 1 0 17808 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_173
timestamp 1698175906
transform 1 0 20720 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_177
timestamp 1698175906
transform 1 0 21168 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_193
timestamp 1698175906
transform 1 0 22960 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_201
timestamp 1698175906
transform 1 0 23856 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_208
timestamp 1698175906
transform 1 0 24640 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_216
timestamp 1698175906
transform 1 0 25536 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_231
timestamp 1698175906
transform 1 0 27216 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_238
timestamp 1698175906
transform 1 0 28000 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_242
timestamp 1698175906
transform 1 0 28448 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_244
timestamp 1698175906
transform 1 0 28672 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_247
timestamp 1698175906
transform 1 0 29008 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_311
timestamp 1698175906
transform 1 0 36176 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_317
timestamp 1698175906
transform 1 0 36848 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_321
timestamp 1698175906
transform 1 0 37296 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_2
timestamp 1698175906
transform 1 0 1568 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_66
timestamp 1698175906
transform 1 0 8736 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_72
timestamp 1698175906
transform 1 0 9408 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_80
timestamp 1698175906
transform 1 0 10304 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_84
timestamp 1698175906
transform 1 0 10752 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_115
timestamp 1698175906
transform 1 0 14224 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_119
timestamp 1698175906
transform 1 0 14672 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_135
timestamp 1698175906
transform 1 0 16464 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_139
timestamp 1698175906
transform 1 0 16912 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_142
timestamp 1698175906
transform 1 0 17248 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_150
timestamp 1698175906
transform 1 0 18144 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_160
timestamp 1698175906
transform 1 0 19264 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_168
timestamp 1698175906
transform 1 0 20160 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_172
timestamp 1698175906
transform 1 0 20608 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_174
timestamp 1698175906
transform 1 0 20832 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_181
timestamp 1698175906
transform 1 0 21616 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_197
timestamp 1698175906
transform 1 0 23408 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_205
timestamp 1698175906
transform 1 0 24304 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_209
timestamp 1698175906
transform 1 0 24752 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_212
timestamp 1698175906
transform 1 0 25088 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_236
timestamp 1698175906
transform 1 0 27776 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_268
timestamp 1698175906
transform 1 0 31360 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_276
timestamp 1698175906
transform 1 0 32256 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_282
timestamp 1698175906
transform 1 0 32928 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_314
timestamp 1698175906
transform 1 0 36512 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_322
timestamp 1698175906
transform 1 0 37408 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_2
timestamp 1698175906
transform 1 0 1568 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698175906
transform 1 0 5152 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_37
timestamp 1698175906
transform 1 0 5488 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_101
timestamp 1698175906
transform 1 0 12656 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_107
timestamp 1698175906
transform 1 0 13328 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_115
timestamp 1698175906
transform 1 0 14224 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_145
timestamp 1698175906
transform 1 0 17584 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_149
timestamp 1698175906
transform 1 0 18032 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_153
timestamp 1698175906
transform 1 0 18480 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_160
timestamp 1698175906
transform 1 0 19264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_162
timestamp 1698175906
transform 1 0 19488 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_177
timestamp 1698175906
transform 1 0 21168 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_179
timestamp 1698175906
transform 1 0 21392 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_188
timestamp 1698175906
transform 1 0 22400 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_192
timestamp 1698175906
transform 1 0 22848 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_205
timestamp 1698175906
transform 1 0 24304 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_221
timestamp 1698175906
transform 1 0 26096 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_229
timestamp 1698175906
transform 1 0 26992 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_238
timestamp 1698175906
transform 1 0 28000 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_242
timestamp 1698175906
transform 1 0 28448 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_244
timestamp 1698175906
transform 1 0 28672 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_247
timestamp 1698175906
transform 1 0 29008 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_311
timestamp 1698175906
transform 1 0 36176 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_317
timestamp 1698175906
transform 1 0 36848 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_28
timestamp 1698175906
transform 1 0 4480 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_60
timestamp 1698175906
transform 1 0 8064 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_68
timestamp 1698175906
transform 1 0 8960 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_72
timestamp 1698175906
transform 1 0 9408 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_137
timestamp 1698175906
transform 1 0 16688 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_139
timestamp 1698175906
transform 1 0 16912 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_142
timestamp 1698175906
transform 1 0 17248 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_158
timestamp 1698175906
transform 1 0 19040 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_182
timestamp 1698175906
transform 1 0 21728 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_197
timestamp 1698175906
transform 1 0 23408 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_219
timestamp 1698175906
transform 1 0 25872 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_221
timestamp 1698175906
transform 1 0 26096 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_253
timestamp 1698175906
transform 1 0 29680 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_269
timestamp 1698175906
transform 1 0 31472 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_277
timestamp 1698175906
transform 1 0 32368 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_279
timestamp 1698175906
transform 1 0 32592 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_282
timestamp 1698175906
transform 1 0 32928 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_314
timestamp 1698175906
transform 1 0 36512 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_322
timestamp 1698175906
transform 1 0 37408 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_2
timestamp 1698175906
transform 1 0 1568 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698175906
transform 1 0 5152 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_37
timestamp 1698175906
transform 1 0 5488 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_101
timestamp 1698175906
transform 1 0 12656 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_107
timestamp 1698175906
transform 1 0 13328 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_111
timestamp 1698175906
transform 1 0 13776 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_121
timestamp 1698175906
transform 1 0 14896 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_125
timestamp 1698175906
transform 1 0 15344 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_133
timestamp 1698175906
transform 1 0 16240 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_147
timestamp 1698175906
transform 1 0 17808 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_151
timestamp 1698175906
transform 1 0 18256 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_167
timestamp 1698175906
transform 1 0 20048 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_201
timestamp 1698175906
transform 1 0 23856 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_209
timestamp 1698175906
transform 1 0 24752 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_224
timestamp 1698175906
transform 1 0 26432 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_241
timestamp 1698175906
transform 1 0 28336 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_247
timestamp 1698175906
transform 1 0 29008 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_311
timestamp 1698175906
transform 1 0 36176 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_317
timestamp 1698175906
transform 1 0 36848 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_2
timestamp 1698175906
transform 1 0 1568 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_66
timestamp 1698175906
transform 1 0 8736 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_72
timestamp 1698175906
transform 1 0 9408 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_104
timestamp 1698175906
transform 1 0 12992 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_108
timestamp 1698175906
transform 1 0 13440 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_110
timestamp 1698175906
transform 1 0 13664 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_113
timestamp 1698175906
transform 1 0 14000 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_121
timestamp 1698175906
transform 1 0 14896 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_125
timestamp 1698175906
transform 1 0 15344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_127
timestamp 1698175906
transform 1 0 15568 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_135
timestamp 1698175906
transform 1 0 16464 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_139
timestamp 1698175906
transform 1 0 16912 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_142
timestamp 1698175906
transform 1 0 17248 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_146
timestamp 1698175906
transform 1 0 17696 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_175
timestamp 1698175906
transform 1 0 20944 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_206
timestamp 1698175906
transform 1 0 24416 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_212
timestamp 1698175906
transform 1 0 25088 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_214
timestamp 1698175906
transform 1 0 25312 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_221
timestamp 1698175906
transform 1 0 26096 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_254
timestamp 1698175906
transform 1 0 29792 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_270
timestamp 1698175906
transform 1 0 31584 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_278
timestamp 1698175906
transform 1 0 32480 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_282
timestamp 1698175906
transform 1 0 32928 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_346
timestamp 1698175906
transform 1 0 40096 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_348
timestamp 1698175906
transform 1 0 40320 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_2
timestamp 1698175906
transform 1 0 1568 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698175906
transform 1 0 5152 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_37
timestamp 1698175906
transform 1 0 5488 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_101
timestamp 1698175906
transform 1 0 12656 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_107
timestamp 1698175906
transform 1 0 13328 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_177
timestamp 1698175906
transform 1 0 21168 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_179
timestamp 1698175906
transform 1 0 21392 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_187
timestamp 1698175906
transform 1 0 22288 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_241
timestamp 1698175906
transform 1 0 28336 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_247
timestamp 1698175906
transform 1 0 29008 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_311
timestamp 1698175906
transform 1 0 36176 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_317
timestamp 1698175906
transform 1 0 36848 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_321
timestamp 1698175906
transform 1 0 37296 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_28
timestamp 1698175906
transform 1 0 4480 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_60
timestamp 1698175906
transform 1 0 8064 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_68
timestamp 1698175906
transform 1 0 8960 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_72
timestamp 1698175906
transform 1 0 9408 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_80
timestamp 1698175906
transform 1 0 10304 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_111
timestamp 1698175906
transform 1 0 13776 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_137
timestamp 1698175906
transform 1 0 16688 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_139
timestamp 1698175906
transform 1 0 16912 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_142
timestamp 1698175906
transform 1 0 17248 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_144
timestamp 1698175906
transform 1 0 17472 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_209
timestamp 1698175906
transform 1 0 24752 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_235
timestamp 1698175906
transform 1 0 27664 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_267
timestamp 1698175906
transform 1 0 31248 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_275
timestamp 1698175906
transform 1 0 32144 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_279
timestamp 1698175906
transform 1 0 32592 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_282
timestamp 1698175906
transform 1 0 32928 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_346
timestamp 1698175906
transform 1 0 40096 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_348
timestamp 1698175906
transform 1 0 40320 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_28
timestamp 1698175906
transform 1 0 4480 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_32
timestamp 1698175906
transform 1 0 4928 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698175906
transform 1 0 5152 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_37
timestamp 1698175906
transform 1 0 5488 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_69
timestamp 1698175906
transform 1 0 9072 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_73
timestamp 1698175906
transform 1 0 9520 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_104
timestamp 1698175906
transform 1 0 12992 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_113
timestamp 1698175906
transform 1 0 14000 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_115
timestamp 1698175906
transform 1 0 14224 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_135
timestamp 1698175906
transform 1 0 16464 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_137
timestamp 1698175906
transform 1 0 16688 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_172
timestamp 1698175906
transform 1 0 20608 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_174
timestamp 1698175906
transform 1 0 20832 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_214
timestamp 1698175906
transform 1 0 25312 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_247
timestamp 1698175906
transform 1 0 29008 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_251
timestamp 1698175906
transform 1 0 29456 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_317
timestamp 1698175906
transform 1 0 36848 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_28
timestamp 1698175906
transform 1 0 4480 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_60
timestamp 1698175906
transform 1 0 8064 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_68
timestamp 1698175906
transform 1 0 8960 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_72
timestamp 1698175906
transform 1 0 9408 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_88
timestamp 1698175906
transform 1 0 11200 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_102
timestamp 1698175906
transform 1 0 12768 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_106
timestamp 1698175906
transform 1 0 13216 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_122
timestamp 1698175906
transform 1 0 15008 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_128
timestamp 1698175906
transform 1 0 15680 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_136
timestamp 1698175906
transform 1 0 16576 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_142
timestamp 1698175906
transform 1 0 17248 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_177
timestamp 1698175906
transform 1 0 21168 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_181
timestamp 1698175906
transform 1 0 21616 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_207
timestamp 1698175906
transform 1 0 24528 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_209
timestamp 1698175906
transform 1 0 24752 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_218
timestamp 1698175906
transform 1 0 25760 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_255
timestamp 1698175906
transform 1 0 29904 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_271
timestamp 1698175906
transform 1 0 31696 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_279
timestamp 1698175906
transform 1 0 32592 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_282
timestamp 1698175906
transform 1 0 32928 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_314
timestamp 1698175906
transform 1 0 36512 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_322
timestamp 1698175906
transform 1 0 37408 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_28
timestamp 1698175906
transform 1 0 4480 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_32
timestamp 1698175906
transform 1 0 4928 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698175906
transform 1 0 5152 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_37
timestamp 1698175906
transform 1 0 5488 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_101
timestamp 1698175906
transform 1 0 12656 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_107
timestamp 1698175906
transform 1 0 13328 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_111
timestamp 1698175906
transform 1 0 13776 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_113
timestamp 1698175906
transform 1 0 14000 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_129
timestamp 1698175906
transform 1 0 15792 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_145
timestamp 1698175906
transform 1 0 17584 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_147
timestamp 1698175906
transform 1 0 17808 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_160
timestamp 1698175906
transform 1 0 19264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_162
timestamp 1698175906
transform 1 0 19488 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_174
timestamp 1698175906
transform 1 0 20832 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_184
timestamp 1698175906
transform 1 0 21952 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_241
timestamp 1698175906
transform 1 0 28336 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_247
timestamp 1698175906
transform 1 0 29008 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_311
timestamp 1698175906
transform 1 0 36176 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_317
timestamp 1698175906
transform 1 0 36848 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_321
timestamp 1698175906
transform 1 0 37296 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_28
timestamp 1698175906
transform 1 0 4480 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_60
timestamp 1698175906
transform 1 0 8064 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_68
timestamp 1698175906
transform 1 0 8960 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_72
timestamp 1698175906
transform 1 0 9408 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_88
timestamp 1698175906
transform 1 0 11200 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_92
timestamp 1698175906
transform 1 0 11648 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_132
timestamp 1698175906
transform 1 0 16128 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_136
timestamp 1698175906
transform 1 0 16576 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_142
timestamp 1698175906
transform 1 0 17248 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_152
timestamp 1698175906
transform 1 0 18368 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_156
timestamp 1698175906
transform 1 0 18816 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_158
timestamp 1698175906
transform 1 0 19040 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_188
timestamp 1698175906
transform 1 0 22400 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_192
timestamp 1698175906
transform 1 0 22848 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_201
timestamp 1698175906
transform 1 0 23856 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_209
timestamp 1698175906
transform 1 0 24752 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_212
timestamp 1698175906
transform 1 0 25088 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_220
timestamp 1698175906
transform 1 0 25984 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_233
timestamp 1698175906
transform 1 0 27440 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_237
timestamp 1698175906
transform 1 0 27888 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_269
timestamp 1698175906
transform 1 0 31472 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_277
timestamp 1698175906
transform 1 0 32368 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_279
timestamp 1698175906
transform 1 0 32592 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_282
timestamp 1698175906
transform 1 0 32928 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_314
timestamp 1698175906
transform 1 0 36512 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_322
timestamp 1698175906
transform 1 0 37408 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_2
timestamp 1698175906
transform 1 0 1568 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698175906
transform 1 0 5152 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_37
timestamp 1698175906
transform 1 0 5488 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_101
timestamp 1698175906
transform 1 0 12656 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_107
timestamp 1698175906
transform 1 0 13328 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_150
timestamp 1698175906
transform 1 0 18144 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_162
timestamp 1698175906
transform 1 0 19488 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_170
timestamp 1698175906
transform 1 0 20384 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_174
timestamp 1698175906
transform 1 0 20832 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_177
timestamp 1698175906
transform 1 0 21168 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_241
timestamp 1698175906
transform 1 0 28336 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_247
timestamp 1698175906
transform 1 0 29008 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_311
timestamp 1698175906
transform 1 0 36176 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_317
timestamp 1698175906
transform 1 0 36848 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_28
timestamp 1698175906
transform 1 0 4480 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_60
timestamp 1698175906
transform 1 0 8064 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_68
timestamp 1698175906
transform 1 0 8960 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_72
timestamp 1698175906
transform 1 0 9408 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_88
timestamp 1698175906
transform 1 0 11200 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_125
timestamp 1698175906
transform 1 0 15344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_129
timestamp 1698175906
transform 1 0 15792 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_137
timestamp 1698175906
transform 1 0 16688 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_139
timestamp 1698175906
transform 1 0 16912 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_142
timestamp 1698175906
transform 1 0 17248 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_153
timestamp 1698175906
transform 1 0 18480 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_161
timestamp 1698175906
transform 1 0 19376 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_165
timestamp 1698175906
transform 1 0 19824 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_212
timestamp 1698175906
transform 1 0 25088 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_216
timestamp 1698175906
transform 1 0 25536 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_282
timestamp 1698175906
transform 1 0 32928 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_346
timestamp 1698175906
transform 1 0 40096 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_348
timestamp 1698175906
transform 1 0 40320 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_2
timestamp 1698175906
transform 1 0 1568 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698175906
transform 1 0 5152 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_37
timestamp 1698175906
transform 1 0 5488 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_101
timestamp 1698175906
transform 1 0 12656 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_107
timestamp 1698175906
transform 1 0 13328 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_123
timestamp 1698175906
transform 1 0 15120 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_127
timestamp 1698175906
transform 1 0 15568 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_129
timestamp 1698175906
transform 1 0 15792 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_185
timestamp 1698175906
transform 1 0 22064 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_217
timestamp 1698175906
transform 1 0 25648 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_233
timestamp 1698175906
transform 1 0 27440 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_241
timestamp 1698175906
transform 1 0 28336 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_247
timestamp 1698175906
transform 1 0 29008 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_311
timestamp 1698175906
transform 1 0 36176 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_317
timestamp 1698175906
transform 1 0 36848 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_2
timestamp 1698175906
transform 1 0 1568 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_66
timestamp 1698175906
transform 1 0 8736 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_72
timestamp 1698175906
transform 1 0 9408 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_136
timestamp 1698175906
transform 1 0 16576 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_142
timestamp 1698175906
transform 1 0 17248 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_158
timestamp 1698175906
transform 1 0 19040 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_195
timestamp 1698175906
transform 1 0 23184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_199
timestamp 1698175906
transform 1 0 23632 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_207
timestamp 1698175906
transform 1 0 24528 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_209
timestamp 1698175906
transform 1 0 24752 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_212
timestamp 1698175906
transform 1 0 25088 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_276
timestamp 1698175906
transform 1 0 32256 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_282
timestamp 1698175906
transform 1 0 32928 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_346
timestamp 1698175906
transform 1 0 40096 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_348
timestamp 1698175906
transform 1 0 40320 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_2
timestamp 1698175906
transform 1 0 1568 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698175906
transform 1 0 5152 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_37
timestamp 1698175906
transform 1 0 5488 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_101
timestamp 1698175906
transform 1 0 12656 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_107
timestamp 1698175906
transform 1 0 13328 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_171
timestamp 1698175906
transform 1 0 20496 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_177
timestamp 1698175906
transform 1 0 21168 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_181
timestamp 1698175906
transform 1 0 21616 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_186
timestamp 1698175906
transform 1 0 22176 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_218
timestamp 1698175906
transform 1 0 25760 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_234
timestamp 1698175906
transform 1 0 27552 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_242
timestamp 1698175906
transform 1 0 28448 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_244
timestamp 1698175906
transform 1 0 28672 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_247
timestamp 1698175906
transform 1 0 29008 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_311
timestamp 1698175906
transform 1 0 36176 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_317
timestamp 1698175906
transform 1 0 36848 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_2
timestamp 1698175906
transform 1 0 1568 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_66
timestamp 1698175906
transform 1 0 8736 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_72
timestamp 1698175906
transform 1 0 9408 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_136
timestamp 1698175906
transform 1 0 16576 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_142
timestamp 1698175906
transform 1 0 17248 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_206
timestamp 1698175906
transform 1 0 24416 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_212
timestamp 1698175906
transform 1 0 25088 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_276
timestamp 1698175906
transform 1 0 32256 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_282
timestamp 1698175906
transform 1 0 32928 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_346
timestamp 1698175906
transform 1 0 40096 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_348
timestamp 1698175906
transform 1 0 40320 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698175906
transform 1 0 1568 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698175906
transform 1 0 5152 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_37
timestamp 1698175906
transform 1 0 5488 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_101
timestamp 1698175906
transform 1 0 12656 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_107
timestamp 1698175906
transform 1 0 13328 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_171
timestamp 1698175906
transform 1 0 20496 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_177
timestamp 1698175906
transform 1 0 21168 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_241
timestamp 1698175906
transform 1 0 28336 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_247
timestamp 1698175906
transform 1 0 29008 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_311
timestamp 1698175906
transform 1 0 36176 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_317
timestamp 1698175906
transform 1 0 36848 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2
timestamp 1698175906
transform 1 0 1568 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_66
timestamp 1698175906
transform 1 0 8736 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_72
timestamp 1698175906
transform 1 0 9408 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_136
timestamp 1698175906
transform 1 0 16576 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_142
timestamp 1698175906
transform 1 0 17248 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_206
timestamp 1698175906
transform 1 0 24416 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_212
timestamp 1698175906
transform 1 0 25088 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_276
timestamp 1698175906
transform 1 0 32256 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_282
timestamp 1698175906
transform 1 0 32928 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_346
timestamp 1698175906
transform 1 0 40096 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_348
timestamp 1698175906
transform 1 0 40320 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_2
timestamp 1698175906
transform 1 0 1568 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698175906
transform 1 0 5152 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_37
timestamp 1698175906
transform 1 0 5488 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_101
timestamp 1698175906
transform 1 0 12656 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_107
timestamp 1698175906
transform 1 0 13328 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_171
timestamp 1698175906
transform 1 0 20496 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_177
timestamp 1698175906
transform 1 0 21168 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_241
timestamp 1698175906
transform 1 0 28336 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_247
timestamp 1698175906
transform 1 0 29008 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_311
timestamp 1698175906
transform 1 0 36176 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_317
timestamp 1698175906
transform 1 0 36848 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2
timestamp 1698175906
transform 1 0 1568 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_66
timestamp 1698175906
transform 1 0 8736 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_72
timestamp 1698175906
transform 1 0 9408 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_136
timestamp 1698175906
transform 1 0 16576 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_142
timestamp 1698175906
transform 1 0 17248 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_206
timestamp 1698175906
transform 1 0 24416 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_212
timestamp 1698175906
transform 1 0 25088 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_276
timestamp 1698175906
transform 1 0 32256 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_282
timestamp 1698175906
transform 1 0 32928 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_346
timestamp 1698175906
transform 1 0 40096 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_348
timestamp 1698175906
transform 1 0 40320 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698175906
transform 1 0 1568 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698175906
transform 1 0 5152 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_37
timestamp 1698175906
transform 1 0 5488 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_101
timestamp 1698175906
transform 1 0 12656 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_107
timestamp 1698175906
transform 1 0 13328 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_171
timestamp 1698175906
transform 1 0 20496 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_177
timestamp 1698175906
transform 1 0 21168 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_241
timestamp 1698175906
transform 1 0 28336 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_247
timestamp 1698175906
transform 1 0 29008 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_311
timestamp 1698175906
transform 1 0 36176 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_317
timestamp 1698175906
transform 1 0 36848 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_2
timestamp 1698175906
transform 1 0 1568 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_66
timestamp 1698175906
transform 1 0 8736 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_72
timestamp 1698175906
transform 1 0 9408 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_136
timestamp 1698175906
transform 1 0 16576 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_142
timestamp 1698175906
transform 1 0 17248 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_206
timestamp 1698175906
transform 1 0 24416 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_212
timestamp 1698175906
transform 1 0 25088 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_276
timestamp 1698175906
transform 1 0 32256 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_282
timestamp 1698175906
transform 1 0 32928 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_346
timestamp 1698175906
transform 1 0 40096 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_348
timestamp 1698175906
transform 1 0 40320 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698175906
transform 1 0 1568 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698175906
transform 1 0 5152 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_37
timestamp 1698175906
transform 1 0 5488 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_101
timestamp 1698175906
transform 1 0 12656 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_107
timestamp 1698175906
transform 1 0 13328 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_171
timestamp 1698175906
transform 1 0 20496 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_177
timestamp 1698175906
transform 1 0 21168 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_241
timestamp 1698175906
transform 1 0 28336 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_247
timestamp 1698175906
transform 1 0 29008 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_311
timestamp 1698175906
transform 1 0 36176 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_317
timestamp 1698175906
transform 1 0 36848 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2
timestamp 1698175906
transform 1 0 1568 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1698175906
transform 1 0 8736 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_72
timestamp 1698175906
transform 1 0 9408 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_136
timestamp 1698175906
transform 1 0 16576 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_142
timestamp 1698175906
transform 1 0 17248 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_206
timestamp 1698175906
transform 1 0 24416 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_212
timestamp 1698175906
transform 1 0 25088 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_276
timestamp 1698175906
transform 1 0 32256 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_282
timestamp 1698175906
transform 1 0 32928 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_346
timestamp 1698175906
transform 1 0 40096 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_348
timestamp 1698175906
transform 1 0 40320 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_6
timestamp 1698175906
transform 1 0 2016 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_22
timestamp 1698175906
transform 1 0 3808 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_30
timestamp 1698175906
transform 1 0 4704 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698175906
transform 1 0 5152 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_37
timestamp 1698175906
transform 1 0 5488 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_101
timestamp 1698175906
transform 1 0 12656 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_107
timestamp 1698175906
transform 1 0 13328 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_171
timestamp 1698175906
transform 1 0 20496 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_177
timestamp 1698175906
transform 1 0 21168 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_241
timestamp 1698175906
transform 1 0 28336 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_247
timestamp 1698175906
transform 1 0 29008 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_311
timestamp 1698175906
transform 1 0 36176 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_317
timestamp 1698175906
transform 1 0 36848 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_2
timestamp 1698175906
transform 1 0 1568 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_66
timestamp 1698175906
transform 1 0 8736 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_72
timestamp 1698175906
transform 1 0 9408 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_136
timestamp 1698175906
transform 1 0 16576 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_142
timestamp 1698175906
transform 1 0 17248 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_150
timestamp 1698175906
transform 1 0 18144 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_155
timestamp 1698175906
transform 1 0 18704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_183
timestamp 1698175906
transform 1 0 21840 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_199
timestamp 1698175906
transform 1 0 23632 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_207
timestamp 1698175906
transform 1 0 24528 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_209
timestamp 1698175906
transform 1 0 24752 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_238
timestamp 1698175906
transform 1 0 28000 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_270
timestamp 1698175906
transform 1 0 31584 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_278
timestamp 1698175906
transform 1 0 32480 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_282
timestamp 1698175906
transform 1 0 32928 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_346
timestamp 1698175906
transform 1 0 40096 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_348
timestamp 1698175906
transform 1 0 40320 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_2
timestamp 1698175906
transform 1 0 1568 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_36
timestamp 1698175906
transform 1 0 5376 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_70
timestamp 1698175906
transform 1 0 9184 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_104
timestamp 1698175906
transform 1 0 12992 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_138
timestamp 1698175906
transform 1 0 16800 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_142
timestamp 1698175906
transform 1 0 17248 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_172
timestamp 1698175906
transform 1 0 20608 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_176
timestamp 1698175906
transform 1 0 21056 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_236
timestamp 1698175906
transform 1 0 27776 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_240
timestamp 1698175906
transform 1 0 28224 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_274
timestamp 1698175906
transform 1 0 32032 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_308
timestamp 1698175906
transform 1 0 35840 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_342
timestamp 1698175906
transform 1 0 39648 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_346
timestamp 1698175906
transform 1 0 40096 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_348
timestamp 1698175906
transform 1 0 40320 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita28_24 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 27776 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita28_25
timestamp 1698175906
transform -1 0 2016 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita28_26
timestamp 1698175906
transform -1 0 18704 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 4480 0 1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output2
timestamp 1698175906
transform 1 0 24976 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output3
timestamp 1698175906
transform 1 0 17472 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output4
timestamp 1698175906
transform 1 0 25088 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output5
timestamp 1698175906
transform 1 0 37520 0 1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output6
timestamp 1698175906
transform 1 0 37520 0 1 15680
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output7
timestamp 1698175906
transform -1 0 4480 0 1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output8
timestamp 1698175906
transform -1 0 4480 0 -1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output9
timestamp 1698175906
transform 1 0 18928 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output10
timestamp 1698175906
transform -1 0 4480 0 -1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output11
timestamp 1698175906
transform 1 0 24416 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output12
timestamp 1698175906
transform 1 0 37520 0 -1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output13
timestamp 1698175906
transform -1 0 4480 0 -1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output14
timestamp 1698175906
transform 1 0 16912 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output15
timestamp 1698175906
transform 1 0 37520 0 -1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output16
timestamp 1698175906
transform 1 0 37520 0 1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output17
timestamp 1698175906
transform 1 0 37520 0 -1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output18
timestamp 1698175906
transform 1 0 37520 0 -1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output19
timestamp 1698175906
transform 1 0 21280 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output20
timestamp 1698175906
transform 1 0 37520 0 -1 15680
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output21
timestamp 1698175906
transform 1 0 17248 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output22
timestamp 1698175906
transform -1 0 4480 0 -1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output23
timestamp 1698175906
transform -1 0 4480 0 -1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_45 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698175906
transform -1 0 40656 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_46
timestamp 1698175906
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698175906
transform -1 0 40656 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_47
timestamp 1698175906
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698175906
transform -1 0 40656 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_48
timestamp 1698175906
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698175906
transform -1 0 40656 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_49
timestamp 1698175906
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698175906
transform -1 0 40656 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_50
timestamp 1698175906
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698175906
transform -1 0 40656 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_51
timestamp 1698175906
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698175906
transform -1 0 40656 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_52
timestamp 1698175906
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698175906
transform -1 0 40656 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_53
timestamp 1698175906
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698175906
transform -1 0 40656 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_54
timestamp 1698175906
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698175906
transform -1 0 40656 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_55
timestamp 1698175906
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698175906
transform -1 0 40656 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_56
timestamp 1698175906
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698175906
transform -1 0 40656 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_57
timestamp 1698175906
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698175906
transform -1 0 40656 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_58
timestamp 1698175906
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698175906
transform -1 0 40656 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_59
timestamp 1698175906
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698175906
transform -1 0 40656 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_60
timestamp 1698175906
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698175906
transform -1 0 40656 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_61
timestamp 1698175906
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698175906
transform -1 0 40656 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_62
timestamp 1698175906
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698175906
transform -1 0 40656 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_63
timestamp 1698175906
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698175906
transform -1 0 40656 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_64
timestamp 1698175906
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698175906
transform -1 0 40656 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_65
timestamp 1698175906
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698175906
transform -1 0 40656 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_66
timestamp 1698175906
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698175906
transform -1 0 40656 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_67
timestamp 1698175906
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698175906
transform -1 0 40656 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_68
timestamp 1698175906
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698175906
transform -1 0 40656 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_69
timestamp 1698175906
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698175906
transform -1 0 40656 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_70
timestamp 1698175906
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698175906
transform -1 0 40656 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_71
timestamp 1698175906
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698175906
transform -1 0 40656 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_72
timestamp 1698175906
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698175906
transform -1 0 40656 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_73
timestamp 1698175906
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698175906
transform -1 0 40656 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_74
timestamp 1698175906
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698175906
transform -1 0 40656 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_75
timestamp 1698175906
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698175906
transform -1 0 40656 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_76
timestamp 1698175906
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698175906
transform -1 0 40656 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_77
timestamp 1698175906
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698175906
transform -1 0 40656 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_78
timestamp 1698175906
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698175906
transform -1 0 40656 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_79
timestamp 1698175906
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698175906
transform -1 0 40656 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_80
timestamp 1698175906
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698175906
transform -1 0 40656 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_81
timestamp 1698175906
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698175906
transform -1 0 40656 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_82
timestamp 1698175906
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698175906
transform -1 0 40656 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_83
timestamp 1698175906
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698175906
transform -1 0 40656 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_84
timestamp 1698175906
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698175906
transform -1 0 40656 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_85
timestamp 1698175906
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698175906
transform -1 0 40656 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_86
timestamp 1698175906
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698175906
transform -1 0 40656 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_87
timestamp 1698175906
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698175906
transform -1 0 40656 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_88
timestamp 1698175906
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698175906
transform -1 0 40656 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_89
timestamp 1698175906
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698175906
transform -1 0 40656 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_90 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_91
timestamp 1698175906
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_92
timestamp 1698175906
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_93
timestamp 1698175906
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_94
timestamp 1698175906
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_95
timestamp 1698175906
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_96
timestamp 1698175906
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_97
timestamp 1698175906
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_98
timestamp 1698175906
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_99
timestamp 1698175906
transform 1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_100
timestamp 1698175906
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_101
timestamp 1698175906
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_102
timestamp 1698175906
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_103
timestamp 1698175906
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_104
timestamp 1698175906
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_105
timestamp 1698175906
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_106
timestamp 1698175906
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_107
timestamp 1698175906
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_108
timestamp 1698175906
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_109
timestamp 1698175906
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_110
timestamp 1698175906
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_111
timestamp 1698175906
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_112
timestamp 1698175906
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_113
timestamp 1698175906
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_114
timestamp 1698175906
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_115
timestamp 1698175906
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_116
timestamp 1698175906
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_117
timestamp 1698175906
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_118
timestamp 1698175906
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_119
timestamp 1698175906
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_120
timestamp 1698175906
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_121
timestamp 1698175906
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_122
timestamp 1698175906
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_123
timestamp 1698175906
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_124
timestamp 1698175906
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_125
timestamp 1698175906
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_126
timestamp 1698175906
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_127
timestamp 1698175906
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_128
timestamp 1698175906
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_129
timestamp 1698175906
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_130
timestamp 1698175906
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_131
timestamp 1698175906
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_132
timestamp 1698175906
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_133
timestamp 1698175906
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_134
timestamp 1698175906
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_135
timestamp 1698175906
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_136
timestamp 1698175906
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_137
timestamp 1698175906
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_138
timestamp 1698175906
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_139
timestamp 1698175906
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_140
timestamp 1698175906
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_141
timestamp 1698175906
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_142
timestamp 1698175906
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_143
timestamp 1698175906
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_144
timestamp 1698175906
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_145
timestamp 1698175906
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_146
timestamp 1698175906
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_147
timestamp 1698175906
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_148
timestamp 1698175906
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_149
timestamp 1698175906
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_150
timestamp 1698175906
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_151
timestamp 1698175906
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_152
timestamp 1698175906
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_153
timestamp 1698175906
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_154
timestamp 1698175906
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_155
timestamp 1698175906
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_156
timestamp 1698175906
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_157
timestamp 1698175906
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_158
timestamp 1698175906
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_159
timestamp 1698175906
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_160
timestamp 1698175906
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_161
timestamp 1698175906
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_162
timestamp 1698175906
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_163
timestamp 1698175906
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_164
timestamp 1698175906
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_165
timestamp 1698175906
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_166
timestamp 1698175906
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_167
timestamp 1698175906
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_168
timestamp 1698175906
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_169
timestamp 1698175906
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_170
timestamp 1698175906
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_171
timestamp 1698175906
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_172
timestamp 1698175906
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_173
timestamp 1698175906
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_174
timestamp 1698175906
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_175
timestamp 1698175906
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_176
timestamp 1698175906
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_177
timestamp 1698175906
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_178
timestamp 1698175906
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_179
timestamp 1698175906
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_180
timestamp 1698175906
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_181
timestamp 1698175906
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_182
timestamp 1698175906
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_183
timestamp 1698175906
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_184
timestamp 1698175906
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_185
timestamp 1698175906
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_186
timestamp 1698175906
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_187
timestamp 1698175906
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_188
timestamp 1698175906
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_189
timestamp 1698175906
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_190
timestamp 1698175906
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_191
timestamp 1698175906
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_192
timestamp 1698175906
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_193
timestamp 1698175906
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_194
timestamp 1698175906
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_195
timestamp 1698175906
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_196
timestamp 1698175906
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_197
timestamp 1698175906
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_198
timestamp 1698175906
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_199
timestamp 1698175906
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_200
timestamp 1698175906
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_201
timestamp 1698175906
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_202
timestamp 1698175906
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_203
timestamp 1698175906
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_204
timestamp 1698175906
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_205
timestamp 1698175906
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_206
timestamp 1698175906
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_207
timestamp 1698175906
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_208
timestamp 1698175906
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_209
timestamp 1698175906
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_210
timestamp 1698175906
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_211
timestamp 1698175906
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_212
timestamp 1698175906
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_213
timestamp 1698175906
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_214
timestamp 1698175906
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_215
timestamp 1698175906
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_216
timestamp 1698175906
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_217
timestamp 1698175906
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_218
timestamp 1698175906
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_219
timestamp 1698175906
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_220
timestamp 1698175906
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_221
timestamp 1698175906
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_222
timestamp 1698175906
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_223
timestamp 1698175906
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_224
timestamp 1698175906
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_225
timestamp 1698175906
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_226
timestamp 1698175906
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_227
timestamp 1698175906
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_228
timestamp 1698175906
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_229
timestamp 1698175906
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_230
timestamp 1698175906
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_231
timestamp 1698175906
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_232
timestamp 1698175906
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_233
timestamp 1698175906
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_234
timestamp 1698175906
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_235
timestamp 1698175906
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_236
timestamp 1698175906
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_237
timestamp 1698175906
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_238
timestamp 1698175906
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_239
timestamp 1698175906
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_240
timestamp 1698175906
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_241
timestamp 1698175906
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_242
timestamp 1698175906
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_243
timestamp 1698175906
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_244
timestamp 1698175906
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_245
timestamp 1698175906
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_246
timestamp 1698175906
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_247
timestamp 1698175906
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_248
timestamp 1698175906
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_249
timestamp 1698175906
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_250
timestamp 1698175906
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_251
timestamp 1698175906
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_252
timestamp 1698175906
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_253
timestamp 1698175906
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_254
timestamp 1698175906
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_255
timestamp 1698175906
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_256
timestamp 1698175906
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_257
timestamp 1698175906
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_258
timestamp 1698175906
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_259
timestamp 1698175906
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_260
timestamp 1698175906
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_261
timestamp 1698175906
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_262
timestamp 1698175906
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_263
timestamp 1698175906
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_264
timestamp 1698175906
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_265
timestamp 1698175906
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_266
timestamp 1698175906
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_267
timestamp 1698175906
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_268
timestamp 1698175906
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_269
timestamp 1698175906
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_270
timestamp 1698175906
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_271
timestamp 1698175906
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_272
timestamp 1698175906
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_273
timestamp 1698175906
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_274
timestamp 1698175906
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_275
timestamp 1698175906
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_276
timestamp 1698175906
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_277
timestamp 1698175906
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_278
timestamp 1698175906
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_279
timestamp 1698175906
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_280
timestamp 1698175906
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_281
timestamp 1698175906
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_282
timestamp 1698175906
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_283
timestamp 1698175906
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_284
timestamp 1698175906
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_285
timestamp 1698175906
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_286
timestamp 1698175906
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_287
timestamp 1698175906
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_288
timestamp 1698175906
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_289
timestamp 1698175906
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_290
timestamp 1698175906
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_291
timestamp 1698175906
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_292
timestamp 1698175906
transform 1 0 32704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_293
timestamp 1698175906
transform 1 0 5152 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_294
timestamp 1698175906
transform 1 0 8960 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_295
timestamp 1698175906
transform 1 0 12768 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_296
timestamp 1698175906
transform 1 0 16576 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_297
timestamp 1698175906
transform 1 0 20384 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_298
timestamp 1698175906
transform 1 0 24192 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_299
timestamp 1698175906
transform 1 0 28000 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_300
timestamp 1698175906
transform 1 0 31808 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_301
timestamp 1698175906
transform 1 0 35616 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_302
timestamp 1698175906
transform 1 0 39424 0 1 37632
box -86 -86 310 870
<< labels >>
flabel metal3 s 0 28224 800 28336 0 FreeSans 448 0 0 0 clk
port 0 nsew signal input
flabel metal3 s 0 23520 800 23632 0 FreeSans 448 0 0 0 segm[0]
port 1 nsew signal tristate
flabel metal2 s 24864 0 24976 800 0 FreeSans 448 90 0 0 segm[10]
port 2 nsew signal tristate
flabel metal2 s 17472 41200 17584 42000 0 FreeSans 448 90 0 0 segm[11]
port 3 nsew signal tristate
flabel metal2 s 24864 41200 24976 42000 0 FreeSans 448 90 0 0 segm[12]
port 4 nsew signal tristate
flabel metal3 s 41200 23520 42000 23632 0 FreeSans 448 0 0 0 segm[13]
port 5 nsew signal tristate
flabel metal2 s 26880 41200 26992 42000 0 FreeSans 448 90 0 0 segm[1]
port 6 nsew signal tristate
flabel metal3 s 41200 15456 42000 15568 0 FreeSans 448 0 0 0 segm[2]
port 7 nsew signal tristate
flabel metal3 s 0 22176 800 22288 0 FreeSans 448 0 0 0 segm[3]
port 8 nsew signal tristate
flabel metal3 s 0 36288 800 36400 0 FreeSans 448 0 0 0 segm[4]
port 9 nsew signal tristate
flabel metal2 s 18144 41200 18256 42000 0 FreeSans 448 90 0 0 segm[5]
port 10 nsew signal tristate
flabel metal3 s 0 24192 800 24304 0 FreeSans 448 0 0 0 segm[6]
port 11 nsew signal tristate
flabel metal2 s 18816 41200 18928 42000 0 FreeSans 448 90 0 0 segm[7]
port 12 nsew signal tristate
flabel metal3 s 0 21504 800 21616 0 FreeSans 448 0 0 0 segm[8]
port 13 nsew signal tristate
flabel metal2 s 22848 41200 22960 42000 0 FreeSans 448 90 0 0 segm[9]
port 14 nsew signal tristate
flabel metal3 s 41200 24192 42000 24304 0 FreeSans 448 0 0 0 sel[0]
port 15 nsew signal tristate
flabel metal3 s 0 25536 800 25648 0 FreeSans 448 0 0 0 sel[10]
port 16 nsew signal tristate
flabel metal2 s 16800 0 16912 800 0 FreeSans 448 90 0 0 sel[11]
port 17 nsew signal tristate
flabel metal3 s 41200 22848 42000 22960 0 FreeSans 448 0 0 0 sel[1]
port 18 nsew signal tristate
flabel metal3 s 41200 20160 42000 20272 0 FreeSans 448 0 0 0 sel[2]
port 19 nsew signal tristate
flabel metal3 s 41200 18144 42000 18256 0 FreeSans 448 0 0 0 sel[3]
port 20 nsew signal tristate
flabel metal3 s 41200 16128 42000 16240 0 FreeSans 448 0 0 0 sel[4]
port 21 nsew signal tristate
flabel metal2 s 22176 41200 22288 42000 0 FreeSans 448 90 0 0 sel[5]
port 22 nsew signal tristate
flabel metal3 s 41200 14784 42000 14896 0 FreeSans 448 0 0 0 sel[6]
port 23 nsew signal tristate
flabel metal2 s 16128 0 16240 800 0 FreeSans 448 90 0 0 sel[7]
port 24 nsew signal tristate
flabel metal3 s 0 18144 800 18256 0 FreeSans 448 0 0 0 sel[8]
port 25 nsew signal tristate
flabel metal3 s 0 22848 800 22960 0 FreeSans 448 0 0 0 sel[9]
port 26 nsew signal tristate
flabel metal4 s 4448 3076 4768 38476 0 FreeSans 1280 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 35168 3076 35488 38476 0 FreeSans 1280 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 19808 3076 20128 38476 0 FreeSans 1280 90 0 0 vss
port 28 nsew ground bidirectional
rlabel metal1 21000 38416 21000 38416 0 vdd
rlabel metal1 21000 37632 21000 37632 0 vss
rlabel metal2 26264 15848 26264 15848 0 _000_
rlabel metal3 23968 23800 23968 23800 0 _001_
rlabel metal3 14000 22232 14000 22232 0 _002_
rlabel metal2 14168 24248 14168 24248 0 _003_
rlabel metal3 13552 21448 13552 21448 0 _004_
rlabel metal2 22960 14616 22960 14616 0 _005_
rlabel metal3 22792 23576 22792 23576 0 _006_
rlabel metal2 27552 23240 27552 23240 0 _007_
rlabel metal2 14392 25928 14392 25928 0 _008_
rlabel metal2 14616 15064 14616 15064 0 _009_
rlabel metal3 17920 25592 17920 25592 0 _010_
rlabel metal3 20328 27944 20328 27944 0 _011_
rlabel metal2 16072 26208 16072 26208 0 _012_
rlabel metal2 14280 14504 14280 14504 0 _013_
rlabel metal2 13272 17640 13272 17640 0 _014_
rlabel metal2 27384 16240 27384 16240 0 _015_
rlabel metal2 19880 24304 19880 24304 0 _016_
rlabel metal2 27384 18592 27384 18592 0 _017_
rlabel metal2 27496 19600 27496 19600 0 _018_
rlabel metal2 14448 20328 14448 20328 0 _019_
rlabel metal2 12152 19264 12152 19264 0 _020_
rlabel metal2 18648 14840 18648 14840 0 _021_
rlabel metal2 20440 13216 20440 13216 0 _022_
rlabel metal2 26488 22008 26488 22008 0 _023_
rlabel metal2 19432 14056 19432 14056 0 _024_
rlabel metal2 20104 13216 20104 13216 0 _025_
rlabel metal2 26264 22064 26264 22064 0 _026_
rlabel metal2 27160 21168 27160 21168 0 _027_
rlabel metal3 26824 21560 26824 21560 0 _028_
rlabel metal2 26152 17136 26152 17136 0 _029_
rlabel metal2 26656 15960 26656 15960 0 _030_
rlabel metal2 23240 23744 23240 23744 0 _031_
rlabel metal2 27048 23408 27048 23408 0 _032_
rlabel metal2 27608 23688 27608 23688 0 _033_
rlabel metal3 27020 24024 27020 24024 0 _034_
rlabel metal3 20496 24136 20496 24136 0 _035_
rlabel metal2 22232 23660 22232 23660 0 _036_
rlabel metal2 15792 21672 15792 21672 0 _037_
rlabel metal2 15848 22736 15848 22736 0 _038_
rlabel metal2 15624 22400 15624 22400 0 _039_
rlabel metal2 14392 23912 14392 23912 0 _040_
rlabel metal2 14504 23576 14504 23576 0 _041_
rlabel metal2 21952 20776 21952 20776 0 _042_
rlabel metal2 14728 21728 14728 21728 0 _043_
rlabel metal2 23128 22680 23128 22680 0 _044_
rlabel metal2 22904 16128 22904 16128 0 _045_
rlabel metal3 24416 15288 24416 15288 0 _046_
rlabel metal2 22344 23604 22344 23604 0 _047_
rlabel metal2 23576 23912 23576 23912 0 _048_
rlabel metal2 28056 24192 28056 24192 0 _049_
rlabel metal2 18984 24696 18984 24696 0 _050_
rlabel metal2 14504 25088 14504 25088 0 _051_
rlabel metal3 14924 25368 14924 25368 0 _052_
rlabel metal2 16744 14168 16744 14168 0 _053_
rlabel metal2 15848 14112 15848 14112 0 _054_
rlabel metal2 19656 26824 19656 26824 0 _055_
rlabel metal2 20552 27776 20552 27776 0 _056_
rlabel metal2 20328 27328 20328 27328 0 _057_
rlabel metal3 21336 27160 21336 27160 0 _058_
rlabel metal2 17752 24080 17752 24080 0 _059_
rlabel metal3 17080 26488 17080 26488 0 _060_
rlabel metal2 15624 12600 15624 12600 0 _061_
rlabel metal2 14952 19096 14952 19096 0 _062_
rlabel metal2 14616 18760 14616 18760 0 _063_
rlabel metal2 25928 18816 25928 18816 0 _064_
rlabel metal2 27944 23520 27944 23520 0 _065_
rlabel metal2 22904 18816 22904 18816 0 _066_
rlabel metal2 23800 16744 23800 16744 0 _067_
rlabel metal2 27608 16800 27608 16800 0 _068_
rlabel metal2 27720 16576 27720 16576 0 _069_
rlabel metal2 19656 18760 19656 18760 0 _070_
rlabel metal3 17136 19992 17136 19992 0 _071_
rlabel metal2 27160 16408 27160 16408 0 _072_
rlabel metal2 21448 17752 21448 17752 0 _073_
rlabel metal2 25144 22680 25144 22680 0 _074_
rlabel metal3 15960 12824 15960 12824 0 _075_
rlabel metal2 20552 21224 20552 21224 0 _076_
rlabel metal2 26040 19880 26040 19880 0 _077_
rlabel metal2 21896 18424 21896 18424 0 _078_
rlabel metal3 18200 20104 18200 20104 0 _079_
rlabel metal2 19320 17976 19320 17976 0 _080_
rlabel metal2 20160 22344 20160 22344 0 _081_
rlabel metal2 20440 23968 20440 23968 0 _082_
rlabel metal2 22456 19768 22456 19768 0 _083_
rlabel metal3 20664 22232 20664 22232 0 _084_
rlabel metal2 20496 22568 20496 22568 0 _085_
rlabel metal3 18200 22120 18200 22120 0 _086_
rlabel metal2 14504 21784 14504 21784 0 _087_
rlabel metal2 17976 22344 17976 22344 0 _088_
rlabel metal2 22344 23128 22344 23128 0 _089_
rlabel metal2 15064 20048 15064 20048 0 _090_
rlabel metal2 24136 22176 24136 22176 0 _091_
rlabel metal2 23128 19992 23128 19992 0 _092_
rlabel metal2 23800 21672 23800 21672 0 _093_
rlabel metal2 27832 20664 27832 20664 0 _094_
rlabel metal2 28000 17640 28000 17640 0 _095_
rlabel metal2 27160 19096 27160 19096 0 _096_
rlabel metal2 27048 19488 27048 19488 0 _097_
rlabel metal2 25592 19824 25592 19824 0 _098_
rlabel metal3 26152 19208 26152 19208 0 _099_
rlabel metal2 14728 20664 14728 20664 0 _100_
rlabel metal2 13832 20496 13832 20496 0 _101_
rlabel metal2 17976 19992 17976 19992 0 _102_
rlabel metal2 14168 22232 14168 22232 0 _103_
rlabel metal2 19152 16072 19152 16072 0 _104_
rlabel metal2 19544 15624 19544 15624 0 _105_
rlabel metal2 20384 14840 20384 14840 0 _106_
rlabel metal2 14952 22400 14952 22400 0 _107_
rlabel metal3 2478 28280 2478 28280 0 clk
rlabel metal2 22904 21112 22904 21112 0 clknet_0_clk
rlabel metal2 14952 24640 14952 24640 0 clknet_1_0__leaf_clk
rlabel metal3 21000 27832 21000 27832 0 clknet_1_1__leaf_clk
rlabel metal2 22456 18760 22456 18760 0 dut28.count\[0\]
rlabel metal2 14280 18256 14280 18256 0 dut28.count\[1\]
rlabel metal2 21112 17248 21112 17248 0 dut28.count\[2\]
rlabel metal2 23184 13608 23184 13608 0 dut28.count\[3\]
rlabel metal2 12264 23632 12264 23632 0 net1
rlabel metal3 6356 21560 6356 21560 0 net10
rlabel metal2 23016 28224 23016 28224 0 net11
rlabel metal2 37912 24248 37912 24248 0 net12
rlabel metal2 12264 26208 12264 26208 0 net13
rlabel metal2 17080 5964 17080 5964 0 net14
rlabel metal2 28616 22512 28616 22512 0 net15
rlabel metal2 29624 19488 29624 19488 0 net16
rlabel metal2 27720 17920 27720 17920 0 net17
rlabel metal2 27720 15512 27720 15512 0 net18
rlabel metal3 21896 24584 21896 24584 0 net19
rlabel metal2 25144 14616 25144 14616 0 net2
rlabel metal2 37688 14560 37688 14560 0 net20
rlabel metal2 16072 12152 16072 12152 0 net21
rlabel metal3 6356 18424 6356 18424 0 net22
rlabel metal2 4312 23072 4312 23072 0 net23
rlabel metal2 27496 38248 27496 38248 0 net24
rlabel metal3 1246 36344 1246 36344 0 net25
rlabel metal2 18312 37464 18312 37464 0 net26
rlabel metal2 17920 25592 17920 25592 0 net3
rlabel metal2 25256 32060 25256 32060 0 net4
rlabel metal2 29736 23464 29736 23464 0 net5
rlabel metal2 28280 15176 28280 15176 0 net6
rlabel metal2 9912 22400 9912 22400 0 net7
rlabel metal2 12040 24640 12040 24640 0 net8
rlabel metal2 19656 27160 19656 27160 0 net9
rlabel metal3 1358 23576 1358 23576 0 segm[0]
rlabel metal2 24920 2198 24920 2198 0 segm[10]
rlabel metal2 17528 39746 17528 39746 0 segm[11]
rlabel metal2 24920 39354 24920 39354 0 segm[12]
rlabel metal2 40040 23800 40040 23800 0 segm[13]
rlabel metal2 40040 15848 40040 15848 0 segm[2]
rlabel metal3 1358 22232 1358 22232 0 segm[3]
rlabel metal3 1358 24248 1358 24248 0 segm[6]
rlabel metal3 19488 37464 19488 37464 0 segm[7]
rlabel metal3 1358 21560 1358 21560 0 segm[8]
rlabel metal2 22904 39746 22904 39746 0 segm[9]
rlabel metal2 40040 24360 40040 24360 0 sel[0]
rlabel metal3 1358 25592 1358 25592 0 sel[10]
rlabel metal2 16856 2086 16856 2086 0 sel[11]
rlabel metal3 40642 22904 40642 22904 0 sel[1]
rlabel metal2 40040 20552 40040 20552 0 sel[2]
rlabel metal3 40642 18200 40642 18200 0 sel[3]
rlabel metal2 39928 16464 39928 16464 0 sel[4]
rlabel metal2 22232 39746 22232 39746 0 sel[5]
rlabel metal2 40040 15008 40040 15008 0 sel[6]
rlabel metal2 16184 2478 16184 2478 0 sel[7]
rlabel metal3 1358 18200 1358 18200 0 sel[8]
rlabel metal3 1358 22904 1358 22904 0 sel[9]
<< properties >>
string FIXED_BBOX 0 0 42000 42000
<< end >>
