magic
tech gf180mcuD
magscale 1 10
timestamp 1699645710
<< metal1 >>
rect 1344 38442 40656 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 40656 38442
rect 1344 38356 40656 38390
rect 22094 38274 22146 38286
rect 22094 38210 22146 38222
rect 26126 38274 26178 38286
rect 26126 38210 26178 38222
rect 21074 37998 21086 38050
rect 21138 37998 21150 38050
rect 25330 37998 25342 38050
rect 25394 37998 25406 38050
rect 29150 37938 29202 37950
rect 29150 37874 29202 37886
rect 1344 37658 40656 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 40656 37658
rect 1344 37572 40656 37606
rect 20750 37490 20802 37502
rect 20750 37426 20802 37438
rect 19730 37214 19742 37266
rect 19794 37214 19806 37266
rect 1344 36874 40656 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 40656 36874
rect 1344 36788 40656 36822
rect 1344 36090 40656 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 40656 36090
rect 1344 36004 40656 36038
rect 1344 35306 40656 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 40656 35306
rect 1344 35220 40656 35254
rect 1344 34522 40656 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 40656 34522
rect 1344 34436 40656 34470
rect 1344 33738 40656 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 40656 33738
rect 1344 33652 40656 33686
rect 1344 32954 40656 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 40656 32954
rect 1344 32868 40656 32902
rect 1344 32170 40656 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 40656 32170
rect 1344 32084 40656 32118
rect 1344 31386 40656 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 40656 31386
rect 1344 31300 40656 31334
rect 1344 30602 40656 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 40656 30602
rect 1344 30516 40656 30550
rect 1344 29818 40656 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 40656 29818
rect 1344 29732 40656 29766
rect 1344 29034 40656 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 40656 29034
rect 1344 28948 40656 28982
rect 20078 28642 20130 28654
rect 20078 28578 20130 28590
rect 1344 28250 40656 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 40656 28250
rect 1344 28164 40656 28198
rect 21870 27858 21922 27870
rect 21298 27806 21310 27858
rect 21362 27806 21374 27858
rect 21870 27794 21922 27806
rect 25678 27746 25730 27758
rect 18386 27694 18398 27746
rect 18450 27694 18462 27746
rect 20514 27694 20526 27746
rect 20578 27694 20590 27746
rect 25678 27682 25730 27694
rect 1344 27466 40656 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 40656 27466
rect 1344 27380 40656 27414
rect 1934 27186 1986 27198
rect 20638 27186 20690 27198
rect 40014 27186 40066 27198
rect 19842 27134 19854 27186
rect 19906 27134 19918 27186
rect 25330 27134 25342 27186
rect 25394 27134 25406 27186
rect 28578 27134 28590 27186
rect 28642 27134 28654 27186
rect 1934 27122 1986 27134
rect 20638 27122 20690 27134
rect 40014 27122 40066 27134
rect 20862 27074 20914 27086
rect 4274 27022 4286 27074
rect 4338 27022 4350 27074
rect 17042 27022 17054 27074
rect 17106 27022 17118 27074
rect 17714 27022 17726 27074
rect 17778 27022 17790 27074
rect 20862 27010 20914 27022
rect 21646 27074 21698 27086
rect 21646 27010 21698 27022
rect 21758 27074 21810 27086
rect 21758 27010 21810 27022
rect 21982 27074 22034 27086
rect 22418 27022 22430 27074
rect 22482 27022 22494 27074
rect 25666 27022 25678 27074
rect 25730 27022 25742 27074
rect 37650 27022 37662 27074
rect 37714 27022 37726 27074
rect 21982 27010 22034 27022
rect 14702 26962 14754 26974
rect 14702 26898 14754 26910
rect 15150 26962 15202 26974
rect 15150 26898 15202 26910
rect 20190 26962 20242 26974
rect 20190 26898 20242 26910
rect 20414 26962 20466 26974
rect 20414 26898 20466 26910
rect 21310 26962 21362 26974
rect 23202 26910 23214 26962
rect 23266 26910 23278 26962
rect 26450 26910 26462 26962
rect 26514 26910 26526 26962
rect 21310 26898 21362 26910
rect 14590 26850 14642 26862
rect 14590 26786 14642 26798
rect 14814 26850 14866 26862
rect 14814 26786 14866 26798
rect 14926 26850 14978 26862
rect 14926 26786 14978 26798
rect 15822 26850 15874 26862
rect 15822 26786 15874 26798
rect 1344 26682 40656 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 40656 26682
rect 1344 26596 40656 26630
rect 15934 26514 15986 26526
rect 19854 26514 19906 26526
rect 18834 26462 18846 26514
rect 18898 26462 18910 26514
rect 15934 26450 15986 26462
rect 19854 26450 19906 26462
rect 20862 26514 20914 26526
rect 20862 26450 20914 26462
rect 22990 26514 23042 26526
rect 22990 26450 23042 26462
rect 24446 26514 24498 26526
rect 24446 26450 24498 26462
rect 16158 26402 16210 26414
rect 14802 26350 14814 26402
rect 14866 26350 14878 26402
rect 16158 26338 16210 26350
rect 20750 26402 20802 26414
rect 24558 26402 24610 26414
rect 23986 26350 23998 26402
rect 24050 26350 24062 26402
rect 20750 26338 20802 26350
rect 24558 26338 24610 26350
rect 26686 26402 26738 26414
rect 27794 26350 27806 26402
rect 27858 26350 27870 26402
rect 26686 26338 26738 26350
rect 16270 26290 16322 26302
rect 15474 26238 15486 26290
rect 15538 26238 15550 26290
rect 16270 26226 16322 26238
rect 16718 26290 16770 26302
rect 19630 26290 19682 26302
rect 19058 26238 19070 26290
rect 19122 26238 19134 26290
rect 16718 26226 16770 26238
rect 19630 26226 19682 26238
rect 19742 26290 19794 26302
rect 19742 26226 19794 26238
rect 19966 26290 20018 26302
rect 20638 26290 20690 26302
rect 20178 26238 20190 26290
rect 20242 26238 20254 26290
rect 19966 26226 20018 26238
rect 20638 26226 20690 26238
rect 20974 26290 21026 26302
rect 22878 26290 22930 26302
rect 21186 26238 21198 26290
rect 21250 26238 21262 26290
rect 22642 26238 22654 26290
rect 22706 26238 22718 26290
rect 20974 26226 21026 26238
rect 22878 26226 22930 26238
rect 23102 26290 23154 26302
rect 23102 26226 23154 26238
rect 23214 26290 23266 26302
rect 23214 26226 23266 26238
rect 23662 26290 23714 26302
rect 23662 26226 23714 26238
rect 24222 26290 24274 26302
rect 27570 26238 27582 26290
rect 27634 26238 27646 26290
rect 37650 26238 37662 26290
rect 37714 26238 37726 26290
rect 24222 26226 24274 26238
rect 25342 26178 25394 26190
rect 12674 26126 12686 26178
rect 12738 26126 12750 26178
rect 39890 26126 39902 26178
rect 39954 26126 39966 26178
rect 25342 26114 25394 26126
rect 26574 26066 26626 26078
rect 26574 26002 26626 26014
rect 1344 25898 40656 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 40656 25898
rect 1344 25812 40656 25846
rect 16942 25618 16994 25630
rect 16482 25566 16494 25618
rect 16546 25566 16558 25618
rect 16942 25554 16994 25566
rect 20190 25618 20242 25630
rect 20190 25554 20242 25566
rect 23102 25618 23154 25630
rect 23102 25554 23154 25566
rect 25118 25618 25170 25630
rect 25118 25554 25170 25566
rect 17278 25506 17330 25518
rect 13682 25454 13694 25506
rect 13746 25454 13758 25506
rect 17278 25442 17330 25454
rect 17838 25506 17890 25518
rect 17838 25442 17890 25454
rect 19294 25506 19346 25518
rect 25006 25506 25058 25518
rect 19954 25454 19966 25506
rect 20018 25454 20030 25506
rect 24770 25454 24782 25506
rect 24834 25454 24846 25506
rect 19294 25442 19346 25454
rect 25006 25442 25058 25454
rect 20302 25394 20354 25406
rect 14354 25342 14366 25394
rect 14418 25342 14430 25394
rect 19618 25342 19630 25394
rect 19682 25342 19694 25394
rect 20302 25330 20354 25342
rect 25454 25394 25506 25406
rect 25454 25330 25506 25342
rect 22318 25282 22370 25294
rect 21970 25230 21982 25282
rect 22034 25230 22046 25282
rect 22318 25218 22370 25230
rect 22766 25282 22818 25294
rect 22766 25218 22818 25230
rect 22990 25282 23042 25294
rect 22990 25218 23042 25230
rect 23214 25282 23266 25294
rect 23214 25218 23266 25230
rect 25230 25282 25282 25294
rect 25230 25218 25282 25230
rect 1344 25114 40656 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 40656 25114
rect 1344 25028 40656 25062
rect 15374 24946 15426 24958
rect 15374 24882 15426 24894
rect 17502 24946 17554 24958
rect 17502 24882 17554 24894
rect 19182 24946 19234 24958
rect 19182 24882 19234 24894
rect 22542 24946 22594 24958
rect 22542 24882 22594 24894
rect 22766 24946 22818 24958
rect 22766 24882 22818 24894
rect 15486 24834 15538 24846
rect 17390 24834 17442 24846
rect 16370 24782 16382 24834
rect 16434 24782 16446 24834
rect 15486 24770 15538 24782
rect 17390 24770 17442 24782
rect 20974 24834 21026 24846
rect 20974 24770 21026 24782
rect 22430 24834 22482 24846
rect 22430 24770 22482 24782
rect 17614 24722 17666 24734
rect 16594 24670 16606 24722
rect 16658 24670 16670 24722
rect 17614 24658 17666 24670
rect 17950 24722 18002 24734
rect 20862 24722 20914 24734
rect 20402 24670 20414 24722
rect 20466 24670 20478 24722
rect 17950 24658 18002 24670
rect 20862 24658 20914 24670
rect 19070 24610 19122 24622
rect 19070 24546 19122 24558
rect 25566 24610 25618 24622
rect 25566 24546 25618 24558
rect 15262 24498 15314 24510
rect 15262 24434 15314 24446
rect 20638 24498 20690 24510
rect 20638 24434 20690 24446
rect 1344 24330 40656 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 40656 24330
rect 1344 24244 40656 24278
rect 13918 24162 13970 24174
rect 13918 24098 13970 24110
rect 23774 24162 23826 24174
rect 23774 24098 23826 24110
rect 18958 24050 19010 24062
rect 18050 23998 18062 24050
rect 18114 23998 18126 24050
rect 18958 23986 19010 23998
rect 19630 24050 19682 24062
rect 19630 23986 19682 23998
rect 23438 24050 23490 24062
rect 40014 24050 40066 24062
rect 28578 23998 28590 24050
rect 28642 23998 28654 24050
rect 23438 23986 23490 23998
rect 40014 23986 40066 23998
rect 24894 23938 24946 23950
rect 13906 23886 13918 23938
rect 13970 23886 13982 23938
rect 18722 23886 18734 23938
rect 18786 23886 18798 23938
rect 19842 23886 19854 23938
rect 19906 23886 19918 23938
rect 24894 23874 24946 23886
rect 25118 23938 25170 23950
rect 25666 23886 25678 23938
rect 25730 23886 25742 23938
rect 37650 23886 37662 23938
rect 37714 23886 37726 23938
rect 25118 23874 25170 23886
rect 13582 23826 13634 23838
rect 13582 23762 13634 23774
rect 18398 23826 18450 23838
rect 18398 23762 18450 23774
rect 19070 23826 19122 23838
rect 19070 23762 19122 23774
rect 19518 23826 19570 23838
rect 25230 23826 25282 23838
rect 20626 23774 20638 23826
rect 20690 23774 20702 23826
rect 19518 23762 19570 23774
rect 25230 23762 25282 23774
rect 25342 23826 25394 23838
rect 26450 23774 26462 23826
rect 26514 23774 26526 23826
rect 25342 23762 25394 23774
rect 18174 23714 18226 23726
rect 18174 23650 18226 23662
rect 20302 23714 20354 23726
rect 20302 23650 20354 23662
rect 23662 23714 23714 23726
rect 23662 23650 23714 23662
rect 1344 23546 40656 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 40656 23546
rect 1344 23460 40656 23494
rect 16606 23378 16658 23390
rect 16606 23314 16658 23326
rect 19406 23266 19458 23278
rect 21310 23266 21362 23278
rect 20402 23214 20414 23266
rect 20466 23214 20478 23266
rect 19406 23202 19458 23214
rect 21310 23202 21362 23214
rect 21534 23266 21586 23278
rect 21534 23202 21586 23214
rect 16270 23154 16322 23166
rect 10882 23102 10894 23154
rect 10946 23102 10958 23154
rect 14802 23102 14814 23154
rect 14866 23102 14878 23154
rect 16270 23090 16322 23102
rect 17726 23154 17778 23166
rect 17726 23090 17778 23102
rect 18398 23154 18450 23166
rect 18398 23090 18450 23102
rect 18622 23154 18674 23166
rect 18622 23090 18674 23102
rect 19070 23154 19122 23166
rect 19070 23090 19122 23102
rect 19742 23154 19794 23166
rect 23214 23154 23266 23166
rect 20178 23102 20190 23154
rect 20242 23102 20254 23154
rect 22978 23102 22990 23154
rect 23042 23102 23054 23154
rect 19742 23090 19794 23102
rect 23214 23090 23266 23102
rect 23998 23154 24050 23166
rect 23998 23090 24050 23102
rect 24446 23154 24498 23166
rect 24446 23090 24498 23102
rect 24558 23154 24610 23166
rect 25890 23102 25902 23154
rect 25954 23102 25966 23154
rect 37650 23102 37662 23154
rect 37714 23102 37726 23154
rect 24558 23090 24610 23102
rect 14142 23042 14194 23054
rect 17502 23042 17554 23054
rect 11666 22990 11678 23042
rect 11730 22990 11742 23042
rect 13794 22990 13806 23042
rect 13858 22990 13870 23042
rect 14466 22990 14478 23042
rect 14530 22990 14542 23042
rect 14142 22978 14194 22990
rect 17502 22978 17554 22990
rect 18846 23042 18898 23054
rect 18846 22978 18898 22990
rect 24222 23042 24274 23054
rect 24222 22978 24274 22990
rect 25342 23042 25394 23054
rect 26674 22990 26686 23042
rect 26738 22990 26750 23042
rect 28802 22990 28814 23042
rect 28866 22990 28878 23042
rect 25342 22978 25394 22990
rect 21646 22930 21698 22942
rect 18050 22878 18062 22930
rect 18114 22878 18126 22930
rect 21646 22866 21698 22878
rect 23326 22930 23378 22942
rect 40014 22930 40066 22942
rect 25442 22878 25454 22930
rect 25506 22927 25518 22930
rect 25666 22927 25678 22930
rect 25506 22881 25678 22927
rect 25506 22878 25518 22881
rect 25666 22878 25678 22881
rect 25730 22878 25742 22930
rect 23326 22866 23378 22878
rect 40014 22866 40066 22878
rect 1344 22762 40656 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 40656 22762
rect 1344 22676 40656 22710
rect 21534 22594 21586 22606
rect 21534 22530 21586 22542
rect 19742 22482 19794 22494
rect 10770 22430 10782 22482
rect 10834 22430 10846 22482
rect 12898 22430 12910 22482
rect 12962 22430 12974 22482
rect 19742 22418 19794 22430
rect 20302 22482 20354 22494
rect 20302 22418 20354 22430
rect 25790 22482 25842 22494
rect 25790 22418 25842 22430
rect 26350 22482 26402 22494
rect 26350 22418 26402 22430
rect 13918 22370 13970 22382
rect 10098 22318 10110 22370
rect 10162 22318 10174 22370
rect 13918 22306 13970 22318
rect 14366 22370 14418 22382
rect 17390 22370 17442 22382
rect 22878 22370 22930 22382
rect 16258 22318 16270 22370
rect 16322 22318 16334 22370
rect 16930 22318 16942 22370
rect 16994 22318 17006 22370
rect 19506 22318 19518 22370
rect 19570 22318 19582 22370
rect 14366 22306 14418 22318
rect 17390 22306 17442 22318
rect 22878 22306 22930 22318
rect 23102 22370 23154 22382
rect 23662 22370 23714 22382
rect 23426 22318 23438 22370
rect 23490 22318 23502 22370
rect 23102 22306 23154 22318
rect 23662 22306 23714 22318
rect 23886 22370 23938 22382
rect 24334 22370 24386 22382
rect 24098 22318 24110 22370
rect 24162 22318 24174 22370
rect 23886 22306 23938 22318
rect 24334 22306 24386 22318
rect 24782 22370 24834 22382
rect 24782 22306 24834 22318
rect 24894 22370 24946 22382
rect 24894 22306 24946 22318
rect 25566 22370 25618 22382
rect 25566 22306 25618 22318
rect 26574 22370 26626 22382
rect 26574 22306 26626 22318
rect 26686 22370 26738 22382
rect 26686 22306 26738 22318
rect 13582 22258 13634 22270
rect 18510 22258 18562 22270
rect 15922 22206 15934 22258
rect 15986 22206 15998 22258
rect 13582 22194 13634 22206
rect 18510 22194 18562 22206
rect 21310 22258 21362 22270
rect 21310 22194 21362 22206
rect 22542 22258 22594 22270
rect 22542 22194 22594 22206
rect 25342 22258 25394 22270
rect 25342 22194 25394 22206
rect 25902 22258 25954 22270
rect 25902 22194 25954 22206
rect 26238 22258 26290 22270
rect 26238 22194 26290 22206
rect 17502 22146 17554 22158
rect 22766 22146 22818 22158
rect 16818 22094 16830 22146
rect 16882 22094 16894 22146
rect 21858 22094 21870 22146
rect 21922 22094 21934 22146
rect 17502 22082 17554 22094
rect 22766 22082 22818 22094
rect 23774 22146 23826 22158
rect 23774 22082 23826 22094
rect 24670 22146 24722 22158
rect 24670 22082 24722 22094
rect 1344 21978 40656 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 40656 21978
rect 1344 21892 40656 21926
rect 13134 21810 13186 21822
rect 16494 21810 16546 21822
rect 15138 21758 15150 21810
rect 15202 21758 15214 21810
rect 16146 21758 16158 21810
rect 16210 21758 16222 21810
rect 13134 21746 13186 21758
rect 16494 21746 16546 21758
rect 26014 21810 26066 21822
rect 26014 21746 26066 21758
rect 14814 21698 14866 21710
rect 25230 21698 25282 21710
rect 14130 21646 14142 21698
rect 14194 21646 14206 21698
rect 15810 21646 15822 21698
rect 15874 21646 15886 21698
rect 14814 21634 14866 21646
rect 25230 21634 25282 21646
rect 25566 21698 25618 21710
rect 25566 21634 25618 21646
rect 26238 21698 26290 21710
rect 26238 21634 26290 21646
rect 17838 21586 17890 21598
rect 24558 21586 24610 21598
rect 14354 21534 14366 21586
rect 14418 21534 14430 21586
rect 15586 21534 15598 21586
rect 15650 21534 15662 21586
rect 18162 21534 18174 21586
rect 18226 21534 18238 21586
rect 23762 21534 23774 21586
rect 23826 21534 23838 21586
rect 24322 21534 24334 21586
rect 24386 21534 24398 21586
rect 17838 21522 17890 21534
rect 24558 21522 24610 21534
rect 25790 21586 25842 21598
rect 25790 21522 25842 21534
rect 26350 21586 26402 21598
rect 37650 21534 37662 21586
rect 37714 21534 37726 21586
rect 26350 21522 26402 21534
rect 24446 21474 24498 21486
rect 21634 21422 21646 21474
rect 21698 21422 21710 21474
rect 24446 21410 24498 21422
rect 25342 21474 25394 21486
rect 25342 21410 25394 21422
rect 40014 21362 40066 21374
rect 23986 21310 23998 21362
rect 24050 21310 24062 21362
rect 40014 21298 40066 21310
rect 1344 21194 40656 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 40656 21194
rect 1344 21108 40656 21142
rect 19182 21026 19234 21038
rect 19182 20962 19234 20974
rect 1934 20914 1986 20926
rect 1934 20850 1986 20862
rect 18622 20914 18674 20926
rect 18622 20850 18674 20862
rect 14702 20802 14754 20814
rect 4162 20750 4174 20802
rect 4226 20750 4238 20802
rect 14702 20738 14754 20750
rect 16942 20802 16994 20814
rect 16942 20738 16994 20750
rect 17502 20802 17554 20814
rect 18846 20802 18898 20814
rect 20526 20802 20578 20814
rect 18050 20750 18062 20802
rect 18114 20750 18126 20802
rect 19618 20750 19630 20802
rect 19682 20750 19694 20802
rect 20178 20750 20190 20802
rect 20242 20750 20254 20802
rect 17502 20738 17554 20750
rect 18846 20738 18898 20750
rect 20526 20738 20578 20750
rect 20862 20802 20914 20814
rect 21634 20750 21646 20802
rect 21698 20750 21710 20802
rect 20862 20738 20914 20750
rect 25666 20638 25678 20690
rect 25730 20638 25742 20690
rect 15026 20526 15038 20578
rect 15090 20526 15102 20578
rect 18274 20526 18286 20578
rect 18338 20526 18350 20578
rect 1344 20410 40656 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 40656 20410
rect 1344 20324 40656 20358
rect 13134 20242 13186 20254
rect 13134 20178 13186 20190
rect 15374 20242 15426 20254
rect 15374 20178 15426 20190
rect 15598 20242 15650 20254
rect 15598 20178 15650 20190
rect 14366 20130 14418 20142
rect 14366 20066 14418 20078
rect 14478 20130 14530 20142
rect 14478 20066 14530 20078
rect 15486 20130 15538 20142
rect 15486 20066 15538 20078
rect 16270 20130 16322 20142
rect 16270 20066 16322 20078
rect 18846 20130 18898 20142
rect 18846 20066 18898 20078
rect 21310 20130 21362 20142
rect 21310 20066 21362 20078
rect 22430 20130 22482 20142
rect 22430 20066 22482 20078
rect 22654 20130 22706 20142
rect 22654 20066 22706 20078
rect 22990 20130 23042 20142
rect 22990 20066 23042 20078
rect 23774 20130 23826 20142
rect 23986 20078 23998 20130
rect 24050 20078 24062 20130
rect 26450 20078 26462 20130
rect 26514 20078 26526 20130
rect 23774 20066 23826 20078
rect 14702 20018 14754 20030
rect 4274 19966 4286 20018
rect 4338 19966 4350 20018
rect 13906 19966 13918 20018
rect 13970 19966 13982 20018
rect 14702 19954 14754 19966
rect 14926 20018 14978 20030
rect 14926 19954 14978 19966
rect 16382 20018 16434 20030
rect 16382 19954 16434 19966
rect 16606 20018 16658 20030
rect 19630 20018 19682 20030
rect 22318 20018 22370 20030
rect 16818 19966 16830 20018
rect 16882 19966 16894 20018
rect 19394 19966 19406 20018
rect 19458 19966 19470 20018
rect 20514 19966 20526 20018
rect 20578 19966 20590 20018
rect 16606 19954 16658 19966
rect 19630 19954 19682 19966
rect 22318 19954 22370 19966
rect 22878 20018 22930 20030
rect 22878 19954 22930 19966
rect 24222 20018 24274 20030
rect 24222 19954 24274 19966
rect 24670 20018 24722 20030
rect 25666 19966 25678 20018
rect 25730 19966 25742 20018
rect 37650 19966 37662 20018
rect 37714 19966 37726 20018
rect 24670 19954 24722 19966
rect 11790 19906 11842 19918
rect 20974 19906 21026 19918
rect 24446 19906 24498 19918
rect 14354 19854 14366 19906
rect 14418 19854 14430 19906
rect 16258 19854 16270 19906
rect 16322 19854 16334 19906
rect 20178 19854 20190 19906
rect 20242 19854 20254 19906
rect 21746 19854 21758 19906
rect 21810 19854 21822 19906
rect 11790 19842 11842 19854
rect 20974 19842 21026 19854
rect 24446 19842 24498 19854
rect 24558 19906 24610 19918
rect 24558 19842 24610 19854
rect 25342 19906 25394 19918
rect 28578 19854 28590 19906
rect 28642 19854 28654 19906
rect 25342 19842 25394 19854
rect 1934 19794 1986 19806
rect 1934 19730 1986 19742
rect 11902 19794 11954 19806
rect 11902 19730 11954 19742
rect 22990 19794 23042 19806
rect 22990 19730 23042 19742
rect 40014 19794 40066 19806
rect 40014 19730 40066 19742
rect 1344 19626 40656 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 40656 19626
rect 1344 19540 40656 19574
rect 15150 19458 15202 19470
rect 15150 19394 15202 19406
rect 1934 19346 1986 19358
rect 9874 19294 9886 19346
rect 9938 19294 9950 19346
rect 12114 19294 12126 19346
rect 12178 19294 12190 19346
rect 14802 19294 14814 19346
rect 14866 19294 14878 19346
rect 17042 19294 17054 19346
rect 17106 19294 17118 19346
rect 26450 19294 26462 19346
rect 26514 19294 26526 19346
rect 28578 19294 28590 19346
rect 28642 19294 28654 19346
rect 1934 19282 1986 19294
rect 22206 19234 22258 19246
rect 24446 19234 24498 19246
rect 4274 19182 4286 19234
rect 4338 19182 4350 19234
rect 12898 19182 12910 19234
rect 12962 19182 12974 19234
rect 13682 19182 13694 19234
rect 13746 19182 13758 19234
rect 19842 19182 19854 19234
rect 19906 19182 19918 19234
rect 23986 19182 23998 19234
rect 24050 19182 24062 19234
rect 22206 19170 22258 19182
rect 24446 19170 24498 19182
rect 24558 19234 24610 19246
rect 25666 19182 25678 19234
rect 25730 19182 25742 19234
rect 24558 19170 24610 19182
rect 13458 19070 13470 19122
rect 13522 19070 13534 19122
rect 14926 19010 14978 19022
rect 24222 19010 24274 19022
rect 21858 18958 21870 19010
rect 21922 18958 21934 19010
rect 14926 18946 14978 18958
rect 24222 18946 24274 18958
rect 24334 19010 24386 19022
rect 24334 18946 24386 18958
rect 25342 19010 25394 19022
rect 25342 18946 25394 18958
rect 1344 18842 40656 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 40656 18842
rect 1344 18756 40656 18790
rect 20750 18674 20802 18686
rect 12450 18622 12462 18674
rect 12514 18622 12526 18674
rect 20402 18622 20414 18674
rect 20466 18622 20478 18674
rect 20750 18610 20802 18622
rect 21086 18674 21138 18686
rect 21410 18622 21422 18674
rect 21474 18622 21486 18674
rect 21086 18610 21138 18622
rect 23998 18562 24050 18574
rect 23998 18498 24050 18510
rect 24222 18562 24274 18574
rect 24222 18498 24274 18510
rect 17502 18450 17554 18462
rect 4274 18398 4286 18450
rect 4338 18398 4350 18450
rect 12674 18398 12686 18450
rect 12738 18398 12750 18450
rect 16594 18398 16606 18450
rect 16658 18398 16670 18450
rect 17502 18386 17554 18398
rect 19630 18450 19682 18462
rect 19630 18386 19682 18398
rect 23662 18450 23714 18462
rect 23662 18386 23714 18398
rect 27918 18450 27970 18462
rect 27918 18386 27970 18398
rect 28030 18450 28082 18462
rect 37650 18398 37662 18450
rect 37714 18398 37726 18450
rect 28030 18386 28082 18398
rect 23774 18338 23826 18350
rect 13682 18286 13694 18338
rect 13746 18286 13758 18338
rect 15810 18286 15822 18338
rect 15874 18286 15886 18338
rect 19170 18286 19182 18338
rect 19234 18286 19246 18338
rect 23774 18274 23826 18286
rect 1934 18226 1986 18238
rect 1934 18162 1986 18174
rect 40014 18226 40066 18238
rect 40014 18162 40066 18174
rect 1344 18058 40656 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 40656 18058
rect 1344 17972 40656 18006
rect 15374 17890 15426 17902
rect 15374 17826 15426 17838
rect 20638 17890 20690 17902
rect 20638 17826 20690 17838
rect 1934 17778 1986 17790
rect 1934 17714 1986 17726
rect 15262 17778 15314 17790
rect 21298 17726 21310 17778
rect 21362 17726 21374 17778
rect 23986 17726 23998 17778
rect 24050 17726 24062 17778
rect 26114 17726 26126 17778
rect 26178 17726 26190 17778
rect 15262 17714 15314 17726
rect 15710 17666 15762 17678
rect 4274 17614 4286 17666
rect 4338 17614 4350 17666
rect 15026 17614 15038 17666
rect 15090 17614 15102 17666
rect 15710 17602 15762 17614
rect 15934 17666 15986 17678
rect 15934 17602 15986 17614
rect 16382 17666 16434 17678
rect 18958 17666 19010 17678
rect 17602 17614 17614 17666
rect 17666 17614 17678 17666
rect 16382 17602 16434 17614
rect 18958 17602 19010 17614
rect 19294 17666 19346 17678
rect 19294 17602 19346 17614
rect 19630 17666 19682 17678
rect 20750 17666 20802 17678
rect 20066 17614 20078 17666
rect 20130 17614 20142 17666
rect 22194 17614 22206 17666
rect 22258 17614 22270 17666
rect 23202 17614 23214 17666
rect 23266 17614 23278 17666
rect 19630 17602 19682 17614
rect 20750 17602 20802 17614
rect 14254 17554 14306 17566
rect 14254 17490 14306 17502
rect 14478 17554 14530 17566
rect 14478 17490 14530 17502
rect 20302 17554 20354 17566
rect 20302 17490 20354 17502
rect 21422 17554 21474 17566
rect 21422 17490 21474 17502
rect 21646 17554 21698 17566
rect 21646 17490 21698 17502
rect 14366 17442 14418 17454
rect 14366 17378 14418 17390
rect 15822 17442 15874 17454
rect 19182 17442 19234 17454
rect 26574 17442 26626 17454
rect 17378 17390 17390 17442
rect 17442 17390 17454 17442
rect 21970 17390 21982 17442
rect 22034 17390 22046 17442
rect 15822 17378 15874 17390
rect 19182 17378 19234 17390
rect 26574 17378 26626 17390
rect 1344 17274 40656 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 40656 17274
rect 1344 17188 40656 17222
rect 14478 17106 14530 17118
rect 14478 17042 14530 17054
rect 14590 17106 14642 17118
rect 14590 17042 14642 17054
rect 15374 17106 15426 17118
rect 15374 17042 15426 17054
rect 17614 17106 17666 17118
rect 17614 17042 17666 17054
rect 24446 16994 24498 17006
rect 13234 16942 13246 16994
rect 13298 16942 13310 16994
rect 18722 16942 18734 16994
rect 18786 16942 18798 16994
rect 22866 16942 22878 16994
rect 22930 16991 22942 16994
rect 23202 16991 23214 16994
rect 22930 16945 23214 16991
rect 22930 16942 22942 16945
rect 23202 16942 23214 16945
rect 23266 16942 23278 16994
rect 24446 16930 24498 16942
rect 14366 16882 14418 16894
rect 14018 16830 14030 16882
rect 14082 16830 14094 16882
rect 14914 16830 14926 16882
rect 14978 16830 14990 16882
rect 17938 16830 17950 16882
rect 18002 16830 18014 16882
rect 23314 16830 23326 16882
rect 23378 16830 23390 16882
rect 14366 16818 14418 16830
rect 23550 16770 23602 16782
rect 11106 16718 11118 16770
rect 11170 16718 11182 16770
rect 20850 16718 20862 16770
rect 20914 16718 20926 16770
rect 23550 16706 23602 16718
rect 24222 16770 24274 16782
rect 24222 16706 24274 16718
rect 24334 16770 24386 16782
rect 24334 16706 24386 16718
rect 23774 16658 23826 16670
rect 23774 16594 23826 16606
rect 23886 16658 23938 16670
rect 23886 16594 23938 16606
rect 1344 16490 40656 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 40656 16490
rect 1344 16404 40656 16438
rect 18510 16322 18562 16334
rect 18510 16258 18562 16270
rect 14254 16210 14306 16222
rect 26238 16210 26290 16222
rect 19394 16158 19406 16210
rect 19458 16158 19470 16210
rect 23650 16158 23662 16210
rect 23714 16158 23726 16210
rect 25778 16158 25790 16210
rect 25842 16158 25854 16210
rect 14254 16146 14306 16158
rect 26238 16146 26290 16158
rect 22866 16046 22878 16098
rect 22930 16046 22942 16098
rect 18398 15986 18450 15998
rect 18398 15922 18450 15934
rect 19518 15986 19570 15998
rect 19518 15922 19570 15934
rect 19742 15986 19794 15998
rect 19742 15922 19794 15934
rect 16382 15874 16434 15886
rect 16034 15822 16046 15874
rect 16098 15822 16110 15874
rect 16382 15810 16434 15822
rect 18510 15874 18562 15886
rect 18510 15810 18562 15822
rect 1344 15706 40656 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 40656 15706
rect 1344 15620 40656 15654
rect 16606 15538 16658 15550
rect 16606 15474 16658 15486
rect 17502 15538 17554 15550
rect 17502 15474 17554 15486
rect 20190 15538 20242 15550
rect 20190 15474 20242 15486
rect 20302 15538 20354 15550
rect 20302 15474 20354 15486
rect 20638 15538 20690 15550
rect 20638 15474 20690 15486
rect 21198 15538 21250 15550
rect 21198 15474 21250 15486
rect 15374 15426 15426 15438
rect 15374 15362 15426 15374
rect 22990 15426 23042 15438
rect 22990 15362 23042 15374
rect 15150 15314 15202 15326
rect 19070 15314 19122 15326
rect 15586 15262 15598 15314
rect 15650 15262 15662 15314
rect 15810 15262 15822 15314
rect 15874 15262 15886 15314
rect 15150 15250 15202 15262
rect 19070 15250 19122 15262
rect 19406 15314 19458 15326
rect 20414 15314 20466 15326
rect 19842 15262 19854 15314
rect 19906 15262 19918 15314
rect 19406 15250 19458 15262
rect 20414 15250 20466 15262
rect 22542 15314 22594 15326
rect 22542 15250 22594 15262
rect 23102 15314 23154 15326
rect 23102 15250 23154 15262
rect 14366 15202 14418 15214
rect 14366 15138 14418 15150
rect 15262 15202 15314 15214
rect 15262 15138 15314 15150
rect 19182 15202 19234 15214
rect 19182 15138 19234 15150
rect 22766 15202 22818 15214
rect 22766 15138 22818 15150
rect 14254 15090 14306 15102
rect 14254 15026 14306 15038
rect 19518 15090 19570 15102
rect 19518 15026 19570 15038
rect 1344 14922 40656 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 40656 14922
rect 1344 14836 40656 14870
rect 17054 14754 17106 14766
rect 17054 14690 17106 14702
rect 22542 14754 22594 14766
rect 22542 14690 22594 14702
rect 22094 14642 22146 14654
rect 14242 14590 14254 14642
rect 14306 14590 14318 14642
rect 16370 14590 16382 14642
rect 16434 14590 16446 14642
rect 18610 14590 18622 14642
rect 18674 14590 18686 14642
rect 20738 14590 20750 14642
rect 20802 14590 20814 14642
rect 22094 14578 22146 14590
rect 17502 14530 17554 14542
rect 22430 14530 22482 14542
rect 13570 14478 13582 14530
rect 13634 14478 13646 14530
rect 16818 14478 16830 14530
rect 16882 14478 16894 14530
rect 17826 14478 17838 14530
rect 17890 14478 17902 14530
rect 23986 14478 23998 14530
rect 24050 14478 24062 14530
rect 17502 14466 17554 14478
rect 22430 14466 22482 14478
rect 17266 14366 17278 14418
rect 17330 14366 17342 14418
rect 22542 14306 22594 14318
rect 17042 14254 17054 14306
rect 17106 14254 17118 14306
rect 24210 14254 24222 14306
rect 24274 14254 24286 14306
rect 22542 14242 22594 14254
rect 1344 14138 40656 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 40656 14138
rect 1344 14052 40656 14086
rect 17390 13970 17442 13982
rect 17390 13906 17442 13918
rect 25342 13970 25394 13982
rect 25342 13906 25394 13918
rect 14690 13806 14702 13858
rect 14754 13806 14766 13858
rect 18834 13806 18846 13858
rect 18898 13806 18910 13858
rect 22530 13806 22542 13858
rect 22594 13806 22606 13858
rect 13906 13694 13918 13746
rect 13970 13694 13982 13746
rect 18050 13694 18062 13746
rect 18114 13694 18126 13746
rect 21858 13694 21870 13746
rect 21922 13694 21934 13746
rect 17502 13634 17554 13646
rect 16818 13582 16830 13634
rect 16882 13582 16894 13634
rect 20962 13582 20974 13634
rect 21026 13582 21038 13634
rect 24658 13582 24670 13634
rect 24722 13582 24734 13634
rect 17502 13570 17554 13582
rect 1344 13354 40656 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 40656 13354
rect 1344 13268 40656 13302
rect 20190 13186 20242 13198
rect 20190 13122 20242 13134
rect 17166 13074 17218 13086
rect 17166 13010 17218 13022
rect 17838 13074 17890 13086
rect 17838 13010 17890 13022
rect 20302 12962 20354 12974
rect 20302 12898 20354 12910
rect 24222 12738 24274 12750
rect 23874 12686 23886 12738
rect 23938 12686 23950 12738
rect 24222 12674 24274 12686
rect 1344 12570 40656 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 40656 12570
rect 1344 12484 40656 12518
rect 40238 12290 40290 12302
rect 40238 12226 40290 12238
rect 1344 11786 40656 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 40656 11786
rect 1344 11700 40656 11734
rect 1344 11002 40656 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 40656 11002
rect 1344 10916 40656 10950
rect 1344 10218 40656 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 40656 10218
rect 1344 10132 40656 10166
rect 1344 9434 40656 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 40656 9434
rect 1344 9348 40656 9382
rect 1344 8650 40656 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 40656 8650
rect 1344 8564 40656 8598
rect 1344 7866 40656 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 40656 7866
rect 1344 7780 40656 7814
rect 1344 7082 40656 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 40656 7082
rect 1344 6996 40656 7030
rect 1344 6298 40656 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 40656 6298
rect 1344 6212 40656 6246
rect 1344 5514 40656 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 40656 5514
rect 1344 5428 40656 5462
rect 16718 5234 16770 5246
rect 16718 5170 16770 5182
rect 24782 5234 24834 5246
rect 24782 5170 24834 5182
rect 15698 5070 15710 5122
rect 15762 5070 15774 5122
rect 23762 5070 23774 5122
rect 23826 5070 23838 5122
rect 1344 4730 40656 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 40656 4730
rect 1344 4644 40656 4678
rect 20402 4286 20414 4338
rect 20466 4286 20478 4338
rect 25442 4286 25454 4338
rect 25506 4286 25518 4338
rect 21422 4114 21474 4126
rect 21422 4050 21474 4062
rect 26238 4114 26290 4126
rect 26238 4050 26290 4062
rect 1344 3946 40656 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 40656 3946
rect 1344 3860 40656 3894
rect 22094 3666 22146 3678
rect 22094 3602 22146 3614
rect 25566 3666 25618 3678
rect 25566 3602 25618 3614
rect 29374 3666 29426 3678
rect 29374 3602 29426 3614
rect 17042 3502 17054 3554
rect 17106 3502 17118 3554
rect 21074 3502 21086 3554
rect 21138 3502 21150 3554
rect 24546 3502 24558 3554
rect 24610 3502 24622 3554
rect 28578 3502 28590 3554
rect 28642 3502 28654 3554
rect 18062 3330 18114 3342
rect 18062 3266 18114 3278
rect 1344 3162 40656 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 40656 3162
rect 1344 3076 40656 3110
<< via1 >>
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 22094 38222 22146 38274
rect 26126 38222 26178 38274
rect 21086 37998 21138 38050
rect 25342 37998 25394 38050
rect 29150 37886 29202 37938
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 20750 37438 20802 37490
rect 19742 37214 19794 37266
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 20078 28590 20130 28642
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 21310 27806 21362 27858
rect 21870 27806 21922 27858
rect 18398 27694 18450 27746
rect 20526 27694 20578 27746
rect 25678 27694 25730 27746
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 1934 27134 1986 27186
rect 19854 27134 19906 27186
rect 20638 27134 20690 27186
rect 25342 27134 25394 27186
rect 28590 27134 28642 27186
rect 40014 27134 40066 27186
rect 4286 27022 4338 27074
rect 17054 27022 17106 27074
rect 17726 27022 17778 27074
rect 20862 27022 20914 27074
rect 21646 27022 21698 27074
rect 21758 27022 21810 27074
rect 21982 27022 22034 27074
rect 22430 27022 22482 27074
rect 25678 27022 25730 27074
rect 37662 27022 37714 27074
rect 14702 26910 14754 26962
rect 15150 26910 15202 26962
rect 20190 26910 20242 26962
rect 20414 26910 20466 26962
rect 21310 26910 21362 26962
rect 23214 26910 23266 26962
rect 26462 26910 26514 26962
rect 14590 26798 14642 26850
rect 14814 26798 14866 26850
rect 14926 26798 14978 26850
rect 15822 26798 15874 26850
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 15934 26462 15986 26514
rect 18846 26462 18898 26514
rect 19854 26462 19906 26514
rect 20862 26462 20914 26514
rect 22990 26462 23042 26514
rect 24446 26462 24498 26514
rect 14814 26350 14866 26402
rect 16158 26350 16210 26402
rect 20750 26350 20802 26402
rect 23998 26350 24050 26402
rect 24558 26350 24610 26402
rect 26686 26350 26738 26402
rect 27806 26350 27858 26402
rect 15486 26238 15538 26290
rect 16270 26238 16322 26290
rect 16718 26238 16770 26290
rect 19070 26238 19122 26290
rect 19630 26238 19682 26290
rect 19742 26238 19794 26290
rect 19966 26238 20018 26290
rect 20190 26238 20242 26290
rect 20638 26238 20690 26290
rect 20974 26238 21026 26290
rect 21198 26238 21250 26290
rect 22654 26238 22706 26290
rect 22878 26238 22930 26290
rect 23102 26238 23154 26290
rect 23214 26238 23266 26290
rect 23662 26238 23714 26290
rect 24222 26238 24274 26290
rect 27582 26238 27634 26290
rect 37662 26238 37714 26290
rect 12686 26126 12738 26178
rect 25342 26126 25394 26178
rect 39902 26126 39954 26178
rect 26574 26014 26626 26066
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 16494 25566 16546 25618
rect 16942 25566 16994 25618
rect 20190 25566 20242 25618
rect 23102 25566 23154 25618
rect 25118 25566 25170 25618
rect 13694 25454 13746 25506
rect 17278 25454 17330 25506
rect 17838 25454 17890 25506
rect 19294 25454 19346 25506
rect 19966 25454 20018 25506
rect 24782 25454 24834 25506
rect 25006 25454 25058 25506
rect 14366 25342 14418 25394
rect 19630 25342 19682 25394
rect 20302 25342 20354 25394
rect 25454 25342 25506 25394
rect 21982 25230 22034 25282
rect 22318 25230 22370 25282
rect 22766 25230 22818 25282
rect 22990 25230 23042 25282
rect 23214 25230 23266 25282
rect 25230 25230 25282 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 15374 24894 15426 24946
rect 17502 24894 17554 24946
rect 19182 24894 19234 24946
rect 22542 24894 22594 24946
rect 22766 24894 22818 24946
rect 15486 24782 15538 24834
rect 16382 24782 16434 24834
rect 17390 24782 17442 24834
rect 20974 24782 21026 24834
rect 22430 24782 22482 24834
rect 16606 24670 16658 24722
rect 17614 24670 17666 24722
rect 17950 24670 18002 24722
rect 20414 24670 20466 24722
rect 20862 24670 20914 24722
rect 19070 24558 19122 24610
rect 25566 24558 25618 24610
rect 15262 24446 15314 24498
rect 20638 24446 20690 24498
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 13918 24110 13970 24162
rect 23774 24110 23826 24162
rect 18062 23998 18114 24050
rect 18958 23998 19010 24050
rect 19630 23998 19682 24050
rect 23438 23998 23490 24050
rect 28590 23998 28642 24050
rect 40014 23998 40066 24050
rect 13918 23886 13970 23938
rect 18734 23886 18786 23938
rect 19854 23886 19906 23938
rect 24894 23886 24946 23938
rect 25118 23886 25170 23938
rect 25678 23886 25730 23938
rect 37662 23886 37714 23938
rect 13582 23774 13634 23826
rect 18398 23774 18450 23826
rect 19070 23774 19122 23826
rect 19518 23774 19570 23826
rect 20638 23774 20690 23826
rect 25230 23774 25282 23826
rect 25342 23774 25394 23826
rect 26462 23774 26514 23826
rect 18174 23662 18226 23714
rect 20302 23662 20354 23714
rect 23662 23662 23714 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 16606 23326 16658 23378
rect 19406 23214 19458 23266
rect 20414 23214 20466 23266
rect 21310 23214 21362 23266
rect 21534 23214 21586 23266
rect 10894 23102 10946 23154
rect 14814 23102 14866 23154
rect 16270 23102 16322 23154
rect 17726 23102 17778 23154
rect 18398 23102 18450 23154
rect 18622 23102 18674 23154
rect 19070 23102 19122 23154
rect 19742 23102 19794 23154
rect 20190 23102 20242 23154
rect 22990 23102 23042 23154
rect 23214 23102 23266 23154
rect 23998 23102 24050 23154
rect 24446 23102 24498 23154
rect 24558 23102 24610 23154
rect 25902 23102 25954 23154
rect 37662 23102 37714 23154
rect 11678 22990 11730 23042
rect 13806 22990 13858 23042
rect 14142 22990 14194 23042
rect 14478 22990 14530 23042
rect 17502 22990 17554 23042
rect 18846 22990 18898 23042
rect 24222 22990 24274 23042
rect 25342 22990 25394 23042
rect 26686 22990 26738 23042
rect 28814 22990 28866 23042
rect 18062 22878 18114 22930
rect 21646 22878 21698 22930
rect 23326 22878 23378 22930
rect 25454 22878 25506 22930
rect 25678 22878 25730 22930
rect 40014 22878 40066 22930
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 21534 22542 21586 22594
rect 10782 22430 10834 22482
rect 12910 22430 12962 22482
rect 19742 22430 19794 22482
rect 20302 22430 20354 22482
rect 25790 22430 25842 22482
rect 26350 22430 26402 22482
rect 10110 22318 10162 22370
rect 13918 22318 13970 22370
rect 14366 22318 14418 22370
rect 16270 22318 16322 22370
rect 16942 22318 16994 22370
rect 17390 22318 17442 22370
rect 19518 22318 19570 22370
rect 22878 22318 22930 22370
rect 23102 22318 23154 22370
rect 23438 22318 23490 22370
rect 23662 22318 23714 22370
rect 23886 22318 23938 22370
rect 24110 22318 24162 22370
rect 24334 22318 24386 22370
rect 24782 22318 24834 22370
rect 24894 22318 24946 22370
rect 25566 22318 25618 22370
rect 26574 22318 26626 22370
rect 26686 22318 26738 22370
rect 13582 22206 13634 22258
rect 15934 22206 15986 22258
rect 18510 22206 18562 22258
rect 21310 22206 21362 22258
rect 22542 22206 22594 22258
rect 25342 22206 25394 22258
rect 25902 22206 25954 22258
rect 26238 22206 26290 22258
rect 16830 22094 16882 22146
rect 17502 22094 17554 22146
rect 21870 22094 21922 22146
rect 22766 22094 22818 22146
rect 23774 22094 23826 22146
rect 24670 22094 24722 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 13134 21758 13186 21810
rect 15150 21758 15202 21810
rect 16158 21758 16210 21810
rect 16494 21758 16546 21810
rect 26014 21758 26066 21810
rect 14142 21646 14194 21698
rect 14814 21646 14866 21698
rect 15822 21646 15874 21698
rect 25230 21646 25282 21698
rect 25566 21646 25618 21698
rect 26238 21646 26290 21698
rect 14366 21534 14418 21586
rect 15598 21534 15650 21586
rect 17838 21534 17890 21586
rect 18174 21534 18226 21586
rect 23774 21534 23826 21586
rect 24334 21534 24386 21586
rect 24558 21534 24610 21586
rect 25790 21534 25842 21586
rect 26350 21534 26402 21586
rect 37662 21534 37714 21586
rect 21646 21422 21698 21474
rect 24446 21422 24498 21474
rect 25342 21422 25394 21474
rect 23998 21310 24050 21362
rect 40014 21310 40066 21362
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 19182 20974 19234 21026
rect 1934 20862 1986 20914
rect 18622 20862 18674 20914
rect 4174 20750 4226 20802
rect 14702 20750 14754 20802
rect 16942 20750 16994 20802
rect 17502 20750 17554 20802
rect 18062 20750 18114 20802
rect 18846 20750 18898 20802
rect 19630 20750 19682 20802
rect 20190 20750 20242 20802
rect 20526 20750 20578 20802
rect 20862 20750 20914 20802
rect 21646 20750 21698 20802
rect 25678 20638 25730 20690
rect 15038 20526 15090 20578
rect 18286 20526 18338 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 13134 20190 13186 20242
rect 15374 20190 15426 20242
rect 15598 20190 15650 20242
rect 14366 20078 14418 20130
rect 14478 20078 14530 20130
rect 15486 20078 15538 20130
rect 16270 20078 16322 20130
rect 18846 20078 18898 20130
rect 21310 20078 21362 20130
rect 22430 20078 22482 20130
rect 22654 20078 22706 20130
rect 22990 20078 23042 20130
rect 23774 20078 23826 20130
rect 23998 20078 24050 20130
rect 26462 20078 26514 20130
rect 4286 19966 4338 20018
rect 13918 19966 13970 20018
rect 14702 19966 14754 20018
rect 14926 19966 14978 20018
rect 16382 19966 16434 20018
rect 16606 19966 16658 20018
rect 16830 19966 16882 20018
rect 19406 19966 19458 20018
rect 19630 19966 19682 20018
rect 20526 19966 20578 20018
rect 22318 19966 22370 20018
rect 22878 19966 22930 20018
rect 24222 19966 24274 20018
rect 24670 19966 24722 20018
rect 25678 19966 25730 20018
rect 37662 19966 37714 20018
rect 11790 19854 11842 19906
rect 14366 19854 14418 19906
rect 16270 19854 16322 19906
rect 20190 19854 20242 19906
rect 20974 19854 21026 19906
rect 21758 19854 21810 19906
rect 24446 19854 24498 19906
rect 24558 19854 24610 19906
rect 25342 19854 25394 19906
rect 28590 19854 28642 19906
rect 1934 19742 1986 19794
rect 11902 19742 11954 19794
rect 22990 19742 23042 19794
rect 40014 19742 40066 19794
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 15150 19406 15202 19458
rect 1934 19294 1986 19346
rect 9886 19294 9938 19346
rect 12126 19294 12178 19346
rect 14814 19294 14866 19346
rect 17054 19294 17106 19346
rect 26462 19294 26514 19346
rect 28590 19294 28642 19346
rect 4286 19182 4338 19234
rect 12910 19182 12962 19234
rect 13694 19182 13746 19234
rect 19854 19182 19906 19234
rect 22206 19182 22258 19234
rect 23998 19182 24050 19234
rect 24446 19182 24498 19234
rect 24558 19182 24610 19234
rect 25678 19182 25730 19234
rect 13470 19070 13522 19122
rect 14926 18958 14978 19010
rect 21870 18958 21922 19010
rect 24222 18958 24274 19010
rect 24334 18958 24386 19010
rect 25342 18958 25394 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 12462 18622 12514 18674
rect 20414 18622 20466 18674
rect 20750 18622 20802 18674
rect 21086 18622 21138 18674
rect 21422 18622 21474 18674
rect 23998 18510 24050 18562
rect 24222 18510 24274 18562
rect 4286 18398 4338 18450
rect 12686 18398 12738 18450
rect 16606 18398 16658 18450
rect 17502 18398 17554 18450
rect 19630 18398 19682 18450
rect 23662 18398 23714 18450
rect 27918 18398 27970 18450
rect 28030 18398 28082 18450
rect 37662 18398 37714 18450
rect 13694 18286 13746 18338
rect 15822 18286 15874 18338
rect 19182 18286 19234 18338
rect 23774 18286 23826 18338
rect 1934 18174 1986 18226
rect 40014 18174 40066 18226
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 15374 17838 15426 17890
rect 20638 17838 20690 17890
rect 1934 17726 1986 17778
rect 15262 17726 15314 17778
rect 21310 17726 21362 17778
rect 23998 17726 24050 17778
rect 26126 17726 26178 17778
rect 4286 17614 4338 17666
rect 15038 17614 15090 17666
rect 15710 17614 15762 17666
rect 15934 17614 15986 17666
rect 16382 17614 16434 17666
rect 17614 17614 17666 17666
rect 18958 17614 19010 17666
rect 19294 17614 19346 17666
rect 19630 17614 19682 17666
rect 20078 17614 20130 17666
rect 20750 17614 20802 17666
rect 22206 17614 22258 17666
rect 23214 17614 23266 17666
rect 14254 17502 14306 17554
rect 14478 17502 14530 17554
rect 20302 17502 20354 17554
rect 21422 17502 21474 17554
rect 21646 17502 21698 17554
rect 14366 17390 14418 17442
rect 15822 17390 15874 17442
rect 17390 17390 17442 17442
rect 19182 17390 19234 17442
rect 21982 17390 22034 17442
rect 26574 17390 26626 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 14478 17054 14530 17106
rect 14590 17054 14642 17106
rect 15374 17054 15426 17106
rect 17614 17054 17666 17106
rect 13246 16942 13298 16994
rect 18734 16942 18786 16994
rect 22878 16942 22930 16994
rect 23214 16942 23266 16994
rect 24446 16942 24498 16994
rect 14030 16830 14082 16882
rect 14366 16830 14418 16882
rect 14926 16830 14978 16882
rect 17950 16830 18002 16882
rect 23326 16830 23378 16882
rect 11118 16718 11170 16770
rect 20862 16718 20914 16770
rect 23550 16718 23602 16770
rect 24222 16718 24274 16770
rect 24334 16718 24386 16770
rect 23774 16606 23826 16658
rect 23886 16606 23938 16658
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 18510 16270 18562 16322
rect 14254 16158 14306 16210
rect 19406 16158 19458 16210
rect 23662 16158 23714 16210
rect 25790 16158 25842 16210
rect 26238 16158 26290 16210
rect 22878 16046 22930 16098
rect 18398 15934 18450 15986
rect 19518 15934 19570 15986
rect 19742 15934 19794 15986
rect 16046 15822 16098 15874
rect 16382 15822 16434 15874
rect 18510 15822 18562 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 16606 15486 16658 15538
rect 17502 15486 17554 15538
rect 20190 15486 20242 15538
rect 20302 15486 20354 15538
rect 20638 15486 20690 15538
rect 21198 15486 21250 15538
rect 15374 15374 15426 15426
rect 22990 15374 23042 15426
rect 15150 15262 15202 15314
rect 15598 15262 15650 15314
rect 15822 15262 15874 15314
rect 19070 15262 19122 15314
rect 19406 15262 19458 15314
rect 19854 15262 19906 15314
rect 20414 15262 20466 15314
rect 22542 15262 22594 15314
rect 23102 15262 23154 15314
rect 14366 15150 14418 15202
rect 15262 15150 15314 15202
rect 19182 15150 19234 15202
rect 22766 15150 22818 15202
rect 14254 15038 14306 15090
rect 19518 15038 19570 15090
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 17054 14702 17106 14754
rect 22542 14702 22594 14754
rect 14254 14590 14306 14642
rect 16382 14590 16434 14642
rect 18622 14590 18674 14642
rect 20750 14590 20802 14642
rect 22094 14590 22146 14642
rect 13582 14478 13634 14530
rect 16830 14478 16882 14530
rect 17502 14478 17554 14530
rect 17838 14478 17890 14530
rect 22430 14478 22482 14530
rect 23998 14478 24050 14530
rect 17278 14366 17330 14418
rect 17054 14254 17106 14306
rect 22542 14254 22594 14306
rect 24222 14254 24274 14306
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 17390 13918 17442 13970
rect 25342 13918 25394 13970
rect 14702 13806 14754 13858
rect 18846 13806 18898 13858
rect 22542 13806 22594 13858
rect 13918 13694 13970 13746
rect 18062 13694 18114 13746
rect 21870 13694 21922 13746
rect 16830 13582 16882 13634
rect 17502 13582 17554 13634
rect 20974 13582 21026 13634
rect 24670 13582 24722 13634
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 20190 13134 20242 13186
rect 17166 13022 17218 13074
rect 17838 13022 17890 13074
rect 20302 12910 20354 12962
rect 23886 12686 23938 12738
rect 24222 12686 24274 12738
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 40238 12238 40290 12290
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 16718 5182 16770 5234
rect 24782 5182 24834 5234
rect 15710 5070 15762 5122
rect 23774 5070 23826 5122
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 20414 4286 20466 4338
rect 25454 4286 25506 4338
rect 21422 4062 21474 4114
rect 26238 4062 26290 4114
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 22094 3614 22146 3666
rect 25566 3614 25618 3666
rect 29374 3614 29426 3666
rect 17054 3502 17106 3554
rect 21086 3502 21138 3554
rect 24558 3502 24610 3554
rect 28590 3502 28642 3554
rect 18062 3278 18114 3330
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
<< metal2 >>
rect 19488 41200 19600 42000
rect 20832 41200 20944 42000
rect 24864 41200 24976 42000
rect 28896 41200 29008 42000
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 19516 37492 19572 41200
rect 20860 38276 20916 41200
rect 20860 38210 20916 38220
rect 22092 38276 22148 38286
rect 22092 38182 22148 38220
rect 24892 38276 24948 41200
rect 24892 38210 24948 38220
rect 26124 38276 26180 38286
rect 26124 38182 26180 38220
rect 21084 38050 21140 38062
rect 21084 37998 21086 38050
rect 21138 37998 21140 38050
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 19516 37426 19572 37436
rect 20748 37492 20804 37502
rect 20748 37398 20804 37436
rect 19740 37268 19796 37278
rect 19628 37266 19796 37268
rect 19628 37214 19742 37266
rect 19794 37214 19796 37266
rect 19628 37212 19796 37214
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 17052 28644 17108 28654
rect 4172 27636 4228 27646
rect 1932 27186 1988 27198
rect 1932 27134 1934 27186
rect 1986 27134 1988 27186
rect 1932 26292 1988 27134
rect 1932 26226 1988 26236
rect 4172 21476 4228 27580
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 4284 27076 4340 27086
rect 4284 26982 4340 27020
rect 12684 27076 12740 27086
rect 12684 26404 12740 27020
rect 17052 27074 17108 28588
rect 19628 28084 19684 37212
rect 19740 37202 19796 37212
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 21084 31948 21140 37998
rect 20748 31892 21140 31948
rect 25340 38050 25396 38062
rect 25340 37998 25342 38050
rect 25394 37998 25396 38050
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 20076 28644 20132 28654
rect 20076 28550 20132 28588
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 19628 28028 19908 28084
rect 18396 27748 18452 27758
rect 18396 27654 18452 27692
rect 19852 27188 19908 28028
rect 19628 27186 19908 27188
rect 19628 27134 19854 27186
rect 19906 27134 19908 27186
rect 19628 27132 19908 27134
rect 20524 27746 20580 27758
rect 20524 27694 20526 27746
rect 20578 27694 20580 27746
rect 20524 27188 20580 27694
rect 20748 27748 20804 31892
rect 21308 27860 21364 27870
rect 21868 27860 21924 27870
rect 21308 27858 22484 27860
rect 21308 27806 21310 27858
rect 21362 27806 21870 27858
rect 21922 27806 22484 27858
rect 21308 27804 22484 27806
rect 21308 27794 21364 27804
rect 21868 27794 21924 27804
rect 20636 27188 20692 27198
rect 20524 27186 20692 27188
rect 20524 27134 20638 27186
rect 20690 27134 20692 27186
rect 20524 27132 20692 27134
rect 17052 27022 17054 27074
rect 17106 27022 17108 27074
rect 14700 26962 14756 26974
rect 14700 26910 14702 26962
rect 14754 26910 14756 26962
rect 14588 26850 14644 26862
rect 14588 26798 14590 26850
rect 14642 26798 14644 26850
rect 14588 26516 14644 26798
rect 14700 26628 14756 26910
rect 15148 26964 15204 26974
rect 15148 26962 15428 26964
rect 15148 26910 15150 26962
rect 15202 26910 15428 26962
rect 15148 26908 15428 26910
rect 15148 26898 15204 26908
rect 14700 26562 14756 26572
rect 14812 26850 14868 26862
rect 14812 26798 14814 26850
rect 14866 26798 14868 26850
rect 14588 26450 14644 26460
rect 12684 26178 12740 26348
rect 14812 26402 14868 26798
rect 14812 26350 14814 26402
rect 14866 26350 14868 26402
rect 14812 26338 14868 26350
rect 14924 26850 14980 26862
rect 14924 26798 14926 26850
rect 14978 26798 14980 26850
rect 12684 26126 12686 26178
rect 12738 26126 12740 26178
rect 12684 26114 12740 26126
rect 13692 26292 13748 26302
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 13692 25506 13748 26236
rect 14924 25732 14980 26798
rect 14924 25666 14980 25676
rect 15260 26628 15316 26638
rect 13692 25454 13694 25506
rect 13746 25454 13748 25506
rect 13692 25442 13748 25454
rect 14364 25394 14420 25406
rect 14364 25342 14366 25394
rect 14418 25342 14420 25394
rect 13916 24500 13972 24510
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 13916 24162 13972 24444
rect 13916 24110 13918 24162
rect 13970 24110 13972 24162
rect 13916 24098 13972 24110
rect 13916 23940 13972 23950
rect 13916 23938 14308 23940
rect 13916 23886 13918 23938
rect 13970 23886 14308 23938
rect 13916 23884 14308 23886
rect 13916 23874 13972 23884
rect 13580 23826 13636 23838
rect 13580 23774 13582 23826
rect 13634 23774 13636 23826
rect 10892 23154 10948 23166
rect 10892 23102 10894 23154
rect 10946 23102 10948 23154
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 10780 22596 10836 22606
rect 10780 22482 10836 22540
rect 10780 22430 10782 22482
rect 10834 22430 10836 22482
rect 10780 22418 10836 22430
rect 10108 22372 10164 22382
rect 10108 22278 10164 22316
rect 10892 22372 10948 23102
rect 11676 23044 11732 23054
rect 11676 22950 11732 22988
rect 13580 23044 13636 23774
rect 10892 22306 10948 22316
rect 12908 22482 12964 22494
rect 12908 22430 12910 22482
rect 12962 22430 12964 22482
rect 12908 21700 12964 22430
rect 12908 21634 12964 21644
rect 13132 22372 13188 22382
rect 13132 21810 13188 22316
rect 13580 22258 13636 22988
rect 13804 23044 13860 23054
rect 14140 23044 14196 23054
rect 13804 22950 13860 22988
rect 13916 23042 14196 23044
rect 13916 22990 14142 23042
rect 14194 22990 14196 23042
rect 13916 22988 14196 22990
rect 13916 22370 13972 22988
rect 14140 22978 14196 22988
rect 13916 22318 13918 22370
rect 13970 22318 13972 22370
rect 13916 22306 13972 22318
rect 14252 22260 14308 23884
rect 14364 23604 14420 25342
rect 15260 24724 15316 26572
rect 15372 24946 15428 26908
rect 15820 26852 15876 26862
rect 17052 26852 17108 27022
rect 17724 27076 17780 27086
rect 17724 26982 17780 27020
rect 15484 26292 15540 26302
rect 15820 26292 15876 26796
rect 16940 26796 17052 26852
rect 15932 26516 15988 26526
rect 15932 26422 15988 26460
rect 16156 26404 16212 26414
rect 16156 26310 16212 26348
rect 15540 26236 15876 26292
rect 16268 26292 16324 26302
rect 16716 26292 16772 26302
rect 16268 26290 16772 26292
rect 16268 26238 16270 26290
rect 16322 26238 16718 26290
rect 16770 26238 16772 26290
rect 16268 26236 16772 26238
rect 15484 26198 15540 26236
rect 16268 26226 16324 26236
rect 16492 25618 16548 25630
rect 16492 25566 16494 25618
rect 16546 25566 16548 25618
rect 16492 25508 16548 25566
rect 16548 25452 16660 25508
rect 16492 25442 16548 25452
rect 15372 24894 15374 24946
rect 15426 24894 15428 24946
rect 15372 24882 15428 24894
rect 15484 24834 15540 24846
rect 15484 24782 15486 24834
rect 15538 24782 15540 24834
rect 15484 24724 15540 24782
rect 16380 24834 16436 24846
rect 16380 24782 16382 24834
rect 16434 24782 16436 24834
rect 15260 24668 15540 24724
rect 16156 24724 16212 24734
rect 15260 24500 15316 24510
rect 15260 24406 15316 24444
rect 15372 23828 15428 23838
rect 14364 23538 14420 23548
rect 15260 23772 15372 23828
rect 14812 23154 14868 23166
rect 14812 23102 14814 23154
rect 14866 23102 14868 23154
rect 14476 23044 14532 23054
rect 14476 22950 14532 22988
rect 14364 22372 14420 22382
rect 14364 22278 14420 22316
rect 14812 22372 14868 23102
rect 14812 22306 14868 22316
rect 13580 22206 13582 22258
rect 13634 22206 13636 22258
rect 13580 22194 13636 22206
rect 14140 22204 14252 22260
rect 13132 21758 13134 21810
rect 13186 21758 13188 21810
rect 4172 21410 4228 21420
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 1932 20914 1988 20926
rect 1932 20862 1934 20914
rect 1986 20862 1988 20914
rect 1932 20244 1988 20862
rect 1932 20178 1988 20188
rect 4172 20802 4228 20814
rect 4172 20750 4174 20802
rect 4226 20750 4228 20802
rect 1932 19796 1988 19806
rect 1932 19702 1988 19740
rect 1932 19346 1988 19358
rect 1932 19294 1934 19346
rect 1986 19294 1988 19346
rect 1932 18900 1988 19294
rect 4172 19348 4228 20750
rect 13132 20242 13188 21758
rect 14140 21698 14196 22204
rect 14252 22194 14308 22204
rect 14700 22260 14756 22270
rect 14140 21646 14142 21698
rect 14194 21646 14196 21698
rect 14140 21634 14196 21646
rect 14364 21700 14420 21710
rect 14364 21586 14420 21644
rect 14364 21534 14366 21586
rect 14418 21534 14420 21586
rect 14364 21522 14420 21534
rect 13132 20190 13134 20242
rect 13186 20190 13188 20242
rect 13132 20188 13188 20190
rect 12908 20132 13188 20188
rect 14700 20802 14756 22204
rect 15148 21812 15204 21822
rect 15148 21718 15204 21756
rect 14812 21700 14868 21710
rect 14812 21606 14868 21644
rect 14700 20750 14702 20802
rect 14754 20750 14756 20802
rect 14700 20188 14756 20750
rect 15036 20578 15092 20590
rect 15036 20526 15038 20578
rect 15090 20526 15092 20578
rect 14364 20132 14420 20142
rect 4284 20020 4340 20030
rect 4284 19926 4340 19964
rect 12460 20020 12516 20030
rect 11788 19908 11844 19918
rect 11788 19814 11844 19852
rect 11900 19796 11956 19806
rect 11900 19794 12180 19796
rect 11900 19742 11902 19794
rect 11954 19742 12180 19794
rect 11900 19740 12180 19742
rect 11900 19730 11956 19740
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 4172 19282 4228 19292
rect 9884 19348 9940 19358
rect 9884 19254 9940 19292
rect 12124 19346 12180 19740
rect 12124 19294 12126 19346
rect 12178 19294 12180 19346
rect 12124 19282 12180 19294
rect 4284 19236 4340 19246
rect 4284 19142 4340 19180
rect 1932 18834 1988 18844
rect 12460 18674 12516 19964
rect 12460 18622 12462 18674
rect 12514 18622 12516 18674
rect 12460 18610 12516 18622
rect 12684 19348 12740 19358
rect 4284 18452 4340 18462
rect 4284 18358 4340 18396
rect 12684 18450 12740 19292
rect 12684 18398 12686 18450
rect 12738 18398 12740 18450
rect 12684 18386 12740 18398
rect 12908 19234 12964 20132
rect 14364 20038 14420 20076
rect 14476 20130 14532 20142
rect 14700 20132 14980 20188
rect 14476 20078 14478 20130
rect 14530 20078 14532 20130
rect 13916 20018 13972 20030
rect 13916 19966 13918 20018
rect 13970 19966 13972 20018
rect 13692 19348 13748 19358
rect 12908 19182 12910 19234
rect 12962 19182 12964 19234
rect 12908 18452 12964 19182
rect 13468 19236 13524 19246
rect 13468 19122 13524 19180
rect 13692 19234 13748 19292
rect 13692 19182 13694 19234
rect 13746 19182 13748 19234
rect 13692 19170 13748 19182
rect 13468 19070 13470 19122
rect 13522 19070 13524 19122
rect 13468 19058 13524 19070
rect 13916 19012 13972 19966
rect 14364 19908 14420 19918
rect 14364 19814 14420 19852
rect 14476 19460 14532 20078
rect 14700 20018 14756 20030
rect 14700 19966 14702 20018
rect 14754 19966 14756 20018
rect 14700 19796 14756 19966
rect 14924 20018 14980 20132
rect 14924 19966 14926 20018
rect 14978 19966 14980 20018
rect 14924 19954 14980 19966
rect 15036 19796 15092 20526
rect 14700 19740 15092 19796
rect 15036 19572 15092 19740
rect 15036 19506 15092 19516
rect 15148 19908 15204 19918
rect 14140 19404 14532 19460
rect 15148 19458 15204 19852
rect 15148 19406 15150 19458
rect 15202 19406 15204 19458
rect 14140 19348 14196 19404
rect 15148 19394 15204 19406
rect 14812 19348 14868 19358
rect 14140 19282 14196 19292
rect 14252 19346 14868 19348
rect 14252 19294 14814 19346
rect 14866 19294 14868 19346
rect 14252 19292 14868 19294
rect 13916 18946 13972 18956
rect 12908 18386 12964 18396
rect 14028 18452 14084 18462
rect 13692 18340 13748 18350
rect 13692 18246 13748 18284
rect 1932 18228 1988 18238
rect 1932 18134 1988 18172
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 1932 17778 1988 17790
rect 1932 17726 1934 17778
rect 1986 17726 1988 17778
rect 1932 16884 1988 17726
rect 4284 17668 4340 17678
rect 4284 17574 4340 17612
rect 11116 17668 11172 17678
rect 1932 16818 1988 16828
rect 11116 17108 11172 17612
rect 11116 16770 11172 17052
rect 13244 17444 13300 17454
rect 13244 16994 13300 17388
rect 13244 16942 13246 16994
rect 13298 16942 13300 16994
rect 13244 16930 13300 16942
rect 14028 16884 14084 18396
rect 14252 17554 14308 19292
rect 14812 19282 14868 19292
rect 14924 19012 14980 19022
rect 14924 18918 14980 18956
rect 15260 18452 15316 23772
rect 15372 23762 15428 23772
rect 15372 23604 15428 23614
rect 15372 20242 15428 23548
rect 16156 23604 16212 24668
rect 15596 23044 15652 23054
rect 15596 21586 15652 22988
rect 15932 22372 15988 22382
rect 15932 22258 15988 22316
rect 15932 22206 15934 22258
rect 15986 22206 15988 22258
rect 15932 22194 15988 22206
rect 16156 21810 16212 23548
rect 16268 23154 16324 23166
rect 16268 23102 16270 23154
rect 16322 23102 16324 23154
rect 16268 23044 16324 23102
rect 16268 22370 16324 22988
rect 16268 22318 16270 22370
rect 16322 22318 16324 22370
rect 16268 22306 16324 22318
rect 16380 22372 16436 24782
rect 16604 24722 16660 25452
rect 16604 24670 16606 24722
rect 16658 24670 16660 24722
rect 16604 24658 16660 24670
rect 16716 23828 16772 26236
rect 16940 25620 16996 26796
rect 17052 26786 17108 26796
rect 18844 26628 18900 26638
rect 18844 26514 18900 26572
rect 18844 26462 18846 26514
rect 18898 26462 18900 26514
rect 18844 26450 18900 26462
rect 19068 26292 19124 26302
rect 19068 26198 19124 26236
rect 19628 26290 19684 27132
rect 19852 27122 19908 27132
rect 20636 27122 20692 27132
rect 20188 26962 20244 26974
rect 20188 26910 20190 26962
rect 20242 26910 20244 26962
rect 20188 26740 20244 26910
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20188 26674 20244 26684
rect 20300 26964 20356 26974
rect 19836 26618 20100 26628
rect 19852 26516 19908 26526
rect 20300 26516 20356 26908
rect 19852 26514 20356 26516
rect 19852 26462 19854 26514
rect 19906 26462 20356 26514
rect 19852 26460 20356 26462
rect 20412 26962 20468 26974
rect 20748 26964 20804 27692
rect 20860 27188 20916 27198
rect 20860 27074 20916 27132
rect 21980 27188 22036 27198
rect 20860 27022 20862 27074
rect 20914 27022 20916 27074
rect 20860 27010 20916 27022
rect 21644 27074 21700 27086
rect 21644 27022 21646 27074
rect 21698 27022 21700 27074
rect 20412 26910 20414 26962
rect 20466 26910 20468 26962
rect 20412 26852 20468 26910
rect 19852 26450 19908 26460
rect 19628 26238 19630 26290
rect 19682 26238 19684 26290
rect 19628 26226 19684 26238
rect 19740 26292 19796 26302
rect 19964 26292 20020 26302
rect 17500 25732 17556 25742
rect 16940 25618 17108 25620
rect 16940 25566 16942 25618
rect 16994 25566 17108 25618
rect 16940 25564 17108 25566
rect 16940 25554 16996 25564
rect 16716 23762 16772 23772
rect 16604 23380 16660 23390
rect 16604 23286 16660 23324
rect 16380 22306 16436 22316
rect 16940 22370 16996 22382
rect 16940 22318 16942 22370
rect 16994 22318 16996 22370
rect 16156 21758 16158 21810
rect 16210 21758 16212 21810
rect 15596 21534 15598 21586
rect 15650 21534 15652 21586
rect 15596 21522 15652 21534
rect 15820 21700 15876 21710
rect 15820 20356 15876 21644
rect 15372 20190 15374 20242
rect 15426 20190 15428 20242
rect 15372 20178 15428 20190
rect 15596 20300 15988 20356
rect 15596 20242 15652 20300
rect 15596 20190 15598 20242
rect 15650 20190 15652 20242
rect 15596 20178 15652 20190
rect 15484 20132 15540 20142
rect 15484 20038 15540 20076
rect 15148 18396 15316 18452
rect 15036 17666 15092 17678
rect 15036 17614 15038 17666
rect 15090 17614 15092 17666
rect 14252 17502 14254 17554
rect 14306 17502 14308 17554
rect 14252 17490 14308 17502
rect 14476 17554 14532 17566
rect 14476 17502 14478 17554
rect 14530 17502 14532 17554
rect 14364 17444 14420 17454
rect 14364 17350 14420 17388
rect 14476 17106 14532 17502
rect 14476 17054 14478 17106
rect 14530 17054 14532 17106
rect 14476 17042 14532 17054
rect 14588 17108 14644 17118
rect 14588 17014 14644 17052
rect 11116 16718 11118 16770
rect 11170 16718 11172 16770
rect 11116 16706 11172 16718
rect 13580 16882 14308 16884
rect 13580 16830 14030 16882
rect 14082 16830 14308 16882
rect 13580 16828 14308 16830
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 13580 14532 13636 16828
rect 14028 16818 14084 16828
rect 14252 16210 14308 16828
rect 14364 16882 14420 16894
rect 14364 16830 14366 16882
rect 14418 16830 14420 16882
rect 14364 16772 14420 16830
rect 14924 16884 14980 16894
rect 14924 16790 14980 16828
rect 14364 16706 14420 16716
rect 15036 16772 15092 17614
rect 15148 17108 15204 18396
rect 15820 18340 15876 18350
rect 15260 18338 15876 18340
rect 15260 18286 15822 18338
rect 15874 18286 15876 18338
rect 15260 18284 15876 18286
rect 15260 17778 15316 18284
rect 15820 18274 15876 18284
rect 15932 18116 15988 20300
rect 15708 18060 15988 18116
rect 15372 17892 15428 17902
rect 15596 17892 15652 17902
rect 15372 17890 15596 17892
rect 15372 17838 15374 17890
rect 15426 17838 15596 17890
rect 15372 17836 15596 17838
rect 15372 17826 15428 17836
rect 15596 17826 15652 17836
rect 15260 17726 15262 17778
rect 15314 17726 15316 17778
rect 15260 17714 15316 17726
rect 15708 17666 15764 18060
rect 15708 17614 15710 17666
rect 15762 17614 15764 17666
rect 15708 17602 15764 17614
rect 15932 17668 15988 17678
rect 16156 17668 16212 21758
rect 16492 22148 16548 22158
rect 16492 21810 16548 22092
rect 16828 22146 16884 22158
rect 16828 22094 16830 22146
rect 16882 22094 16884 22146
rect 16828 21924 16884 22094
rect 16828 21858 16884 21868
rect 16492 21758 16494 21810
rect 16546 21758 16548 21810
rect 16492 21746 16548 21758
rect 16940 21812 16996 22318
rect 16940 20802 16996 21756
rect 16940 20750 16942 20802
rect 16994 20750 16996 20802
rect 16940 20738 16996 20750
rect 16268 20132 16324 20142
rect 16268 20038 16324 20076
rect 16380 20018 16436 20030
rect 16380 19966 16382 20018
rect 16434 19966 16436 20018
rect 16268 19906 16324 19918
rect 16268 19854 16270 19906
rect 16322 19854 16324 19906
rect 16268 17892 16324 19854
rect 16380 18228 16436 19966
rect 16604 20020 16660 20030
rect 16604 19926 16660 19964
rect 16828 20018 16884 20030
rect 16828 19966 16830 20018
rect 16882 19966 16884 20018
rect 16828 19908 16884 19966
rect 16828 19842 16884 19852
rect 17052 19348 17108 25564
rect 17276 25508 17332 25518
rect 17276 25414 17332 25452
rect 17388 25172 17444 25182
rect 17388 24834 17444 25116
rect 17500 24946 17556 25676
rect 19740 25620 19796 26236
rect 19516 25564 19796 25620
rect 19852 26290 20020 26292
rect 19852 26238 19966 26290
rect 20018 26238 20020 26290
rect 19852 26236 20020 26238
rect 17836 25508 17892 25518
rect 18172 25508 18228 25518
rect 17836 25506 18172 25508
rect 17836 25454 17838 25506
rect 17890 25454 18172 25506
rect 17836 25452 18172 25454
rect 17836 25442 17892 25452
rect 17500 24894 17502 24946
rect 17554 24894 17556 24946
rect 17500 24882 17556 24894
rect 17388 24782 17390 24834
rect 17442 24782 17444 24834
rect 17388 24770 17444 24782
rect 17612 24724 17668 24734
rect 17612 24630 17668 24668
rect 17948 24722 18004 24734
rect 17948 24670 17950 24722
rect 18002 24670 18004 24722
rect 17948 24052 18004 24670
rect 17948 23986 18004 23996
rect 18060 24050 18116 24062
rect 18060 23998 18062 24050
rect 18114 23998 18116 24050
rect 18060 23604 18116 23998
rect 17612 23548 18116 23604
rect 18172 23714 18228 25452
rect 19292 25508 19348 25518
rect 19292 25414 19348 25452
rect 18844 25172 18900 25182
rect 18732 23938 18788 23950
rect 18732 23886 18734 23938
rect 18786 23886 18788 23938
rect 18172 23662 18174 23714
rect 18226 23662 18228 23714
rect 17500 23044 17556 23054
rect 17388 23042 17556 23044
rect 17388 22990 17502 23042
rect 17554 22990 17556 23042
rect 17388 22988 17556 22990
rect 17388 22372 17444 22988
rect 17500 22978 17556 22988
rect 17388 22278 17444 22316
rect 17500 22148 17556 22158
rect 17500 22054 17556 22092
rect 17500 20804 17556 20814
rect 17500 20132 17556 20748
rect 17612 20468 17668 23548
rect 18172 23492 18228 23662
rect 18172 23426 18228 23436
rect 18396 23826 18452 23838
rect 18396 23774 18398 23826
rect 18450 23774 18452 23826
rect 17724 23380 17780 23390
rect 17724 23154 17780 23324
rect 18396 23380 18452 23774
rect 18396 23314 18452 23324
rect 17724 23102 17726 23154
rect 17778 23102 17780 23154
rect 17724 23090 17780 23102
rect 18396 23154 18452 23166
rect 18620 23156 18676 23166
rect 18396 23102 18398 23154
rect 18450 23102 18452 23154
rect 18060 22932 18116 22942
rect 18116 22876 18340 22932
rect 18060 22838 18116 22876
rect 17724 22708 17780 22718
rect 17724 21924 17780 22652
rect 17724 20580 17780 21868
rect 17836 21588 17892 21598
rect 18172 21588 18228 21598
rect 17836 21586 18228 21588
rect 17836 21534 17838 21586
rect 17890 21534 18174 21586
rect 18226 21534 18228 21586
rect 17836 21532 18228 21534
rect 17836 21476 17892 21532
rect 18172 21522 18228 21532
rect 17836 21410 17892 21420
rect 18060 20804 18116 20814
rect 18284 20804 18340 22876
rect 18396 22708 18452 23102
rect 18396 22642 18452 22652
rect 18508 23154 18676 23156
rect 18508 23102 18622 23154
rect 18674 23102 18676 23154
rect 18508 23100 18676 23102
rect 18508 22484 18564 23100
rect 18620 23090 18676 23100
rect 18060 20802 18340 20804
rect 18060 20750 18062 20802
rect 18114 20750 18340 20802
rect 18060 20748 18340 20750
rect 18396 22428 18564 22484
rect 18732 22484 18788 23886
rect 18844 23268 18900 25116
rect 19180 24948 19236 24958
rect 19180 24854 19236 24892
rect 19068 24612 19124 24622
rect 19068 24610 19236 24612
rect 19068 24558 19070 24610
rect 19122 24558 19236 24610
rect 19068 24556 19236 24558
rect 19068 24546 19124 24556
rect 18956 24052 19012 24062
rect 18956 23958 19012 23996
rect 19068 23826 19124 23838
rect 19068 23774 19070 23826
rect 19122 23774 19124 23826
rect 18844 23212 19012 23268
rect 18844 23042 18900 23054
rect 18844 22990 18846 23042
rect 18898 22990 18900 23042
rect 18844 22596 18900 22990
rect 18844 22530 18900 22540
rect 18060 20738 18116 20748
rect 18284 20580 18340 20590
rect 18396 20580 18452 22428
rect 18620 22372 18676 22382
rect 18508 22260 18564 22270
rect 18508 22166 18564 22204
rect 18620 20914 18676 22316
rect 18732 22148 18788 22428
rect 18956 22372 19012 23212
rect 19068 23156 19124 23774
rect 19180 23380 19236 24556
rect 19516 24052 19572 25564
rect 19628 25396 19684 25406
rect 19628 25302 19684 25340
rect 19852 25284 19908 26236
rect 19964 26226 20020 26236
rect 20188 26292 20244 26302
rect 20188 25618 20244 26236
rect 20188 25566 20190 25618
rect 20242 25566 20244 25618
rect 20188 25554 20244 25566
rect 19964 25508 20020 25518
rect 19964 25414 20020 25452
rect 19852 25218 19908 25228
rect 20300 25394 20356 25406
rect 20300 25342 20302 25394
rect 20354 25342 20356 25394
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 20300 24948 20356 25342
rect 20412 25396 20468 26796
rect 20636 26908 20804 26964
rect 21308 26964 21364 26974
rect 20636 26290 20692 26908
rect 21308 26870 21364 26908
rect 21644 26852 21700 27022
rect 21756 27076 21812 27086
rect 21756 26982 21812 27020
rect 21980 27074 22036 27132
rect 21980 27022 21982 27074
rect 22034 27022 22036 27074
rect 21980 26964 22036 27022
rect 22428 27076 22484 27804
rect 25340 27186 25396 37998
rect 28924 37940 28980 41200
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 29148 37940 29204 37950
rect 28924 37938 29204 37940
rect 28924 37886 29150 37938
rect 29202 37886 29204 37938
rect 28924 37884 29204 37886
rect 29148 37874 29204 37884
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 25340 27134 25342 27186
rect 25394 27134 25396 27186
rect 22428 26982 22484 27020
rect 25228 27076 25284 27086
rect 23212 26964 23268 26974
rect 21980 26898 22036 26908
rect 22988 26962 23268 26964
rect 22988 26910 23214 26962
rect 23266 26910 23268 26962
rect 22988 26908 23268 26910
rect 21644 26786 21700 26796
rect 20860 26740 20916 26750
rect 20860 26514 20916 26684
rect 20860 26462 20862 26514
rect 20914 26462 20916 26514
rect 20860 26450 20916 26462
rect 22988 26514 23044 26908
rect 23212 26898 23268 26908
rect 23996 26964 24052 26974
rect 22988 26462 22990 26514
rect 23042 26462 23044 26514
rect 22988 26450 23044 26462
rect 20748 26404 20804 26414
rect 20748 26310 20804 26348
rect 23996 26402 24052 26908
rect 25116 26964 25172 26974
rect 24444 26516 24500 26526
rect 24444 26422 24500 26460
rect 23996 26350 23998 26402
rect 24050 26350 24052 26402
rect 20636 26238 20638 26290
rect 20690 26238 20692 26290
rect 20636 26226 20692 26238
rect 20972 26292 21028 26302
rect 20972 26198 21028 26236
rect 21196 26290 21252 26302
rect 21196 26238 21198 26290
rect 21250 26238 21252 26290
rect 20412 25330 20468 25340
rect 20972 25732 21028 25742
rect 20300 24882 20356 24892
rect 20860 24948 20916 24958
rect 20412 24724 20468 24734
rect 20300 24722 20468 24724
rect 20300 24670 20414 24722
rect 20466 24670 20468 24722
rect 20300 24668 20468 24670
rect 19852 24500 19908 24510
rect 19628 24052 19684 24062
rect 19516 24050 19684 24052
rect 19516 23998 19630 24050
rect 19682 23998 19684 24050
rect 19516 23996 19684 23998
rect 19628 23986 19684 23996
rect 19852 23938 19908 24444
rect 19852 23886 19854 23938
rect 19906 23886 19908 23938
rect 19852 23874 19908 23886
rect 19180 23314 19236 23324
rect 19516 23826 19572 23838
rect 19516 23774 19518 23826
rect 19570 23774 19572 23826
rect 19404 23268 19460 23278
rect 19068 23154 19236 23156
rect 19068 23102 19070 23154
rect 19122 23102 19236 23154
rect 19068 23100 19236 23102
rect 19068 23090 19124 23100
rect 18732 22082 18788 22092
rect 18844 22316 19012 22372
rect 18844 21028 18900 22316
rect 18620 20862 18622 20914
rect 18674 20862 18676 20914
rect 18620 20850 18676 20862
rect 18732 20972 18900 21028
rect 19180 21026 19236 23100
rect 19180 20974 19182 21026
rect 19234 20974 19236 21026
rect 17724 20524 18116 20580
rect 17612 20412 17780 20468
rect 17556 20076 17668 20132
rect 17500 20066 17556 20076
rect 16828 19346 17108 19348
rect 16828 19294 17054 19346
rect 17106 19294 17108 19346
rect 16828 19292 17108 19294
rect 16604 18452 16660 18462
rect 16828 18452 16884 19292
rect 17052 19282 17108 19292
rect 16660 18396 16884 18452
rect 17500 18452 17556 18462
rect 16604 18358 16660 18396
rect 16380 18162 16436 18172
rect 16268 17826 16324 17836
rect 15932 17666 16212 17668
rect 15932 17614 15934 17666
rect 15986 17614 16212 17666
rect 15932 17612 16212 17614
rect 16380 17666 16436 17678
rect 16380 17614 16382 17666
rect 16434 17614 16436 17666
rect 15932 17602 15988 17612
rect 15820 17442 15876 17454
rect 15820 17390 15822 17442
rect 15874 17390 15876 17442
rect 15372 17108 15428 17118
rect 15148 17106 15428 17108
rect 15148 17054 15374 17106
rect 15426 17054 15428 17106
rect 15148 17052 15428 17054
rect 15148 16884 15204 17052
rect 15372 17042 15428 17052
rect 15148 16818 15204 16828
rect 14252 16158 14254 16210
rect 14306 16158 14308 16210
rect 14252 16146 14308 16158
rect 15036 15316 15092 16716
rect 15372 15426 15428 15438
rect 15372 15374 15374 15426
rect 15426 15374 15428 15426
rect 15148 15316 15204 15326
rect 15036 15260 15148 15316
rect 15148 15222 15204 15260
rect 14364 15204 14420 15214
rect 14364 15110 14420 15148
rect 15260 15204 15316 15242
rect 15260 15138 15316 15148
rect 14252 15090 14308 15102
rect 14252 15038 14254 15090
rect 14306 15038 14308 15090
rect 14252 14642 14308 15038
rect 14252 14590 14254 14642
rect 14306 14590 14308 14642
rect 14252 14578 14308 14590
rect 15372 14644 15428 15374
rect 15596 15314 15652 15326
rect 15596 15262 15598 15314
rect 15650 15262 15652 15314
rect 15596 15204 15652 15262
rect 15820 15314 15876 17390
rect 15820 15262 15822 15314
rect 15874 15262 15876 15314
rect 15820 15250 15876 15262
rect 16044 15874 16100 15886
rect 16044 15822 16046 15874
rect 16098 15822 16100 15874
rect 16044 15316 16100 15822
rect 16380 15874 16436 17614
rect 17388 17442 17444 17454
rect 17388 17390 17390 17442
rect 17442 17390 17444 17442
rect 17388 15988 17444 17390
rect 17388 15922 17444 15932
rect 17500 17108 17556 18396
rect 17612 17666 17668 20076
rect 17724 19908 17780 20412
rect 17724 19842 17780 19852
rect 17612 17614 17614 17666
rect 17666 17614 17668 17666
rect 17612 17602 17668 17614
rect 17612 17108 17668 17118
rect 17500 17106 18004 17108
rect 17500 17054 17614 17106
rect 17666 17054 18004 17106
rect 17500 17052 18004 17054
rect 16380 15822 16382 15874
rect 16434 15822 16436 15874
rect 16380 15540 16436 15822
rect 16380 15474 16436 15484
rect 16604 15540 16660 15550
rect 17500 15540 17556 17052
rect 17612 17042 17668 17052
rect 17948 16882 18004 17052
rect 17948 16830 17950 16882
rect 18002 16830 18004 16882
rect 17948 16818 18004 16830
rect 16604 15538 17892 15540
rect 16604 15486 16606 15538
rect 16658 15486 17502 15538
rect 17554 15486 17892 15538
rect 16604 15484 17892 15486
rect 16604 15474 16660 15484
rect 17500 15474 17556 15484
rect 16044 15250 16100 15260
rect 16828 15316 16884 15326
rect 15596 15138 15652 15148
rect 16380 14644 16436 14654
rect 15372 14642 16436 14644
rect 15372 14590 16382 14642
rect 16434 14590 16436 14642
rect 15372 14588 16436 14590
rect 13580 14530 13972 14532
rect 13580 14478 13582 14530
rect 13634 14478 13972 14530
rect 13580 14476 13972 14478
rect 13580 14466 13636 14476
rect 13916 13746 13972 14476
rect 14700 14308 14756 14318
rect 14700 13858 14756 14252
rect 14700 13806 14702 13858
rect 14754 13806 14756 13858
rect 14700 13794 14756 13806
rect 13916 13694 13918 13746
rect 13970 13694 13972 13746
rect 13916 13682 13972 13694
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 16380 8428 16436 14588
rect 16828 14530 16884 15260
rect 17500 15204 17556 15214
rect 17052 15092 17108 15102
rect 17052 14754 17108 15036
rect 17052 14702 17054 14754
rect 17106 14702 17108 14754
rect 17052 14690 17108 14702
rect 16828 14478 16830 14530
rect 16882 14478 16884 14530
rect 16828 14466 16884 14478
rect 17500 14530 17556 15148
rect 17500 14478 17502 14530
rect 17554 14478 17556 14530
rect 17500 14466 17556 14478
rect 17836 14532 17892 15484
rect 18060 15148 18116 20524
rect 18284 20578 18564 20580
rect 18284 20526 18286 20578
rect 18338 20526 18564 20578
rect 18284 20524 18564 20526
rect 18284 20514 18340 20524
rect 18508 18452 18564 20524
rect 18732 20132 18788 20972
rect 19180 20962 19236 20974
rect 18844 20804 18900 20814
rect 19404 20804 19460 23212
rect 19516 22708 19572 23774
rect 20300 23714 20356 24668
rect 20412 24658 20468 24668
rect 20860 24722 20916 24892
rect 20972 24834 21028 25676
rect 21196 25284 21252 26238
rect 22652 26290 22708 26302
rect 22652 26238 22654 26290
rect 22706 26238 22708 26290
rect 22652 25732 22708 26238
rect 22652 25666 22708 25676
rect 22876 26290 22932 26302
rect 22876 26238 22878 26290
rect 22930 26238 22932 26290
rect 22876 25508 22932 26238
rect 23100 26292 23156 26302
rect 23100 26198 23156 26236
rect 23212 26290 23268 26302
rect 23212 26238 23214 26290
rect 23266 26238 23268 26290
rect 23100 25620 23156 25630
rect 23212 25620 23268 26238
rect 23660 26290 23716 26302
rect 23660 26238 23662 26290
rect 23714 26238 23716 26290
rect 23660 25732 23716 26238
rect 23660 25666 23716 25676
rect 23100 25618 23268 25620
rect 23100 25566 23102 25618
rect 23154 25566 23268 25618
rect 23100 25564 23268 25566
rect 23100 25554 23156 25564
rect 22540 25452 22932 25508
rect 22540 25396 22596 25452
rect 21196 25218 21252 25228
rect 21980 25284 22036 25294
rect 21980 25190 22036 25228
rect 22316 25284 22372 25294
rect 22316 25282 22484 25284
rect 22316 25230 22318 25282
rect 22370 25230 22484 25282
rect 22316 25228 22484 25230
rect 22316 25218 22372 25228
rect 22428 24836 22484 25228
rect 22540 24946 22596 25340
rect 23772 25396 23828 25406
rect 22540 24894 22542 24946
rect 22594 24894 22596 24946
rect 22540 24882 22596 24894
rect 22764 25282 22820 25294
rect 22764 25230 22766 25282
rect 22818 25230 22820 25282
rect 22764 24946 22820 25230
rect 22988 25284 23044 25294
rect 22988 25190 23044 25228
rect 23212 25282 23268 25294
rect 23212 25230 23214 25282
rect 23266 25230 23268 25282
rect 22764 24894 22766 24946
rect 22818 24894 22820 24946
rect 22764 24882 22820 24894
rect 20972 24782 20974 24834
rect 21026 24782 21028 24834
rect 20972 24770 21028 24782
rect 22204 24834 22484 24836
rect 22204 24782 22430 24834
rect 22482 24782 22484 24834
rect 22204 24780 22484 24782
rect 20860 24670 20862 24722
rect 20914 24670 20916 24722
rect 20860 24658 20916 24670
rect 20636 24500 20692 24510
rect 20300 23662 20302 23714
rect 20354 23662 20356 23714
rect 19836 23548 20100 23558
rect 19516 22642 19572 22652
rect 19628 23492 19684 23502
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 19628 22484 19684 23436
rect 20188 23380 20244 23390
rect 19740 23156 19796 23166
rect 19740 23154 19908 23156
rect 19740 23102 19742 23154
rect 19794 23102 19908 23154
rect 19740 23100 19908 23102
rect 19740 23090 19796 23100
rect 19740 22484 19796 22494
rect 19628 22482 19796 22484
rect 19628 22430 19742 22482
rect 19794 22430 19796 22482
rect 19628 22428 19796 22430
rect 19740 22418 19796 22428
rect 19516 22372 19572 22382
rect 19516 22278 19572 22316
rect 19852 22148 19908 23100
rect 20188 23154 20244 23324
rect 20300 23268 20356 23662
rect 20524 24444 20636 24500
rect 20300 23202 20356 23212
rect 20412 23266 20468 23278
rect 20412 23214 20414 23266
rect 20466 23214 20468 23266
rect 20188 23102 20190 23154
rect 20242 23102 20244 23154
rect 20188 23090 20244 23102
rect 20300 22596 20356 22606
rect 20300 22482 20356 22540
rect 20300 22430 20302 22482
rect 20354 22430 20356 22482
rect 20300 22418 20356 22430
rect 20412 22148 20468 23214
rect 19628 22092 19908 22148
rect 20188 22092 20412 22148
rect 19628 21924 19684 22092
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 19628 21858 19684 21868
rect 18844 20802 19460 20804
rect 18844 20750 18846 20802
rect 18898 20750 19460 20802
rect 18844 20748 19460 20750
rect 19628 20804 19684 20814
rect 18844 20738 18900 20748
rect 19404 20580 19460 20590
rect 18844 20132 18900 20142
rect 18732 20130 18900 20132
rect 18732 20078 18846 20130
rect 18898 20078 18900 20130
rect 18732 20076 18900 20078
rect 18732 20020 18788 20076
rect 18844 20066 18900 20076
rect 19404 20020 19460 20524
rect 18732 19954 18788 19964
rect 19180 20018 19460 20020
rect 19180 19966 19406 20018
rect 19458 19966 19460 20018
rect 19180 19964 19460 19966
rect 18508 18386 18564 18396
rect 19180 18338 19236 19964
rect 19404 19954 19460 19964
rect 19628 20018 19684 20748
rect 20188 20802 20244 22092
rect 20412 22082 20468 22092
rect 20188 20750 20190 20802
rect 20242 20750 20244 20802
rect 20188 20738 20244 20750
rect 20300 21812 20356 21822
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 19628 19966 19630 20018
rect 19682 19966 19684 20018
rect 19628 19954 19684 19966
rect 19852 20244 19908 20254
rect 19852 19234 19908 20188
rect 20188 19908 20244 19918
rect 20300 19908 20356 21756
rect 20524 20802 20580 24444
rect 20636 24406 20692 24444
rect 20636 23828 20692 23838
rect 20636 23734 20692 23772
rect 21308 23268 21364 23278
rect 21532 23268 21588 23278
rect 21308 23174 21364 23212
rect 21420 23266 21588 23268
rect 21420 23214 21534 23266
rect 21586 23214 21588 23266
rect 21420 23212 21588 23214
rect 21420 22372 21476 23212
rect 21532 23202 21588 23212
rect 21532 22932 21588 22942
rect 21532 22594 21588 22876
rect 21532 22542 21534 22594
rect 21586 22542 21588 22594
rect 21532 22530 21588 22542
rect 21644 22930 21700 22942
rect 21644 22878 21646 22930
rect 21698 22878 21700 22930
rect 21308 22260 21364 22270
rect 21420 22260 21476 22316
rect 21644 22372 21700 22878
rect 21644 22306 21700 22316
rect 21308 22258 21476 22260
rect 21308 22206 21310 22258
rect 21362 22206 21476 22258
rect 21308 22204 21476 22206
rect 21308 22194 21364 22204
rect 20524 20750 20526 20802
rect 20578 20750 20580 20802
rect 20524 20580 20580 20750
rect 20860 22036 20916 22046
rect 20860 20802 20916 21980
rect 20860 20750 20862 20802
rect 20914 20750 20916 20802
rect 20860 20738 20916 20750
rect 20524 20514 20580 20524
rect 21308 20132 21364 20142
rect 20524 20130 21364 20132
rect 20524 20078 21310 20130
rect 21362 20078 21364 20130
rect 20524 20076 21364 20078
rect 20524 20018 20580 20076
rect 20524 19966 20526 20018
rect 20578 19966 20580 20018
rect 20524 19954 20580 19966
rect 20188 19906 20356 19908
rect 20188 19854 20190 19906
rect 20242 19854 20356 19906
rect 20188 19852 20356 19854
rect 20188 19842 20244 19852
rect 19852 19182 19854 19234
rect 19906 19182 19908 19234
rect 19852 19170 19908 19182
rect 20412 19796 20468 19806
rect 20412 19012 20468 19740
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 20412 18674 20468 18956
rect 20748 18676 20804 20076
rect 21308 20066 21364 20076
rect 20972 19908 21028 19918
rect 21420 19908 21476 22204
rect 21868 22146 21924 22158
rect 21868 22094 21870 22146
rect 21922 22094 21924 22146
rect 21644 21474 21700 21486
rect 21644 21422 21646 21474
rect 21698 21422 21700 21474
rect 21644 20802 21700 21422
rect 21644 20750 21646 20802
rect 21698 20750 21700 20802
rect 21644 20244 21700 20750
rect 21868 20804 21924 22094
rect 21868 20738 21924 20748
rect 21644 20178 21700 20188
rect 21756 19908 21812 19918
rect 21420 19906 21812 19908
rect 21420 19854 21758 19906
rect 21810 19854 21812 19906
rect 21420 19852 21812 19854
rect 20972 19814 21028 19852
rect 21756 19842 21812 19852
rect 22204 19908 22260 24780
rect 22428 24770 22484 24780
rect 23212 23380 23268 25230
rect 23772 24162 23828 25340
rect 23772 24110 23774 24162
rect 23826 24110 23828 24162
rect 23772 24098 23828 24110
rect 23884 25284 23940 25294
rect 23436 24052 23492 24062
rect 23436 23958 23492 23996
rect 22764 23324 23268 23380
rect 23660 23714 23716 23726
rect 23660 23662 23662 23714
rect 23714 23662 23716 23714
rect 22652 22372 22708 22382
rect 22540 22258 22596 22270
rect 22540 22206 22542 22258
rect 22594 22206 22596 22258
rect 22540 22148 22596 22206
rect 22540 22082 22596 22092
rect 22652 21812 22708 22316
rect 22540 21756 22708 21812
rect 22764 22146 22820 23324
rect 22988 23154 23044 23166
rect 22988 23102 22990 23154
rect 23042 23102 23044 23154
rect 22876 22484 22932 22494
rect 22988 22484 23044 23102
rect 22932 22428 23044 22484
rect 23100 23156 23156 23166
rect 22876 22370 22932 22428
rect 22876 22318 22878 22370
rect 22930 22318 22932 22370
rect 22876 22306 22932 22318
rect 23100 22372 23156 23100
rect 23212 23156 23268 23166
rect 23212 23154 23604 23156
rect 23212 23102 23214 23154
rect 23266 23102 23604 23154
rect 23212 23100 23604 23102
rect 23212 23090 23268 23100
rect 23324 22930 23380 22942
rect 23324 22878 23326 22930
rect 23378 22878 23380 22930
rect 23100 22370 23268 22372
rect 23100 22318 23102 22370
rect 23154 22318 23268 22370
rect 23100 22316 23268 22318
rect 23100 22306 23156 22316
rect 22764 22094 22766 22146
rect 22818 22094 22820 22146
rect 22428 20132 22484 20142
rect 21420 19236 21476 19246
rect 21084 18676 21140 18686
rect 20412 18622 20414 18674
rect 20466 18622 20468 18674
rect 20412 18610 20468 18622
rect 20524 18674 21140 18676
rect 20524 18622 20750 18674
rect 20802 18622 21086 18674
rect 21138 18622 21140 18674
rect 20524 18620 21140 18622
rect 19180 18286 19182 18338
rect 19234 18286 19236 18338
rect 19180 18274 19236 18286
rect 19292 18452 19348 18462
rect 18956 17668 19012 17678
rect 18508 17666 19012 17668
rect 18508 17614 18958 17666
rect 19010 17614 19012 17666
rect 18508 17612 19012 17614
rect 18508 16322 18564 17612
rect 18956 17602 19012 17612
rect 19292 17666 19348 18396
rect 19628 18452 19684 18462
rect 19628 18358 19684 18396
rect 20524 18340 20580 18620
rect 20748 18610 20804 18620
rect 21084 18610 21140 18620
rect 21420 18674 21476 19180
rect 22204 19234 22260 19852
rect 22204 19182 22206 19234
rect 22258 19182 22260 19234
rect 22204 19170 22260 19182
rect 22316 20018 22372 20030
rect 22316 19966 22318 20018
rect 22370 19966 22372 20018
rect 21420 18622 21422 18674
rect 21474 18622 21476 18674
rect 20300 18284 20580 18340
rect 20636 18452 20692 18462
rect 19628 17780 19684 17790
rect 19628 17668 19684 17724
rect 19292 17614 19294 17666
rect 19346 17614 19348 17666
rect 19292 17556 19348 17614
rect 19292 17490 19348 17500
rect 19516 17666 19684 17668
rect 19516 17614 19630 17666
rect 19682 17614 19684 17666
rect 19516 17612 19684 17614
rect 19180 17442 19236 17454
rect 19180 17390 19182 17442
rect 19234 17390 19236 17442
rect 19180 17108 19236 17390
rect 18732 17052 19236 17108
rect 18732 16994 18788 17052
rect 18732 16942 18734 16994
rect 18786 16942 18788 16994
rect 18732 16930 18788 16942
rect 18508 16270 18510 16322
rect 18562 16270 18564 16322
rect 18508 16258 18564 16270
rect 19404 16212 19460 16222
rect 18620 16210 19460 16212
rect 18620 16158 19406 16210
rect 19458 16158 19460 16210
rect 18620 16156 19460 16158
rect 18396 15988 18452 15998
rect 18396 15204 18452 15932
rect 18508 15874 18564 15886
rect 18508 15822 18510 15874
rect 18562 15822 18564 15874
rect 18508 15540 18564 15822
rect 18508 15474 18564 15484
rect 18060 15092 18228 15148
rect 18396 15138 18452 15148
rect 18172 15026 18228 15036
rect 18620 14642 18676 16156
rect 19404 16146 19460 16156
rect 19516 15986 19572 17612
rect 19628 17602 19684 17612
rect 20076 17668 20132 17678
rect 20076 17574 20132 17612
rect 20300 17554 20356 18284
rect 20636 17892 20692 18396
rect 20636 17798 20692 17836
rect 21308 17780 21364 17790
rect 21308 17686 21364 17724
rect 20748 17668 20804 17678
rect 20804 17612 20916 17668
rect 20748 17574 20804 17612
rect 20300 17502 20302 17554
rect 20354 17502 20356 17554
rect 20300 17490 20356 17502
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 20636 16884 20692 16894
rect 19516 15934 19518 15986
rect 19570 15934 19572 15986
rect 19516 15922 19572 15934
rect 19740 15988 19796 15998
rect 19740 15986 20356 15988
rect 19740 15934 19742 15986
rect 19794 15934 20356 15986
rect 19740 15932 20356 15934
rect 19740 15922 19796 15932
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 20188 15540 20244 15550
rect 20188 15446 20244 15484
rect 20300 15538 20356 15932
rect 20300 15486 20302 15538
rect 20354 15486 20356 15538
rect 20300 15474 20356 15486
rect 20636 15540 20692 16828
rect 20860 16770 20916 17612
rect 21420 17554 21476 18622
rect 21868 19010 21924 19022
rect 21868 18958 21870 19010
rect 21922 18958 21924 19010
rect 21420 17502 21422 17554
rect 21474 17502 21476 17554
rect 21420 17490 21476 17502
rect 21644 17556 21700 17566
rect 21644 17462 21700 17500
rect 20860 16718 20862 16770
rect 20914 16718 20916 16770
rect 20860 16706 20916 16718
rect 21868 16660 21924 18958
rect 22204 17892 22260 17902
rect 22204 17666 22260 17836
rect 22204 17614 22206 17666
rect 22258 17614 22260 17666
rect 22204 17602 22260 17614
rect 22316 17556 22372 19966
rect 22428 19572 22484 20076
rect 22540 19908 22596 21756
rect 22652 21588 22708 21598
rect 22652 20130 22708 21532
rect 22764 21364 22820 22094
rect 23212 21924 23268 22316
rect 23324 22148 23380 22878
rect 23548 22484 23604 23100
rect 23660 22596 23716 23662
rect 23884 22708 23940 25228
rect 23996 23940 24052 26350
rect 24556 26404 24612 26414
rect 24612 26348 24836 26404
rect 24556 26310 24612 26348
rect 24220 26292 24276 26302
rect 24220 26198 24276 26236
rect 24780 25506 24836 26348
rect 24780 25454 24782 25506
rect 24834 25454 24836 25506
rect 24780 25442 24836 25454
rect 25004 26068 25060 26078
rect 25004 25506 25060 26012
rect 25116 25618 25172 26908
rect 25228 26180 25284 27020
rect 25340 26516 25396 27134
rect 25676 27746 25732 27758
rect 25676 27694 25678 27746
rect 25730 27694 25732 27746
rect 25676 27076 25732 27694
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 25676 26982 25732 27020
rect 28588 27188 28644 27198
rect 26460 26964 26516 26974
rect 26460 26870 26516 26908
rect 25340 26450 25396 26460
rect 26684 26516 26740 26526
rect 26684 26402 26740 26460
rect 26684 26350 26686 26402
rect 26738 26350 26740 26402
rect 26684 26338 26740 26350
rect 27580 26516 27636 26526
rect 27580 26290 27636 26460
rect 28588 26516 28644 27132
rect 40012 27186 40068 27198
rect 40012 27134 40014 27186
rect 40066 27134 40068 27186
rect 37660 27076 37716 27086
rect 37660 26982 37716 27020
rect 28588 26450 28644 26460
rect 39900 26852 39956 26862
rect 27804 26404 27860 26414
rect 27804 26310 27860 26348
rect 27580 26238 27582 26290
rect 27634 26238 27636 26290
rect 27580 26226 27636 26238
rect 37660 26292 37716 26302
rect 37660 26198 37716 26236
rect 25340 26180 25396 26190
rect 25228 26178 25396 26180
rect 25228 26126 25342 26178
rect 25394 26126 25396 26178
rect 25228 26124 25396 26126
rect 25116 25566 25118 25618
rect 25170 25566 25172 25618
rect 25116 25554 25172 25566
rect 25004 25454 25006 25506
rect 25058 25454 25060 25506
rect 25004 25442 25060 25454
rect 25116 25396 25172 25406
rect 24892 23940 24948 23950
rect 23996 23938 24948 23940
rect 23996 23886 24894 23938
rect 24946 23886 24948 23938
rect 23996 23884 24948 23886
rect 24892 23716 24948 23884
rect 25116 23938 25172 25340
rect 25228 25282 25284 25294
rect 25228 25230 25230 25282
rect 25282 25230 25284 25282
rect 25228 24052 25284 25230
rect 25340 24612 25396 26124
rect 39900 26178 39956 26796
rect 40012 26292 40068 27134
rect 40012 26226 40068 26236
rect 39900 26126 39902 26178
rect 39954 26126 39956 26178
rect 39900 26114 39956 26126
rect 26572 26068 26628 26078
rect 26572 25974 26628 26012
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 25452 25396 25508 25406
rect 25452 25302 25508 25340
rect 25564 24612 25620 24622
rect 25340 24610 25732 24612
rect 25340 24558 25566 24610
rect 25618 24558 25732 24610
rect 25340 24556 25732 24558
rect 25564 24546 25620 24556
rect 25228 23996 25508 24052
rect 25116 23886 25118 23938
rect 25170 23886 25172 23938
rect 25116 23874 25172 23886
rect 25228 23828 25284 23838
rect 25228 23734 25284 23772
rect 25340 23826 25396 23838
rect 25340 23774 25342 23826
rect 25394 23774 25396 23826
rect 24892 23660 25172 23716
rect 23996 23156 24052 23166
rect 23996 23062 24052 23100
rect 24444 23156 24500 23166
rect 24444 23062 24500 23100
rect 24556 23154 24612 23166
rect 24556 23102 24558 23154
rect 24610 23102 24612 23154
rect 24220 23042 24276 23054
rect 24220 22990 24222 23042
rect 24274 22990 24276 23042
rect 23996 22708 24052 22718
rect 23884 22652 23996 22708
rect 23996 22642 24052 22652
rect 24220 22596 24276 22990
rect 24220 22540 24500 22596
rect 23660 22530 23716 22540
rect 23436 22372 23492 22382
rect 23548 22372 23604 22428
rect 23660 22372 23716 22382
rect 23548 22370 23716 22372
rect 23548 22318 23662 22370
rect 23714 22318 23716 22370
rect 23548 22316 23716 22318
rect 23436 22278 23492 22316
rect 23660 22306 23716 22316
rect 23884 22372 23940 22382
rect 23884 22278 23940 22316
rect 24108 22372 24164 22382
rect 24108 22370 24276 22372
rect 24108 22318 24110 22370
rect 24162 22318 24276 22370
rect 24108 22316 24276 22318
rect 24108 22306 24164 22316
rect 23324 22082 23380 22092
rect 23772 22146 23828 22158
rect 23772 22094 23774 22146
rect 23826 22094 23828 22146
rect 23212 21868 23716 21924
rect 22764 21308 23380 21364
rect 23100 20356 23156 20366
rect 22652 20078 22654 20130
rect 22706 20078 22708 20130
rect 22652 20066 22708 20078
rect 22988 20130 23044 20142
rect 22988 20078 22990 20130
rect 23042 20078 23044 20130
rect 22876 20018 22932 20030
rect 22876 19966 22878 20018
rect 22930 19966 22932 20018
rect 22876 19908 22932 19966
rect 22988 20020 23044 20078
rect 22988 19954 23044 19964
rect 22540 19852 22932 19908
rect 22428 19506 22484 19516
rect 22988 19796 23044 19806
rect 23100 19796 23156 20300
rect 22988 19794 23156 19796
rect 22988 19742 22990 19794
rect 23042 19742 23156 19794
rect 22988 19740 23156 19742
rect 22316 17490 22372 17500
rect 21868 16594 21924 16604
rect 21980 17442 22036 17454
rect 21980 17390 21982 17442
rect 22034 17390 22036 17442
rect 21196 15540 21252 15550
rect 20636 15538 21252 15540
rect 20636 15486 20638 15538
rect 20690 15486 21198 15538
rect 21250 15486 21252 15538
rect 20636 15484 21252 15486
rect 20636 15474 20692 15484
rect 19068 15314 19124 15326
rect 19068 15262 19070 15314
rect 19122 15262 19124 15314
rect 19068 15204 19124 15262
rect 19404 15314 19460 15326
rect 19404 15262 19406 15314
rect 19458 15262 19460 15314
rect 19068 15138 19124 15148
rect 19180 15202 19236 15214
rect 19180 15150 19182 15202
rect 19234 15150 19236 15202
rect 18620 14590 18622 14642
rect 18674 14590 18676 14642
rect 18620 14578 18676 14590
rect 17836 14530 18116 14532
rect 17836 14478 17838 14530
rect 17890 14478 18116 14530
rect 17836 14476 18116 14478
rect 17836 14466 17892 14476
rect 17276 14418 17332 14430
rect 17276 14366 17278 14418
rect 17330 14366 17332 14418
rect 17052 14308 17108 14318
rect 17052 14214 17108 14252
rect 17276 13972 17332 14366
rect 17388 13972 17444 13982
rect 17276 13970 17444 13972
rect 17276 13918 17390 13970
rect 17442 13918 17444 13970
rect 17276 13916 17444 13918
rect 17388 13906 17444 13916
rect 18060 13748 18116 14476
rect 18844 13860 18900 13870
rect 19180 13860 19236 15150
rect 19404 13972 19460 15262
rect 19852 15316 19908 15326
rect 19852 15222 19908 15260
rect 20412 15314 20468 15326
rect 20412 15262 20414 15314
rect 20466 15262 20468 15314
rect 19516 15092 19572 15102
rect 19516 14998 19572 15036
rect 20412 14644 20468 15262
rect 20748 14644 20804 14654
rect 20412 14642 20804 14644
rect 20412 14590 20750 14642
rect 20802 14590 20804 14642
rect 20412 14588 20804 14590
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 19404 13906 19460 13916
rect 20188 13972 20244 13982
rect 18844 13858 19236 13860
rect 18844 13806 18846 13858
rect 18898 13806 19236 13858
rect 18844 13804 19236 13806
rect 18844 13794 18900 13804
rect 17836 13746 18116 13748
rect 17836 13694 18062 13746
rect 18114 13694 18116 13746
rect 17836 13692 18116 13694
rect 15708 8372 16436 8428
rect 16828 13636 16884 13646
rect 17500 13636 17556 13646
rect 16828 13634 17556 13636
rect 16828 13582 16830 13634
rect 16882 13582 17502 13634
rect 17554 13582 17556 13634
rect 16828 13580 17556 13582
rect 16828 8428 16884 13580
rect 17500 13570 17556 13580
rect 17164 13076 17220 13086
rect 17836 13076 17892 13692
rect 18060 13682 18116 13692
rect 20188 13186 20244 13916
rect 20188 13134 20190 13186
rect 20242 13134 20244 13186
rect 20188 13122 20244 13134
rect 17164 13074 17892 13076
rect 17164 13022 17166 13074
rect 17218 13022 17838 13074
rect 17890 13022 17892 13074
rect 17164 13020 17892 13022
rect 17164 13010 17220 13020
rect 17836 13010 17892 13020
rect 20300 12964 20356 12974
rect 20300 12870 20356 12908
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 20748 8428 20804 14588
rect 21196 14644 21252 15484
rect 21980 15540 22036 17390
rect 22876 16994 22932 17006
rect 22876 16942 22878 16994
rect 22930 16942 22932 16994
rect 22876 16098 22932 16942
rect 22876 16046 22878 16098
rect 22930 16046 22932 16098
rect 22876 15988 22932 16046
rect 21980 15474 22036 15484
rect 22428 15932 22932 15988
rect 22428 15148 22484 15932
rect 22988 15426 23044 19740
rect 23212 17666 23268 17678
rect 23212 17614 23214 17666
rect 23266 17614 23268 17666
rect 23212 16994 23268 17614
rect 23212 16942 23214 16994
rect 23266 16942 23268 16994
rect 23212 16884 23268 16942
rect 23212 16818 23268 16828
rect 23324 16882 23380 21308
rect 23548 20132 23604 20142
rect 23548 18676 23604 20076
rect 23660 19796 23716 21868
rect 23772 21586 23828 22094
rect 24220 21812 24276 22316
rect 24332 22370 24388 22382
rect 24332 22318 24334 22370
rect 24386 22318 24388 22370
rect 24332 22260 24388 22318
rect 24444 22372 24500 22540
rect 24444 22306 24500 22316
rect 24332 22194 24388 22204
rect 24556 22036 24612 23102
rect 24892 22596 24948 22606
rect 24668 22484 24724 22494
rect 24724 22428 24836 22484
rect 24668 22418 24724 22428
rect 24780 22370 24836 22428
rect 24780 22318 24782 22370
rect 24834 22318 24836 22370
rect 24780 22306 24836 22318
rect 24892 22372 24948 22540
rect 24892 22370 25060 22372
rect 24892 22318 24894 22370
rect 24946 22318 25060 22370
rect 24892 22316 25060 22318
rect 24892 22306 24948 22316
rect 24668 22260 24724 22270
rect 24668 22146 24724 22204
rect 24668 22094 24670 22146
rect 24722 22094 24724 22146
rect 24668 22082 24724 22094
rect 24556 21970 24612 21980
rect 24220 21746 24276 21756
rect 23772 21534 23774 21586
rect 23826 21534 23828 21586
rect 23772 21522 23828 21534
rect 24332 21700 24388 21710
rect 24332 21586 24388 21644
rect 25004 21700 25060 22316
rect 25116 22260 25172 23660
rect 25340 23268 25396 23774
rect 25452 23380 25508 23996
rect 25676 23938 25732 24556
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 25676 23886 25678 23938
rect 25730 23886 25732 23938
rect 25452 23324 25620 23380
rect 25228 23212 25396 23268
rect 25228 22484 25284 23212
rect 25340 23044 25396 23054
rect 25340 23042 25508 23044
rect 25340 22990 25342 23042
rect 25394 22990 25508 23042
rect 25340 22988 25508 22990
rect 25340 22978 25396 22988
rect 25228 22418 25284 22428
rect 25452 22930 25508 22988
rect 25452 22878 25454 22930
rect 25506 22878 25508 22930
rect 25340 22260 25396 22270
rect 25116 22258 25396 22260
rect 25116 22206 25342 22258
rect 25394 22206 25396 22258
rect 25116 22204 25396 22206
rect 25340 22194 25396 22204
rect 25228 21700 25284 21710
rect 25004 21698 25284 21700
rect 25004 21646 25230 21698
rect 25282 21646 25284 21698
rect 25004 21644 25284 21646
rect 24332 21534 24334 21586
rect 24386 21534 24388 21586
rect 24220 21476 24276 21486
rect 23996 21364 24052 21402
rect 23996 21140 24052 21308
rect 23772 21084 24052 21140
rect 23772 20130 23828 21084
rect 23772 20078 23774 20130
rect 23826 20078 23828 20130
rect 23772 20066 23828 20078
rect 23996 20804 24052 20814
rect 23996 20132 24052 20748
rect 23996 20130 24164 20132
rect 23996 20078 23998 20130
rect 24050 20078 24164 20130
rect 23996 20076 24164 20078
rect 23996 20066 24052 20076
rect 23660 19740 24052 19796
rect 23996 19236 24052 19740
rect 23996 19142 24052 19180
rect 23548 18610 23604 18620
rect 23996 18564 24052 18574
rect 24108 18564 24164 20076
rect 24220 20018 24276 21420
rect 24220 19966 24222 20018
rect 24274 19966 24276 20018
rect 24220 19954 24276 19966
rect 24332 19572 24388 21534
rect 24556 21586 24612 21598
rect 24556 21534 24558 21586
rect 24610 21534 24612 21586
rect 24444 21474 24500 21486
rect 24444 21422 24446 21474
rect 24498 21422 24500 21474
rect 24444 20132 24500 21422
rect 24556 20244 24612 21534
rect 24556 20178 24612 20188
rect 24444 20066 24500 20076
rect 24668 20018 24724 20030
rect 24668 19966 24670 20018
rect 24722 19966 24724 20018
rect 24444 19906 24500 19918
rect 24444 19854 24446 19906
rect 24498 19854 24500 19906
rect 24444 19796 24500 19854
rect 24556 19908 24612 19918
rect 24556 19814 24612 19852
rect 24444 19730 24500 19740
rect 24332 19516 24612 19572
rect 24444 19236 24500 19274
rect 24444 19170 24500 19180
rect 24556 19234 24612 19516
rect 24668 19460 24724 19966
rect 24668 19404 24836 19460
rect 24556 19182 24558 19234
rect 24610 19182 24612 19234
rect 24556 19170 24612 19182
rect 24220 19012 24276 19022
rect 24220 18918 24276 18956
rect 24332 19010 24388 19022
rect 24332 18958 24334 19010
rect 24386 18958 24388 19010
rect 23996 18562 24164 18564
rect 23996 18510 23998 18562
rect 24050 18510 24164 18562
rect 23996 18508 24164 18510
rect 24220 18564 24276 18574
rect 24332 18564 24388 18958
rect 24220 18562 24388 18564
rect 24220 18510 24222 18562
rect 24274 18510 24388 18562
rect 24220 18508 24388 18510
rect 24444 18676 24500 18686
rect 23996 18498 24052 18508
rect 24220 18498 24276 18508
rect 23324 16830 23326 16882
rect 23378 16830 23380 16882
rect 23324 16818 23380 16830
rect 23660 18450 23716 18462
rect 23660 18398 23662 18450
rect 23714 18398 23716 18450
rect 23548 16772 23604 16782
rect 23548 16678 23604 16716
rect 22988 15374 22990 15426
rect 23042 15374 23044 15426
rect 22988 15362 23044 15374
rect 23100 16660 23156 16670
rect 23660 16660 23716 18398
rect 23772 18340 23828 18350
rect 24444 18340 24500 18620
rect 24780 18452 24836 19404
rect 25004 19236 25060 21644
rect 25228 21634 25284 21644
rect 25340 21476 25396 21486
rect 25340 21382 25396 21420
rect 25452 20692 25508 22878
rect 25564 22596 25620 23324
rect 25676 22932 25732 23886
rect 28588 24052 28644 24062
rect 26460 23828 26516 23838
rect 26460 23734 26516 23772
rect 25900 23154 25956 23166
rect 25900 23102 25902 23154
rect 25954 23102 25956 23154
rect 25900 22932 25956 23102
rect 26684 23044 26740 23054
rect 25676 22930 25956 22932
rect 25676 22878 25678 22930
rect 25730 22878 25956 22930
rect 25676 22876 25956 22878
rect 26012 23042 26740 23044
rect 26012 22990 26686 23042
rect 26738 22990 26740 23042
rect 26012 22988 26740 22990
rect 25676 22866 25732 22876
rect 26012 22596 26068 22988
rect 26684 22978 26740 22988
rect 25564 22540 25732 22596
rect 25564 22372 25620 22382
rect 25564 22278 25620 22316
rect 25564 22148 25620 22158
rect 25564 21698 25620 22092
rect 25676 22036 25732 22540
rect 25788 22540 26068 22596
rect 25788 22482 25844 22540
rect 25788 22430 25790 22482
rect 25842 22430 25844 22482
rect 25788 22418 25844 22430
rect 26124 22484 26180 22494
rect 26348 22484 26404 22494
rect 26180 22482 26404 22484
rect 26180 22430 26350 22482
rect 26402 22430 26404 22482
rect 26180 22428 26404 22430
rect 26124 22418 26180 22428
rect 26348 22418 26404 22428
rect 26572 22372 26628 22382
rect 26572 22278 26628 22316
rect 26684 22370 26740 22382
rect 26684 22318 26686 22370
rect 26738 22318 26740 22370
rect 25900 22260 25956 22270
rect 25900 22166 25956 22204
rect 26236 22260 26292 22270
rect 26236 22258 26516 22260
rect 26236 22206 26238 22258
rect 26290 22206 26516 22258
rect 26236 22204 26516 22206
rect 26236 22194 26292 22204
rect 25676 21980 26068 22036
rect 26012 21810 26068 21980
rect 26012 21758 26014 21810
rect 26066 21758 26068 21810
rect 26012 21746 26068 21758
rect 25564 21646 25566 21698
rect 25618 21646 25620 21698
rect 25564 21634 25620 21646
rect 26236 21698 26292 21710
rect 26236 21646 26238 21698
rect 26290 21646 26292 21698
rect 25788 21588 25844 21598
rect 26236 21588 26292 21646
rect 25788 21586 26292 21588
rect 25788 21534 25790 21586
rect 25842 21534 26292 21586
rect 25788 21532 26292 21534
rect 26348 21588 26404 21598
rect 25788 20804 25844 21532
rect 26348 21494 26404 21532
rect 26460 21364 26516 22204
rect 26684 22036 26740 22318
rect 28588 22372 28644 23996
rect 40012 24050 40068 24062
rect 40012 23998 40014 24050
rect 40066 23998 40068 24050
rect 37660 23940 37716 23950
rect 37660 23846 37716 23884
rect 40012 23604 40068 23998
rect 40012 23538 40068 23548
rect 28812 23156 28868 23166
rect 28812 23042 28868 23100
rect 37660 23156 37716 23166
rect 37660 23062 37716 23100
rect 28812 22990 28814 23042
rect 28866 22990 28868 23042
rect 28812 22978 28868 22990
rect 40012 22932 40068 22942
rect 40012 22838 40068 22876
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 28588 22306 28644 22316
rect 26684 21970 26740 21980
rect 25788 20738 25844 20748
rect 26348 21308 26516 21364
rect 28588 21588 28644 21598
rect 25676 20692 25732 20702
rect 25452 20690 25732 20692
rect 25452 20638 25678 20690
rect 25730 20638 25732 20690
rect 25452 20636 25732 20638
rect 25676 20018 25732 20636
rect 25676 19966 25678 20018
rect 25730 19966 25732 20018
rect 25004 19170 25060 19180
rect 25340 19906 25396 19918
rect 25340 19854 25342 19906
rect 25394 19854 25396 19906
rect 24780 18386 24836 18396
rect 25340 19012 25396 19854
rect 25676 19234 25732 19966
rect 26348 19796 26404 21308
rect 26460 20132 26516 20142
rect 26460 20038 26516 20076
rect 26348 19730 26404 19740
rect 26460 19908 26516 19918
rect 26460 19346 26516 19852
rect 28588 19906 28644 21532
rect 37660 21588 37716 21598
rect 37660 21494 37716 21532
rect 40012 21362 40068 21374
rect 40012 21310 40014 21362
rect 40066 21310 40068 21362
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 40012 20916 40068 21310
rect 40012 20850 40068 20860
rect 28588 19854 28590 19906
rect 28642 19854 28644 19906
rect 28588 19842 28644 19854
rect 37660 20018 37716 20030
rect 37660 19966 37662 20018
rect 37714 19966 37716 20018
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 26460 19294 26462 19346
rect 26514 19294 26516 19346
rect 26460 19282 26516 19294
rect 28028 19348 28084 19358
rect 25676 19182 25678 19234
rect 25730 19182 25732 19234
rect 25676 19012 25732 19182
rect 25340 19010 25732 19012
rect 25340 18958 25342 19010
rect 25394 18958 25732 19010
rect 25340 18956 25732 18958
rect 26124 19012 26180 19022
rect 23772 18338 23940 18340
rect 23772 18286 23774 18338
rect 23826 18286 23940 18338
rect 23772 18284 23940 18286
rect 23772 18274 23828 18284
rect 23884 17780 23940 18284
rect 24220 18284 24500 18340
rect 23996 17780 24052 17790
rect 23884 17778 24052 17780
rect 23884 17726 23998 17778
rect 24050 17726 24052 17778
rect 23884 17724 24052 17726
rect 23996 17714 24052 17724
rect 24220 16770 24276 18284
rect 24444 16996 24500 17006
rect 24444 16902 24500 16940
rect 25340 16884 25396 18956
rect 26124 17780 26180 18956
rect 27916 18452 27972 18462
rect 27916 18358 27972 18396
rect 28028 18450 28084 19292
rect 28588 19348 28644 19358
rect 28588 19254 28644 19292
rect 37660 19348 37716 19966
rect 40012 19794 40068 19806
rect 40012 19742 40014 19794
rect 40066 19742 40068 19794
rect 40012 19572 40068 19742
rect 40012 19506 40068 19516
rect 37660 19282 37716 19292
rect 28028 18398 28030 18450
rect 28082 18398 28084 18450
rect 28028 18386 28084 18398
rect 37660 18450 37716 18462
rect 37660 18398 37662 18450
rect 37714 18398 37716 18450
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 26124 17686 26180 17724
rect 37660 17780 37716 18398
rect 40012 18228 40068 18238
rect 40012 18134 40068 18172
rect 37660 17714 37716 17724
rect 26572 17442 26628 17454
rect 26572 17390 26574 17442
rect 26626 17390 26628 17442
rect 24220 16718 24222 16770
rect 24274 16718 24276 16770
rect 24220 16706 24276 16718
rect 24332 16772 24388 16782
rect 24332 16678 24388 16716
rect 23772 16660 23828 16670
rect 23660 16604 23772 16660
rect 22316 15092 22484 15148
rect 22540 15314 22596 15326
rect 22540 15262 22542 15314
rect 22594 15262 22596 15314
rect 21196 14578 21252 14588
rect 22092 14644 22148 14654
rect 22092 14550 22148 14588
rect 21868 13748 21924 13758
rect 22316 13748 22372 15092
rect 22540 14754 22596 15262
rect 23100 15316 23156 16604
rect 23772 16566 23828 16604
rect 23884 16658 23940 16670
rect 23884 16606 23886 16658
rect 23938 16606 23940 16658
rect 23884 16324 23940 16606
rect 23660 16268 23940 16324
rect 23660 16210 23716 16268
rect 23660 16158 23662 16210
rect 23714 16158 23716 16210
rect 23660 16146 23716 16158
rect 23100 15222 23156 15260
rect 22764 15202 22820 15214
rect 22764 15150 22766 15202
rect 22818 15150 22820 15202
rect 22764 15148 22820 15150
rect 22540 14702 22542 14754
rect 22594 14702 22596 14754
rect 22540 14690 22596 14702
rect 22652 15092 22820 15148
rect 22428 14644 22484 14654
rect 22428 14530 22484 14588
rect 22428 14478 22430 14530
rect 22482 14478 22484 14530
rect 22428 14466 22484 14478
rect 22540 14308 22596 14318
rect 22540 14214 22596 14252
rect 22540 13860 22596 13870
rect 22652 13860 22708 15092
rect 22540 13858 22708 13860
rect 22540 13806 22542 13858
rect 22594 13806 22708 13858
rect 22540 13804 22708 13806
rect 23996 14530 24052 14542
rect 23996 14478 23998 14530
rect 24050 14478 24052 14530
rect 23996 14308 24052 14478
rect 22540 13794 22596 13804
rect 21868 13746 22372 13748
rect 21868 13694 21870 13746
rect 21922 13694 22372 13746
rect 21868 13692 22372 13694
rect 21868 13682 21924 13692
rect 20972 13636 21028 13646
rect 20972 13634 21140 13636
rect 20972 13582 20974 13634
rect 21026 13582 21140 13634
rect 20972 13580 21140 13582
rect 20972 13570 21028 13580
rect 16828 8372 17108 8428
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 15484 5236 15540 5246
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 15484 800 15540 5180
rect 15708 5122 15764 8372
rect 16716 5236 16772 5246
rect 16716 5142 16772 5180
rect 15708 5070 15710 5122
rect 15762 5070 15764 5122
rect 15708 5058 15764 5070
rect 17052 3554 17108 8372
rect 20412 8372 20804 8428
rect 21084 12964 21140 13580
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 20412 4338 20468 8372
rect 20412 4286 20414 4338
rect 20466 4286 20468 4338
rect 20412 4274 20468 4286
rect 17052 3502 17054 3554
rect 17106 3502 17108 3554
rect 17052 3490 17108 3502
rect 20188 4116 20244 4126
rect 16828 3444 16884 3454
rect 16828 800 16884 3388
rect 18060 3444 18116 3454
rect 18060 3330 18116 3388
rect 18060 3278 18062 3330
rect 18114 3278 18116 3330
rect 18060 3266 18116 3278
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 20188 800 20244 4060
rect 20860 3668 20916 3678
rect 20860 800 20916 3612
rect 21084 3554 21140 12908
rect 23884 12738 23940 12750
rect 23884 12686 23886 12738
rect 23938 12686 23940 12738
rect 23884 8428 23940 12686
rect 23996 12740 24052 14252
rect 24220 14308 24276 14318
rect 24220 14214 24276 14252
rect 25340 13970 25396 16828
rect 25788 16996 25844 17006
rect 25788 16212 25844 16940
rect 25788 16118 25844 16156
rect 26236 16884 26292 16894
rect 26572 16884 26628 17390
rect 26292 16828 26628 16884
rect 26236 16210 26292 16828
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 26236 16158 26238 16210
rect 26290 16158 26292 16210
rect 26236 16146 26292 16158
rect 28588 16212 28644 16222
rect 25340 13918 25342 13970
rect 25394 13918 25396 13970
rect 25340 13906 25396 13918
rect 25452 14308 25508 14318
rect 24668 13634 24724 13646
rect 24668 13582 24670 13634
rect 24722 13582 24724 13634
rect 24220 12740 24276 12750
rect 24668 12740 24724 13582
rect 23996 12738 24724 12740
rect 23996 12686 24222 12738
rect 24274 12686 24724 12738
rect 23996 12684 24724 12686
rect 23772 8372 23940 8428
rect 24220 8428 24276 12684
rect 24220 8372 24612 8428
rect 23548 5236 23604 5246
rect 21420 4116 21476 4126
rect 21420 4022 21476 4060
rect 22092 3668 22148 3678
rect 22092 3574 22148 3612
rect 21084 3502 21086 3554
rect 21138 3502 21140 3554
rect 21084 3490 21140 3502
rect 22876 3444 22932 3454
rect 22876 800 22932 3388
rect 23548 800 23604 5180
rect 23772 5122 23828 8372
rect 23772 5070 23774 5122
rect 23826 5070 23828 5122
rect 23772 5058 23828 5070
rect 24220 4116 24276 4126
rect 24220 800 24276 4060
rect 24556 3554 24612 8372
rect 24780 5236 24836 5246
rect 24780 5142 24836 5180
rect 25452 4338 25508 14252
rect 25452 4286 25454 4338
rect 25506 4286 25508 4338
rect 25452 4274 25508 4286
rect 26236 4116 26292 4126
rect 26236 4022 26292 4060
rect 24556 3502 24558 3554
rect 24610 3502 24612 3554
rect 24556 3490 24612 3502
rect 24892 3668 24948 3678
rect 24892 800 24948 3612
rect 25564 3666 25620 3678
rect 25564 3614 25566 3666
rect 25618 3614 25620 3666
rect 25564 3444 25620 3614
rect 28588 3554 28644 16156
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 40236 12290 40292 12302
rect 40236 12238 40238 12290
rect 40290 12238 40292 12290
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 40236 11508 40292 12238
rect 40236 11442 40292 11452
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 29372 3668 29428 3678
rect 29372 3574 29428 3612
rect 28588 3502 28590 3554
rect 28642 3502 28644 3554
rect 28588 3490 28644 3502
rect 25564 3378 25620 3388
rect 15456 0 15568 800
rect 16800 0 16912 800
rect 20160 0 20272 800
rect 20832 0 20944 800
rect 22848 0 22960 800
rect 23520 0 23632 800
rect 24192 0 24304 800
rect 24864 0 24976 800
<< via2 >>
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 20860 38220 20916 38276
rect 22092 38274 22148 38276
rect 22092 38222 22094 38274
rect 22094 38222 22146 38274
rect 22146 38222 22148 38274
rect 22092 38220 22148 38222
rect 24892 38220 24948 38276
rect 26124 38274 26180 38276
rect 26124 38222 26126 38274
rect 26126 38222 26178 38274
rect 26178 38222 26180 38274
rect 26124 38220 26180 38222
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 19516 37436 19572 37492
rect 20748 37490 20804 37492
rect 20748 37438 20750 37490
rect 20750 37438 20802 37490
rect 20802 37438 20804 37490
rect 20748 37436 20804 37438
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 17052 28588 17108 28644
rect 4172 27580 4228 27636
rect 1932 26236 1988 26292
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 4284 27074 4340 27076
rect 4284 27022 4286 27074
rect 4286 27022 4338 27074
rect 4338 27022 4340 27074
rect 4284 27020 4340 27022
rect 12684 27020 12740 27076
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 20076 28642 20132 28644
rect 20076 28590 20078 28642
rect 20078 28590 20130 28642
rect 20130 28590 20132 28642
rect 20076 28588 20132 28590
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 18396 27746 18452 27748
rect 18396 27694 18398 27746
rect 18398 27694 18450 27746
rect 18450 27694 18452 27746
rect 18396 27692 18452 27694
rect 20748 27692 20804 27748
rect 14700 26572 14756 26628
rect 14588 26460 14644 26516
rect 12684 26348 12740 26404
rect 13692 26236 13748 26292
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 14924 25676 14980 25732
rect 15260 26572 15316 26628
rect 13916 24444 13972 24500
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 10780 22540 10836 22596
rect 10108 22370 10164 22372
rect 10108 22318 10110 22370
rect 10110 22318 10162 22370
rect 10162 22318 10164 22370
rect 10108 22316 10164 22318
rect 11676 23042 11732 23044
rect 11676 22990 11678 23042
rect 11678 22990 11730 23042
rect 11730 22990 11732 23042
rect 11676 22988 11732 22990
rect 13580 22988 13636 23044
rect 10892 22316 10948 22372
rect 12908 21644 12964 21700
rect 13132 22316 13188 22372
rect 13804 23042 13860 23044
rect 13804 22990 13806 23042
rect 13806 22990 13858 23042
rect 13858 22990 13860 23042
rect 13804 22988 13860 22990
rect 17724 27074 17780 27076
rect 17724 27022 17726 27074
rect 17726 27022 17778 27074
rect 17778 27022 17780 27074
rect 17724 27020 17780 27022
rect 15820 26850 15876 26852
rect 15820 26798 15822 26850
rect 15822 26798 15874 26850
rect 15874 26798 15876 26850
rect 15820 26796 15876 26798
rect 17052 26796 17108 26852
rect 15932 26514 15988 26516
rect 15932 26462 15934 26514
rect 15934 26462 15986 26514
rect 15986 26462 15988 26514
rect 15932 26460 15988 26462
rect 16156 26402 16212 26404
rect 16156 26350 16158 26402
rect 16158 26350 16210 26402
rect 16210 26350 16212 26402
rect 16156 26348 16212 26350
rect 15484 26290 15540 26292
rect 15484 26238 15486 26290
rect 15486 26238 15538 26290
rect 15538 26238 15540 26290
rect 15484 26236 15540 26238
rect 16492 25452 16548 25508
rect 16156 24668 16212 24724
rect 15260 24498 15316 24500
rect 15260 24446 15262 24498
rect 15262 24446 15314 24498
rect 15314 24446 15316 24498
rect 15260 24444 15316 24446
rect 14364 23548 14420 23604
rect 15372 23772 15428 23828
rect 14476 23042 14532 23044
rect 14476 22990 14478 23042
rect 14478 22990 14530 23042
rect 14530 22990 14532 23042
rect 14476 22988 14532 22990
rect 14364 22370 14420 22372
rect 14364 22318 14366 22370
rect 14366 22318 14418 22370
rect 14418 22318 14420 22370
rect 14364 22316 14420 22318
rect 14812 22316 14868 22372
rect 14252 22204 14308 22260
rect 4172 21420 4228 21476
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 1932 20188 1988 20244
rect 1932 19794 1988 19796
rect 1932 19742 1934 19794
rect 1934 19742 1986 19794
rect 1986 19742 1988 19794
rect 1932 19740 1988 19742
rect 14700 22204 14756 22260
rect 14364 21644 14420 21700
rect 15148 21810 15204 21812
rect 15148 21758 15150 21810
rect 15150 21758 15202 21810
rect 15202 21758 15204 21810
rect 15148 21756 15204 21758
rect 14812 21698 14868 21700
rect 14812 21646 14814 21698
rect 14814 21646 14866 21698
rect 14866 21646 14868 21698
rect 14812 21644 14868 21646
rect 4284 20018 4340 20020
rect 4284 19966 4286 20018
rect 4286 19966 4338 20018
rect 4338 19966 4340 20018
rect 4284 19964 4340 19966
rect 12460 19964 12516 20020
rect 11788 19906 11844 19908
rect 11788 19854 11790 19906
rect 11790 19854 11842 19906
rect 11842 19854 11844 19906
rect 11788 19852 11844 19854
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 4172 19292 4228 19348
rect 9884 19346 9940 19348
rect 9884 19294 9886 19346
rect 9886 19294 9938 19346
rect 9938 19294 9940 19346
rect 9884 19292 9940 19294
rect 4284 19234 4340 19236
rect 4284 19182 4286 19234
rect 4286 19182 4338 19234
rect 4338 19182 4340 19234
rect 4284 19180 4340 19182
rect 1932 18844 1988 18900
rect 12684 19292 12740 19348
rect 4284 18450 4340 18452
rect 4284 18398 4286 18450
rect 4286 18398 4338 18450
rect 4338 18398 4340 18450
rect 4284 18396 4340 18398
rect 14364 20130 14420 20132
rect 14364 20078 14366 20130
rect 14366 20078 14418 20130
rect 14418 20078 14420 20130
rect 14364 20076 14420 20078
rect 13692 19292 13748 19348
rect 13468 19180 13524 19236
rect 14364 19906 14420 19908
rect 14364 19854 14366 19906
rect 14366 19854 14418 19906
rect 14418 19854 14420 19906
rect 14364 19852 14420 19854
rect 15036 19516 15092 19572
rect 15148 19852 15204 19908
rect 14140 19292 14196 19348
rect 13916 18956 13972 19012
rect 12908 18396 12964 18452
rect 14028 18396 14084 18452
rect 13692 18338 13748 18340
rect 13692 18286 13694 18338
rect 13694 18286 13746 18338
rect 13746 18286 13748 18338
rect 13692 18284 13748 18286
rect 1932 18226 1988 18228
rect 1932 18174 1934 18226
rect 1934 18174 1986 18226
rect 1986 18174 1988 18226
rect 1932 18172 1988 18174
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 4284 17666 4340 17668
rect 4284 17614 4286 17666
rect 4286 17614 4338 17666
rect 4338 17614 4340 17666
rect 4284 17612 4340 17614
rect 11116 17612 11172 17668
rect 1932 16828 1988 16884
rect 11116 17052 11172 17108
rect 13244 17388 13300 17444
rect 14924 19010 14980 19012
rect 14924 18958 14926 19010
rect 14926 18958 14978 19010
rect 14978 18958 14980 19010
rect 14924 18956 14980 18958
rect 15372 23548 15428 23604
rect 16156 23548 16212 23604
rect 15596 22988 15652 23044
rect 15932 22316 15988 22372
rect 16268 22988 16324 23044
rect 18844 26572 18900 26628
rect 19068 26290 19124 26292
rect 19068 26238 19070 26290
rect 19070 26238 19122 26290
rect 19122 26238 19124 26290
rect 19068 26236 19124 26238
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20188 26684 20244 26740
rect 20300 26908 20356 26964
rect 20044 26628 20100 26630
rect 20860 27132 20916 27188
rect 21980 27132 22036 27188
rect 20412 26796 20468 26852
rect 19740 26290 19796 26292
rect 19740 26238 19742 26290
rect 19742 26238 19794 26290
rect 19794 26238 19796 26290
rect 19740 26236 19796 26238
rect 17500 25676 17556 25732
rect 16716 23772 16772 23828
rect 16604 23378 16660 23380
rect 16604 23326 16606 23378
rect 16606 23326 16658 23378
rect 16658 23326 16660 23378
rect 16604 23324 16660 23326
rect 16380 22316 16436 22372
rect 15820 21698 15876 21700
rect 15820 21646 15822 21698
rect 15822 21646 15874 21698
rect 15874 21646 15876 21698
rect 15820 21644 15876 21646
rect 15484 20130 15540 20132
rect 15484 20078 15486 20130
rect 15486 20078 15538 20130
rect 15538 20078 15540 20130
rect 15484 20076 15540 20078
rect 14364 17442 14420 17444
rect 14364 17390 14366 17442
rect 14366 17390 14418 17442
rect 14418 17390 14420 17442
rect 14364 17388 14420 17390
rect 14588 17106 14644 17108
rect 14588 17054 14590 17106
rect 14590 17054 14642 17106
rect 14642 17054 14644 17106
rect 14588 17052 14644 17054
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 14924 16882 14980 16884
rect 14924 16830 14926 16882
rect 14926 16830 14978 16882
rect 14978 16830 14980 16882
rect 14924 16828 14980 16830
rect 14364 16716 14420 16772
rect 15596 17836 15652 17892
rect 16492 22092 16548 22148
rect 16828 21868 16884 21924
rect 16940 21756 16996 21812
rect 16268 20130 16324 20132
rect 16268 20078 16270 20130
rect 16270 20078 16322 20130
rect 16322 20078 16324 20130
rect 16268 20076 16324 20078
rect 16604 20018 16660 20020
rect 16604 19966 16606 20018
rect 16606 19966 16658 20018
rect 16658 19966 16660 20018
rect 16604 19964 16660 19966
rect 16828 19852 16884 19908
rect 17276 25506 17332 25508
rect 17276 25454 17278 25506
rect 17278 25454 17330 25506
rect 17330 25454 17332 25506
rect 17276 25452 17332 25454
rect 17388 25116 17444 25172
rect 18172 25452 18228 25508
rect 17612 24722 17668 24724
rect 17612 24670 17614 24722
rect 17614 24670 17666 24722
rect 17666 24670 17668 24722
rect 17612 24668 17668 24670
rect 17948 23996 18004 24052
rect 19292 25506 19348 25508
rect 19292 25454 19294 25506
rect 19294 25454 19346 25506
rect 19346 25454 19348 25506
rect 19292 25452 19348 25454
rect 18844 25116 18900 25172
rect 17388 22370 17444 22372
rect 17388 22318 17390 22370
rect 17390 22318 17442 22370
rect 17442 22318 17444 22370
rect 17388 22316 17444 22318
rect 17500 22146 17556 22148
rect 17500 22094 17502 22146
rect 17502 22094 17554 22146
rect 17554 22094 17556 22146
rect 17500 22092 17556 22094
rect 17500 20802 17556 20804
rect 17500 20750 17502 20802
rect 17502 20750 17554 20802
rect 17554 20750 17556 20802
rect 17500 20748 17556 20750
rect 18172 23436 18228 23492
rect 17724 23324 17780 23380
rect 18396 23324 18452 23380
rect 18060 22930 18116 22932
rect 18060 22878 18062 22930
rect 18062 22878 18114 22930
rect 18114 22878 18116 22930
rect 18060 22876 18116 22878
rect 17724 22652 17780 22708
rect 17724 21868 17780 21924
rect 17836 21420 17892 21476
rect 18396 22652 18452 22708
rect 19180 24946 19236 24948
rect 19180 24894 19182 24946
rect 19182 24894 19234 24946
rect 19234 24894 19236 24946
rect 19180 24892 19236 24894
rect 18956 24050 19012 24052
rect 18956 23998 18958 24050
rect 18958 23998 19010 24050
rect 19010 23998 19012 24050
rect 18956 23996 19012 23998
rect 18844 22540 18900 22596
rect 18732 22428 18788 22484
rect 18620 22316 18676 22372
rect 18508 22258 18564 22260
rect 18508 22206 18510 22258
rect 18510 22206 18562 22258
rect 18562 22206 18564 22258
rect 18508 22204 18564 22206
rect 19628 25394 19684 25396
rect 19628 25342 19630 25394
rect 19630 25342 19682 25394
rect 19682 25342 19684 25394
rect 19628 25340 19684 25342
rect 20188 26290 20244 26292
rect 20188 26238 20190 26290
rect 20190 26238 20242 26290
rect 20242 26238 20244 26290
rect 20188 26236 20244 26238
rect 19964 25506 20020 25508
rect 19964 25454 19966 25506
rect 19966 25454 20018 25506
rect 20018 25454 20020 25506
rect 19964 25452 20020 25454
rect 19852 25228 19908 25284
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 21308 26962 21364 26964
rect 21308 26910 21310 26962
rect 21310 26910 21362 26962
rect 21362 26910 21364 26962
rect 21308 26908 21364 26910
rect 21756 27074 21812 27076
rect 21756 27022 21758 27074
rect 21758 27022 21810 27074
rect 21810 27022 21812 27074
rect 21756 27020 21812 27022
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 22428 27074 22484 27076
rect 22428 27022 22430 27074
rect 22430 27022 22482 27074
rect 22482 27022 22484 27074
rect 22428 27020 22484 27022
rect 25228 27020 25284 27076
rect 21980 26908 22036 26964
rect 21644 26796 21700 26852
rect 20860 26684 20916 26740
rect 23996 26908 24052 26964
rect 20748 26402 20804 26404
rect 20748 26350 20750 26402
rect 20750 26350 20802 26402
rect 20802 26350 20804 26402
rect 20748 26348 20804 26350
rect 25116 26908 25172 26964
rect 24444 26514 24500 26516
rect 24444 26462 24446 26514
rect 24446 26462 24498 26514
rect 24498 26462 24500 26514
rect 24444 26460 24500 26462
rect 20972 26290 21028 26292
rect 20972 26238 20974 26290
rect 20974 26238 21026 26290
rect 21026 26238 21028 26290
rect 20972 26236 21028 26238
rect 20412 25340 20468 25396
rect 20972 25676 21028 25732
rect 20300 24892 20356 24948
rect 20860 24892 20916 24948
rect 19852 24444 19908 24500
rect 19180 23324 19236 23380
rect 19404 23266 19460 23268
rect 19404 23214 19406 23266
rect 19406 23214 19458 23266
rect 19458 23214 19460 23266
rect 19404 23212 19460 23214
rect 18732 22092 18788 22148
rect 17500 20076 17556 20132
rect 16604 18450 16660 18452
rect 16604 18398 16606 18450
rect 16606 18398 16658 18450
rect 16658 18398 16660 18450
rect 16604 18396 16660 18398
rect 17500 18450 17556 18452
rect 17500 18398 17502 18450
rect 17502 18398 17554 18450
rect 17554 18398 17556 18450
rect 17500 18396 17556 18398
rect 16380 18172 16436 18228
rect 16268 17836 16324 17892
rect 15148 16828 15204 16884
rect 15036 16716 15092 16772
rect 15148 15314 15204 15316
rect 15148 15262 15150 15314
rect 15150 15262 15202 15314
rect 15202 15262 15204 15314
rect 15148 15260 15204 15262
rect 14364 15202 14420 15204
rect 14364 15150 14366 15202
rect 14366 15150 14418 15202
rect 14418 15150 14420 15202
rect 14364 15148 14420 15150
rect 15260 15202 15316 15204
rect 15260 15150 15262 15202
rect 15262 15150 15314 15202
rect 15314 15150 15316 15202
rect 15260 15148 15316 15150
rect 17388 15932 17444 15988
rect 17724 19852 17780 19908
rect 16380 15484 16436 15540
rect 16044 15260 16100 15316
rect 16828 15260 16884 15316
rect 15596 15148 15652 15204
rect 14700 14252 14756 14308
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 17500 15148 17556 15204
rect 17052 15036 17108 15092
rect 22652 25676 22708 25732
rect 23100 26290 23156 26292
rect 23100 26238 23102 26290
rect 23102 26238 23154 26290
rect 23154 26238 23156 26290
rect 23100 26236 23156 26238
rect 23660 25676 23716 25732
rect 22540 25340 22596 25396
rect 21196 25228 21252 25284
rect 21980 25282 22036 25284
rect 21980 25230 21982 25282
rect 21982 25230 22034 25282
rect 22034 25230 22036 25282
rect 21980 25228 22036 25230
rect 23772 25340 23828 25396
rect 22988 25282 23044 25284
rect 22988 25230 22990 25282
rect 22990 25230 23042 25282
rect 23042 25230 23044 25282
rect 22988 25228 23044 25230
rect 19836 23546 19892 23548
rect 19516 22652 19572 22708
rect 19628 23436 19684 23492
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 20188 23324 20244 23380
rect 19516 22370 19572 22372
rect 19516 22318 19518 22370
rect 19518 22318 19570 22370
rect 19570 22318 19572 22370
rect 19516 22316 19572 22318
rect 20636 24498 20692 24500
rect 20636 24446 20638 24498
rect 20638 24446 20690 24498
rect 20690 24446 20692 24498
rect 20636 24444 20692 24446
rect 20300 23212 20356 23268
rect 20300 22540 20356 22596
rect 20412 22092 20468 22148
rect 19628 21868 19684 21924
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 19628 20802 19684 20804
rect 19628 20750 19630 20802
rect 19630 20750 19682 20802
rect 19682 20750 19684 20802
rect 19628 20748 19684 20750
rect 19404 20524 19460 20580
rect 18732 19964 18788 20020
rect 18508 18396 18564 18452
rect 20300 21756 20356 21812
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 19852 20188 19908 20244
rect 20636 23826 20692 23828
rect 20636 23774 20638 23826
rect 20638 23774 20690 23826
rect 20690 23774 20692 23826
rect 20636 23772 20692 23774
rect 21308 23266 21364 23268
rect 21308 23214 21310 23266
rect 21310 23214 21362 23266
rect 21362 23214 21364 23266
rect 21308 23212 21364 23214
rect 21532 22876 21588 22932
rect 21420 22316 21476 22372
rect 21644 22316 21700 22372
rect 20860 21980 20916 22036
rect 20524 20524 20580 20580
rect 20412 19740 20468 19796
rect 20412 18956 20468 19012
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 20972 19906 21028 19908
rect 20972 19854 20974 19906
rect 20974 19854 21026 19906
rect 21026 19854 21028 19906
rect 20972 19852 21028 19854
rect 21868 20748 21924 20804
rect 21644 20188 21700 20244
rect 23884 25228 23940 25284
rect 23436 24050 23492 24052
rect 23436 23998 23438 24050
rect 23438 23998 23490 24050
rect 23490 23998 23492 24050
rect 23436 23996 23492 23998
rect 22652 22316 22708 22372
rect 22540 22092 22596 22148
rect 22876 22428 22932 22484
rect 23100 23100 23156 23156
rect 22428 20130 22484 20132
rect 22428 20078 22430 20130
rect 22430 20078 22482 20130
rect 22482 20078 22484 20130
rect 22428 20076 22484 20078
rect 22204 19852 22260 19908
rect 21420 19180 21476 19236
rect 19292 18396 19348 18452
rect 19628 18450 19684 18452
rect 19628 18398 19630 18450
rect 19630 18398 19682 18450
rect 19682 18398 19684 18450
rect 19628 18396 19684 18398
rect 20636 18396 20692 18452
rect 19628 17724 19684 17780
rect 19292 17500 19348 17556
rect 18396 15986 18452 15988
rect 18396 15934 18398 15986
rect 18398 15934 18450 15986
rect 18450 15934 18452 15986
rect 18396 15932 18452 15934
rect 18508 15484 18564 15540
rect 18396 15148 18452 15204
rect 18172 15036 18228 15092
rect 20076 17666 20132 17668
rect 20076 17614 20078 17666
rect 20078 17614 20130 17666
rect 20130 17614 20132 17666
rect 20076 17612 20132 17614
rect 20636 17890 20692 17892
rect 20636 17838 20638 17890
rect 20638 17838 20690 17890
rect 20690 17838 20692 17890
rect 20636 17836 20692 17838
rect 21308 17778 21364 17780
rect 21308 17726 21310 17778
rect 21310 17726 21362 17778
rect 21362 17726 21364 17778
rect 21308 17724 21364 17726
rect 20748 17666 20804 17668
rect 20748 17614 20750 17666
rect 20750 17614 20802 17666
rect 20802 17614 20804 17666
rect 20748 17612 20804 17614
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 20636 16828 20692 16884
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 20188 15538 20244 15540
rect 20188 15486 20190 15538
rect 20190 15486 20242 15538
rect 20242 15486 20244 15538
rect 20188 15484 20244 15486
rect 21644 17554 21700 17556
rect 21644 17502 21646 17554
rect 21646 17502 21698 17554
rect 21698 17502 21700 17554
rect 21644 17500 21700 17502
rect 22204 17836 22260 17892
rect 22652 21532 22708 21588
rect 24556 26402 24612 26404
rect 24556 26350 24558 26402
rect 24558 26350 24610 26402
rect 24610 26350 24612 26402
rect 24556 26348 24612 26350
rect 24220 26290 24276 26292
rect 24220 26238 24222 26290
rect 24222 26238 24274 26290
rect 24274 26238 24276 26290
rect 24220 26236 24276 26238
rect 25004 26012 25060 26068
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 25676 27074 25732 27076
rect 25676 27022 25678 27074
rect 25678 27022 25730 27074
rect 25730 27022 25732 27074
rect 25676 27020 25732 27022
rect 28588 27186 28644 27188
rect 28588 27134 28590 27186
rect 28590 27134 28642 27186
rect 28642 27134 28644 27186
rect 28588 27132 28644 27134
rect 26460 26962 26516 26964
rect 26460 26910 26462 26962
rect 26462 26910 26514 26962
rect 26514 26910 26516 26962
rect 26460 26908 26516 26910
rect 25340 26460 25396 26516
rect 26684 26460 26740 26516
rect 27580 26460 27636 26516
rect 37660 27074 37716 27076
rect 37660 27022 37662 27074
rect 37662 27022 37714 27074
rect 37714 27022 37716 27074
rect 37660 27020 37716 27022
rect 28588 26460 28644 26516
rect 39900 26796 39956 26852
rect 27804 26402 27860 26404
rect 27804 26350 27806 26402
rect 27806 26350 27858 26402
rect 27858 26350 27860 26402
rect 27804 26348 27860 26350
rect 37660 26290 37716 26292
rect 37660 26238 37662 26290
rect 37662 26238 37714 26290
rect 37714 26238 37716 26290
rect 37660 26236 37716 26238
rect 25116 25340 25172 25396
rect 40012 26236 40068 26292
rect 26572 26066 26628 26068
rect 26572 26014 26574 26066
rect 26574 26014 26626 26066
rect 26626 26014 26628 26066
rect 26572 26012 26628 26014
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 25452 25394 25508 25396
rect 25452 25342 25454 25394
rect 25454 25342 25506 25394
rect 25506 25342 25508 25394
rect 25452 25340 25508 25342
rect 25228 23826 25284 23828
rect 25228 23774 25230 23826
rect 25230 23774 25282 23826
rect 25282 23774 25284 23826
rect 25228 23772 25284 23774
rect 23996 23154 24052 23156
rect 23996 23102 23998 23154
rect 23998 23102 24050 23154
rect 24050 23102 24052 23154
rect 23996 23100 24052 23102
rect 24444 23154 24500 23156
rect 24444 23102 24446 23154
rect 24446 23102 24498 23154
rect 24498 23102 24500 23154
rect 24444 23100 24500 23102
rect 23996 22652 24052 22708
rect 23660 22540 23716 22596
rect 23548 22428 23604 22484
rect 23436 22370 23492 22372
rect 23436 22318 23438 22370
rect 23438 22318 23490 22370
rect 23490 22318 23492 22370
rect 23436 22316 23492 22318
rect 23884 22370 23940 22372
rect 23884 22318 23886 22370
rect 23886 22318 23938 22370
rect 23938 22318 23940 22370
rect 23884 22316 23940 22318
rect 23324 22092 23380 22148
rect 23100 20300 23156 20356
rect 22988 19964 23044 20020
rect 22428 19516 22484 19572
rect 22316 17500 22372 17556
rect 21868 16604 21924 16660
rect 19068 15148 19124 15204
rect 17052 14306 17108 14308
rect 17052 14254 17054 14306
rect 17054 14254 17106 14306
rect 17106 14254 17108 14306
rect 17052 14252 17108 14254
rect 19852 15314 19908 15316
rect 19852 15262 19854 15314
rect 19854 15262 19906 15314
rect 19906 15262 19908 15314
rect 19852 15260 19908 15262
rect 19516 15090 19572 15092
rect 19516 15038 19518 15090
rect 19518 15038 19570 15090
rect 19570 15038 19572 15090
rect 19516 15036 19572 15038
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 19404 13916 19460 13972
rect 20188 13916 20244 13972
rect 20300 12962 20356 12964
rect 20300 12910 20302 12962
rect 20302 12910 20354 12962
rect 20354 12910 20356 12962
rect 20300 12908 20356 12910
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 21980 15484 22036 15540
rect 23212 16828 23268 16884
rect 23548 20076 23604 20132
rect 24444 22316 24500 22372
rect 24332 22204 24388 22260
rect 24892 22540 24948 22596
rect 24668 22428 24724 22484
rect 24668 22204 24724 22260
rect 24556 21980 24612 22036
rect 24220 21756 24276 21812
rect 24332 21644 24388 21700
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 25228 22428 25284 22484
rect 24220 21420 24276 21476
rect 23996 21362 24052 21364
rect 23996 21310 23998 21362
rect 23998 21310 24050 21362
rect 24050 21310 24052 21362
rect 23996 21308 24052 21310
rect 23996 20748 24052 20804
rect 23996 19234 24052 19236
rect 23996 19182 23998 19234
rect 23998 19182 24050 19234
rect 24050 19182 24052 19234
rect 23996 19180 24052 19182
rect 23548 18620 23604 18676
rect 24556 20188 24612 20244
rect 24444 20076 24500 20132
rect 24556 19906 24612 19908
rect 24556 19854 24558 19906
rect 24558 19854 24610 19906
rect 24610 19854 24612 19906
rect 24556 19852 24612 19854
rect 24444 19740 24500 19796
rect 24444 19234 24500 19236
rect 24444 19182 24446 19234
rect 24446 19182 24498 19234
rect 24498 19182 24500 19234
rect 24444 19180 24500 19182
rect 24220 19010 24276 19012
rect 24220 18958 24222 19010
rect 24222 18958 24274 19010
rect 24274 18958 24276 19010
rect 24220 18956 24276 18958
rect 24444 18620 24500 18676
rect 23548 16770 23604 16772
rect 23548 16718 23550 16770
rect 23550 16718 23602 16770
rect 23602 16718 23604 16770
rect 23548 16716 23604 16718
rect 23100 16604 23156 16660
rect 25340 21474 25396 21476
rect 25340 21422 25342 21474
rect 25342 21422 25394 21474
rect 25394 21422 25396 21474
rect 25340 21420 25396 21422
rect 28588 24050 28644 24052
rect 28588 23998 28590 24050
rect 28590 23998 28642 24050
rect 28642 23998 28644 24050
rect 28588 23996 28644 23998
rect 26460 23826 26516 23828
rect 26460 23774 26462 23826
rect 26462 23774 26514 23826
rect 26514 23774 26516 23826
rect 26460 23772 26516 23774
rect 25564 22370 25620 22372
rect 25564 22318 25566 22370
rect 25566 22318 25618 22370
rect 25618 22318 25620 22370
rect 25564 22316 25620 22318
rect 25564 22092 25620 22148
rect 26124 22428 26180 22484
rect 26572 22370 26628 22372
rect 26572 22318 26574 22370
rect 26574 22318 26626 22370
rect 26626 22318 26628 22370
rect 26572 22316 26628 22318
rect 25900 22258 25956 22260
rect 25900 22206 25902 22258
rect 25902 22206 25954 22258
rect 25954 22206 25956 22258
rect 25900 22204 25956 22206
rect 26348 21586 26404 21588
rect 26348 21534 26350 21586
rect 26350 21534 26402 21586
rect 26402 21534 26404 21586
rect 26348 21532 26404 21534
rect 37660 23938 37716 23940
rect 37660 23886 37662 23938
rect 37662 23886 37714 23938
rect 37714 23886 37716 23938
rect 37660 23884 37716 23886
rect 40012 23548 40068 23604
rect 28812 23100 28868 23156
rect 37660 23154 37716 23156
rect 37660 23102 37662 23154
rect 37662 23102 37714 23154
rect 37714 23102 37716 23154
rect 37660 23100 37716 23102
rect 40012 22930 40068 22932
rect 40012 22878 40014 22930
rect 40014 22878 40066 22930
rect 40066 22878 40068 22930
rect 40012 22876 40068 22878
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 28588 22316 28644 22372
rect 26684 21980 26740 22036
rect 25788 20748 25844 20804
rect 28588 21532 28644 21588
rect 25004 19180 25060 19236
rect 24780 18396 24836 18452
rect 26460 20130 26516 20132
rect 26460 20078 26462 20130
rect 26462 20078 26514 20130
rect 26514 20078 26516 20130
rect 26460 20076 26516 20078
rect 26348 19740 26404 19796
rect 26460 19852 26516 19908
rect 37660 21586 37716 21588
rect 37660 21534 37662 21586
rect 37662 21534 37714 21586
rect 37714 21534 37716 21586
rect 37660 21532 37716 21534
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 40012 20860 40068 20916
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 28028 19292 28084 19348
rect 26124 18956 26180 19012
rect 24444 16994 24500 16996
rect 24444 16942 24446 16994
rect 24446 16942 24498 16994
rect 24498 16942 24500 16994
rect 24444 16940 24500 16942
rect 27916 18450 27972 18452
rect 27916 18398 27918 18450
rect 27918 18398 27970 18450
rect 27970 18398 27972 18450
rect 27916 18396 27972 18398
rect 28588 19346 28644 19348
rect 28588 19294 28590 19346
rect 28590 19294 28642 19346
rect 28642 19294 28644 19346
rect 28588 19292 28644 19294
rect 40012 19516 40068 19572
rect 37660 19292 37716 19348
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 26124 17778 26180 17780
rect 26124 17726 26126 17778
rect 26126 17726 26178 17778
rect 26178 17726 26180 17778
rect 26124 17724 26180 17726
rect 40012 18226 40068 18228
rect 40012 18174 40014 18226
rect 40014 18174 40066 18226
rect 40066 18174 40068 18226
rect 40012 18172 40068 18174
rect 37660 17724 37716 17780
rect 25340 16828 25396 16884
rect 24332 16770 24388 16772
rect 24332 16718 24334 16770
rect 24334 16718 24386 16770
rect 24386 16718 24388 16770
rect 24332 16716 24388 16718
rect 23772 16658 23828 16660
rect 23772 16606 23774 16658
rect 23774 16606 23826 16658
rect 23826 16606 23828 16658
rect 23772 16604 23828 16606
rect 21196 14588 21252 14644
rect 22092 14642 22148 14644
rect 22092 14590 22094 14642
rect 22094 14590 22146 14642
rect 22146 14590 22148 14642
rect 22092 14588 22148 14590
rect 23100 15314 23156 15316
rect 23100 15262 23102 15314
rect 23102 15262 23154 15314
rect 23154 15262 23156 15314
rect 23100 15260 23156 15262
rect 22428 14588 22484 14644
rect 22540 14306 22596 14308
rect 22540 14254 22542 14306
rect 22542 14254 22594 14306
rect 22594 14254 22596 14306
rect 22540 14252 22596 14254
rect 23996 14252 24052 14308
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 15484 5180 15540 5236
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 16716 5234 16772 5236
rect 16716 5182 16718 5234
rect 16718 5182 16770 5234
rect 16770 5182 16772 5234
rect 16716 5180 16772 5182
rect 21084 12908 21140 12964
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 20188 4060 20244 4116
rect 16828 3388 16884 3444
rect 18060 3388 18116 3444
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 20860 3612 20916 3668
rect 24220 14306 24276 14308
rect 24220 14254 24222 14306
rect 24222 14254 24274 14306
rect 24274 14254 24276 14306
rect 24220 14252 24276 14254
rect 25788 16940 25844 16996
rect 25788 16210 25844 16212
rect 25788 16158 25790 16210
rect 25790 16158 25842 16210
rect 25842 16158 25844 16210
rect 25788 16156 25844 16158
rect 26236 16828 26292 16884
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 28588 16156 28644 16212
rect 25452 14252 25508 14308
rect 23548 5180 23604 5236
rect 21420 4114 21476 4116
rect 21420 4062 21422 4114
rect 21422 4062 21474 4114
rect 21474 4062 21476 4114
rect 21420 4060 21476 4062
rect 22092 3666 22148 3668
rect 22092 3614 22094 3666
rect 22094 3614 22146 3666
rect 22146 3614 22148 3666
rect 22092 3612 22148 3614
rect 22876 3388 22932 3444
rect 24220 4060 24276 4116
rect 24780 5234 24836 5236
rect 24780 5182 24782 5234
rect 24782 5182 24834 5234
rect 24834 5182 24836 5234
rect 24780 5180 24836 5182
rect 26236 4114 26292 4116
rect 26236 4062 26238 4114
rect 26238 4062 26290 4114
rect 26290 4062 26292 4114
rect 26236 4060 26292 4062
rect 24892 3612 24948 3668
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 40236 11452 40292 11508
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 29372 3666 29428 3668
rect 29372 3614 29374 3666
rect 29374 3614 29426 3666
rect 29426 3614 29428 3666
rect 29372 3612 29428 3614
rect 25564 3388 25620 3444
<< metal3 >>
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 20850 38220 20860 38276
rect 20916 38220 22092 38276
rect 22148 38220 22158 38276
rect 24882 38220 24892 38276
rect 24948 38220 26124 38276
rect 26180 38220 26190 38276
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 19506 37436 19516 37492
rect 19572 37436 20748 37492
rect 20804 37436 20814 37492
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 17042 28588 17052 28644
rect 17108 28588 20076 28644
rect 20132 28588 20142 28644
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 18386 27692 18396 27748
rect 18452 27692 20748 27748
rect 20804 27692 20814 27748
rect 0 27636 800 27664
rect 0 27580 4172 27636
rect 4228 27580 4238 27636
rect 0 27552 800 27580
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 20850 27132 20860 27188
rect 20916 27132 21980 27188
rect 22036 27132 22046 27188
rect 28578 27132 28588 27188
rect 28644 27132 31948 27188
rect 31892 27076 31948 27132
rect 4274 27020 4284 27076
rect 4340 27020 12684 27076
rect 12740 27020 12750 27076
rect 17714 27020 17724 27076
rect 17780 27020 21756 27076
rect 21812 27020 21822 27076
rect 22418 27020 22428 27076
rect 22484 27020 25228 27076
rect 25284 27020 25676 27076
rect 25732 27020 25742 27076
rect 31892 27020 37660 27076
rect 37716 27020 37726 27076
rect 41200 26964 42000 26992
rect 20290 26908 20300 26964
rect 20356 26908 21308 26964
rect 21364 26908 21374 26964
rect 21970 26908 21980 26964
rect 22036 26908 23996 26964
rect 24052 26908 24062 26964
rect 25106 26908 25116 26964
rect 25172 26908 26460 26964
rect 26516 26908 26526 26964
rect 39900 26908 42000 26964
rect 39900 26852 39956 26908
rect 41200 26880 42000 26908
rect 15810 26796 15820 26852
rect 15876 26796 17052 26852
rect 17108 26796 17118 26852
rect 20402 26796 20412 26852
rect 20468 26796 21644 26852
rect 21700 26796 21710 26852
rect 39890 26796 39900 26852
rect 39956 26796 39966 26852
rect 20178 26684 20188 26740
rect 20244 26684 20860 26740
rect 20916 26684 20926 26740
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 14690 26572 14700 26628
rect 14756 26572 15260 26628
rect 15316 26572 18844 26628
rect 18900 26572 18910 26628
rect 18844 26516 18900 26572
rect 14578 26460 14588 26516
rect 14644 26460 15932 26516
rect 15988 26460 15998 26516
rect 18844 26460 21028 26516
rect 24434 26460 24444 26516
rect 24500 26460 25340 26516
rect 25396 26460 25406 26516
rect 26674 26460 26684 26516
rect 26740 26460 27580 26516
rect 27636 26460 28588 26516
rect 28644 26460 28654 26516
rect 20972 26404 21028 26460
rect 12674 26348 12684 26404
rect 12740 26348 16156 26404
rect 16212 26348 16222 26404
rect 19740 26348 20748 26404
rect 20804 26348 20814 26404
rect 20972 26348 24556 26404
rect 24612 26348 24622 26404
rect 27794 26348 27804 26404
rect 27860 26348 31948 26404
rect 0 26292 800 26320
rect 19740 26292 19796 26348
rect 31892 26292 31948 26348
rect 41200 26292 42000 26320
rect 0 26236 1932 26292
rect 1988 26236 1998 26292
rect 13682 26236 13692 26292
rect 13748 26236 15484 26292
rect 15540 26236 15550 26292
rect 19058 26236 19068 26292
rect 19124 26236 19740 26292
rect 19796 26236 19806 26292
rect 20178 26236 20188 26292
rect 20244 26236 20972 26292
rect 21028 26236 21038 26292
rect 23090 26236 23100 26292
rect 23156 26236 24220 26292
rect 24276 26236 24286 26292
rect 31892 26236 37660 26292
rect 37716 26236 37726 26292
rect 40002 26236 40012 26292
rect 40068 26236 42000 26292
rect 0 26208 800 26236
rect 41200 26208 42000 26236
rect 24994 26012 25004 26068
rect 25060 26012 26572 26068
rect 26628 26012 26638 26068
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 14914 25676 14924 25732
rect 14980 25676 17500 25732
rect 17556 25676 17566 25732
rect 20962 25676 20972 25732
rect 21028 25676 22652 25732
rect 22708 25676 23660 25732
rect 23716 25676 23726 25732
rect 16482 25452 16492 25508
rect 16548 25452 17276 25508
rect 17332 25452 17342 25508
rect 18162 25452 18172 25508
rect 18228 25452 19292 25508
rect 19348 25452 19964 25508
rect 20020 25452 20030 25508
rect 19618 25340 19628 25396
rect 19684 25340 20412 25396
rect 20468 25340 22540 25396
rect 22596 25340 22606 25396
rect 23762 25340 23772 25396
rect 23828 25340 25116 25396
rect 25172 25340 25452 25396
rect 25508 25340 25518 25396
rect 19628 25228 19852 25284
rect 19908 25228 19918 25284
rect 21186 25228 21196 25284
rect 21252 25228 21980 25284
rect 22036 25228 22988 25284
rect 23044 25228 23884 25284
rect 23940 25228 23950 25284
rect 19628 25172 19684 25228
rect 17378 25116 17388 25172
rect 17444 25116 18844 25172
rect 18900 25116 19684 25172
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 19170 24892 19180 24948
rect 19236 24892 20300 24948
rect 20356 24892 20860 24948
rect 20916 24892 20926 24948
rect 16146 24668 16156 24724
rect 16212 24668 17612 24724
rect 17668 24668 17678 24724
rect 13906 24444 13916 24500
rect 13972 24444 15260 24500
rect 15316 24444 15326 24500
rect 19842 24444 19852 24500
rect 19908 24444 20636 24500
rect 20692 24444 20702 24500
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 17938 23996 17948 24052
rect 18004 23996 18956 24052
rect 19012 23996 23436 24052
rect 23492 23996 23502 24052
rect 28578 23996 28588 24052
rect 28644 23996 31948 24052
rect 31892 23940 31948 23996
rect 31892 23884 37660 23940
rect 37716 23884 37726 23940
rect 15362 23772 15372 23828
rect 15428 23772 16716 23828
rect 16772 23772 20636 23828
rect 20692 23772 20702 23828
rect 25218 23772 25228 23828
rect 25284 23772 26460 23828
rect 26516 23772 26526 23828
rect 41200 23604 42000 23632
rect 14354 23548 14364 23604
rect 14420 23548 15372 23604
rect 15428 23548 16156 23604
rect 16212 23548 16222 23604
rect 40002 23548 40012 23604
rect 40068 23548 42000 23604
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 41200 23520 42000 23548
rect 18162 23436 18172 23492
rect 18228 23436 19628 23492
rect 19684 23436 19694 23492
rect 16594 23324 16604 23380
rect 16660 23324 17724 23380
rect 17780 23324 18396 23380
rect 18452 23324 19180 23380
rect 19236 23324 20188 23380
rect 20244 23324 20254 23380
rect 19394 23212 19404 23268
rect 19460 23212 20300 23268
rect 20356 23212 21308 23268
rect 21364 23212 21374 23268
rect 23090 23100 23100 23156
rect 23156 23100 23996 23156
rect 24052 23100 24062 23156
rect 24434 23100 24444 23156
rect 24500 23100 28812 23156
rect 28868 23100 37660 23156
rect 37716 23100 37726 23156
rect 11666 22988 11676 23044
rect 11732 22988 13580 23044
rect 13636 22988 13646 23044
rect 13794 22988 13804 23044
rect 13860 22988 14476 23044
rect 14532 22988 15596 23044
rect 15652 22988 16268 23044
rect 16324 22988 16334 23044
rect 41200 22932 42000 22960
rect 18050 22876 18060 22932
rect 18116 22876 21532 22932
rect 21588 22876 21598 22932
rect 40002 22876 40012 22932
rect 40068 22876 42000 22932
rect 41200 22848 42000 22876
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 17714 22652 17724 22708
rect 17780 22652 18396 22708
rect 18452 22652 19516 22708
rect 19572 22652 19582 22708
rect 23958 22652 23996 22708
rect 24052 22652 24062 22708
rect 10770 22540 10780 22596
rect 10836 22540 18844 22596
rect 18900 22540 18910 22596
rect 20290 22540 20300 22596
rect 20356 22540 23660 22596
rect 23716 22540 24892 22596
rect 24948 22540 24958 22596
rect 18722 22428 18732 22484
rect 18788 22428 22876 22484
rect 22932 22428 22942 22484
rect 23538 22428 23548 22484
rect 23604 22428 24668 22484
rect 24724 22428 24734 22484
rect 25218 22428 25228 22484
rect 25284 22428 26124 22484
rect 26180 22428 26190 22484
rect 10098 22316 10108 22372
rect 10164 22316 10892 22372
rect 10948 22316 13132 22372
rect 13188 22316 14364 22372
rect 14420 22316 14430 22372
rect 14802 22316 14812 22372
rect 14868 22316 15932 22372
rect 15988 22316 16380 22372
rect 16436 22316 17388 22372
rect 17444 22316 17454 22372
rect 18610 22316 18620 22372
rect 18676 22316 19516 22372
rect 19572 22316 21420 22372
rect 21476 22316 21486 22372
rect 21634 22316 21644 22372
rect 21700 22316 22652 22372
rect 22708 22316 23436 22372
rect 23492 22316 23502 22372
rect 23846 22316 23884 22372
rect 23940 22316 23950 22372
rect 24434 22316 24444 22372
rect 24500 22316 25564 22372
rect 25620 22316 25630 22372
rect 26562 22316 26572 22372
rect 26628 22316 28588 22372
rect 28644 22316 28654 22372
rect 23436 22260 23492 22316
rect 14242 22204 14252 22260
rect 14308 22204 14700 22260
rect 14756 22204 18508 22260
rect 18564 22204 18574 22260
rect 23436 22204 24332 22260
rect 24388 22204 24398 22260
rect 24658 22204 24668 22260
rect 24724 22204 25900 22260
rect 25956 22204 25966 22260
rect 16482 22092 16492 22148
rect 16548 22092 17500 22148
rect 17556 22092 18732 22148
rect 18788 22092 18798 22148
rect 20402 22092 20412 22148
rect 20468 22092 22540 22148
rect 22596 22092 23324 22148
rect 23380 22092 25564 22148
rect 25620 22092 25630 22148
rect 20850 21980 20860 22036
rect 20916 21980 24556 22036
rect 24612 21980 26684 22036
rect 26740 21980 26750 22036
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 16818 21868 16828 21924
rect 16884 21868 17724 21924
rect 17780 21868 17790 21924
rect 19618 21868 19628 21924
rect 19684 21868 19694 21924
rect 19628 21812 19684 21868
rect 15138 21756 15148 21812
rect 15204 21756 16940 21812
rect 16996 21756 20300 21812
rect 20356 21756 20366 21812
rect 24210 21756 24220 21812
rect 24276 21756 28644 21812
rect 12898 21644 12908 21700
rect 12964 21644 14364 21700
rect 14420 21644 14812 21700
rect 14868 21644 14878 21700
rect 15810 21644 15820 21700
rect 15876 21644 24332 21700
rect 24388 21644 24398 21700
rect 28588 21588 28644 21756
rect 22642 21532 22652 21588
rect 22708 21532 26348 21588
rect 26404 21532 26414 21588
rect 28578 21532 28588 21588
rect 28644 21532 37660 21588
rect 37716 21532 37726 21588
rect 4162 21420 4172 21476
rect 4228 21420 17836 21476
rect 17892 21420 17902 21476
rect 24210 21420 24220 21476
rect 24276 21420 25340 21476
rect 25396 21420 25406 21476
rect 23958 21308 23996 21364
rect 24052 21308 24062 21364
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 41200 20916 42000 20944
rect 40002 20860 40012 20916
rect 40068 20860 42000 20916
rect 41200 20832 42000 20860
rect 17490 20748 17500 20804
rect 17556 20748 19628 20804
rect 19684 20748 19694 20804
rect 21858 20748 21868 20804
rect 21924 20748 23996 20804
rect 24052 20748 25788 20804
rect 25844 20748 25854 20804
rect 19394 20524 19404 20580
rect 19460 20524 20524 20580
rect 20580 20524 20590 20580
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 23090 20300 23100 20356
rect 23156 20300 23884 20356
rect 23940 20300 23950 20356
rect 0 20244 800 20272
rect 0 20188 1932 20244
rect 1988 20188 1998 20244
rect 19842 20188 19852 20244
rect 19908 20188 21644 20244
rect 21700 20188 21710 20244
rect 24220 20188 24556 20244
rect 24612 20188 24622 20244
rect 0 20160 800 20188
rect 24220 20132 24276 20188
rect 14354 20076 14364 20132
rect 14420 20076 15484 20132
rect 15540 20076 15550 20132
rect 16258 20076 16268 20132
rect 16324 20076 17500 20132
rect 17556 20076 17566 20132
rect 22418 20076 22428 20132
rect 22484 20076 23548 20132
rect 23604 20076 24276 20132
rect 24434 20076 24444 20132
rect 24500 20076 26460 20132
rect 26516 20076 26526 20132
rect 4274 19964 4284 20020
rect 4340 19964 12460 20020
rect 12516 19964 12526 20020
rect 16594 19964 16604 20020
rect 16660 19964 18732 20020
rect 18788 19964 18798 20020
rect 18956 19964 22988 20020
rect 23044 19964 23054 20020
rect 18956 19908 19012 19964
rect 11778 19852 11788 19908
rect 11844 19852 14364 19908
rect 14420 19852 14430 19908
rect 15138 19852 15148 19908
rect 15204 19852 16828 19908
rect 16884 19852 17724 19908
rect 17780 19852 19012 19908
rect 20962 19852 20972 19908
rect 21028 19852 22204 19908
rect 22260 19852 22270 19908
rect 24546 19852 24556 19908
rect 24612 19852 26460 19908
rect 26516 19852 26526 19908
rect 1922 19740 1932 19796
rect 1988 19740 1998 19796
rect 20402 19740 20412 19796
rect 20468 19740 24444 19796
rect 24500 19740 26348 19796
rect 26404 19740 26414 19796
rect 0 19572 800 19600
rect 1932 19572 1988 19740
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 41200 19572 42000 19600
rect 0 19516 1988 19572
rect 15026 19516 15036 19572
rect 15092 19516 22428 19572
rect 22484 19516 22494 19572
rect 40002 19516 40012 19572
rect 40068 19516 42000 19572
rect 0 19488 800 19516
rect 41200 19488 42000 19516
rect 4162 19292 4172 19348
rect 4228 19292 9884 19348
rect 9940 19292 12684 19348
rect 12740 19292 13692 19348
rect 13748 19292 14140 19348
rect 14196 19292 14206 19348
rect 28018 19292 28028 19348
rect 28084 19292 28588 19348
rect 28644 19292 37660 19348
rect 37716 19292 37726 19348
rect 4274 19180 4284 19236
rect 4340 19180 13468 19236
rect 13524 19180 13534 19236
rect 21410 19180 21420 19236
rect 21476 19180 23996 19236
rect 24052 19180 24062 19236
rect 24434 19180 24444 19236
rect 24500 19180 25004 19236
rect 25060 19180 25070 19236
rect 13906 18956 13916 19012
rect 13972 18956 14924 19012
rect 14980 18956 20412 19012
rect 20468 18956 20478 19012
rect 24210 18956 24220 19012
rect 24276 18956 26124 19012
rect 26180 18956 26190 19012
rect 0 18900 800 18928
rect 0 18844 1932 18900
rect 1988 18844 1998 18900
rect 0 18816 800 18844
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 23538 18620 23548 18676
rect 23604 18620 24444 18676
rect 24500 18620 24510 18676
rect 4274 18396 4284 18452
rect 4340 18396 8428 18452
rect 12898 18396 12908 18452
rect 12964 18396 14028 18452
rect 14084 18396 16604 18452
rect 16660 18396 17500 18452
rect 17556 18396 17566 18452
rect 18498 18396 18508 18452
rect 18564 18396 19292 18452
rect 19348 18396 19358 18452
rect 19618 18396 19628 18452
rect 19684 18396 20636 18452
rect 20692 18396 20702 18452
rect 24770 18396 24780 18452
rect 24836 18396 27916 18452
rect 27972 18396 27982 18452
rect 8372 18340 8428 18396
rect 8372 18284 13692 18340
rect 13748 18284 15148 18340
rect 0 18228 800 18256
rect 15092 18228 15148 18284
rect 41200 18228 42000 18256
rect 0 18172 1932 18228
rect 1988 18172 1998 18228
rect 15092 18172 16380 18228
rect 16436 18172 16446 18228
rect 40002 18172 40012 18228
rect 40068 18172 42000 18228
rect 0 18144 800 18172
rect 41200 18144 42000 18172
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 15586 17836 15596 17892
rect 15652 17836 16268 17892
rect 16324 17836 16334 17892
rect 20626 17836 20636 17892
rect 20692 17836 22204 17892
rect 22260 17836 22270 17892
rect 19618 17724 19628 17780
rect 19684 17724 21308 17780
rect 21364 17724 21374 17780
rect 26114 17724 26124 17780
rect 26180 17724 37660 17780
rect 37716 17724 37726 17780
rect 4274 17612 4284 17668
rect 4340 17612 11116 17668
rect 11172 17612 11182 17668
rect 20066 17612 20076 17668
rect 20132 17612 20748 17668
rect 20804 17612 20814 17668
rect 19282 17500 19292 17556
rect 19348 17500 21644 17556
rect 21700 17500 22316 17556
rect 22372 17500 22382 17556
rect 13234 17388 13244 17444
rect 13300 17388 14364 17444
rect 14420 17388 14430 17444
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 11106 17052 11116 17108
rect 11172 17052 14588 17108
rect 14644 17052 14654 17108
rect 24434 16940 24444 16996
rect 24500 16940 25788 16996
rect 25844 16940 25854 16996
rect 0 16884 800 16912
rect 0 16828 1932 16884
rect 1988 16828 1998 16884
rect 14914 16828 14924 16884
rect 14980 16828 15148 16884
rect 15204 16828 20636 16884
rect 20692 16828 20702 16884
rect 23202 16828 23212 16884
rect 23268 16828 25340 16884
rect 25396 16828 26236 16884
rect 26292 16828 26302 16884
rect 0 16800 800 16828
rect 14354 16716 14364 16772
rect 14420 16716 15036 16772
rect 15092 16716 15102 16772
rect 23538 16716 23548 16772
rect 23604 16716 24332 16772
rect 24388 16716 24398 16772
rect 21858 16604 21868 16660
rect 21924 16604 23100 16660
rect 23156 16604 23772 16660
rect 23828 16604 23838 16660
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 25778 16156 25788 16212
rect 25844 16156 28588 16212
rect 28644 16156 28654 16212
rect 17378 15932 17388 15988
rect 17444 15932 18396 15988
rect 18452 15932 18462 15988
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 16370 15484 16380 15540
rect 16436 15484 18508 15540
rect 18564 15484 20188 15540
rect 20244 15484 21980 15540
rect 22036 15484 22046 15540
rect 15138 15260 15148 15316
rect 15204 15260 16044 15316
rect 16100 15260 16828 15316
rect 16884 15260 16894 15316
rect 19842 15260 19852 15316
rect 19908 15260 23100 15316
rect 23156 15260 23166 15316
rect 14354 15148 14364 15204
rect 14420 15148 15260 15204
rect 15316 15148 15326 15204
rect 15586 15148 15596 15204
rect 15652 15148 17500 15204
rect 17556 15148 18396 15204
rect 18452 15148 19068 15204
rect 19124 15148 19134 15204
rect 17042 15036 17052 15092
rect 17108 15036 18172 15092
rect 18228 15036 19516 15092
rect 19572 15036 19582 15092
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 21186 14588 21196 14644
rect 21252 14588 22092 14644
rect 22148 14588 22428 14644
rect 22484 14588 22494 14644
rect 14690 14252 14700 14308
rect 14756 14252 17052 14308
rect 17108 14252 17118 14308
rect 22530 14252 22540 14308
rect 22596 14252 23996 14308
rect 24052 14252 24062 14308
rect 24210 14252 24220 14308
rect 24276 14252 25452 14308
rect 25508 14252 25518 14308
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 19394 13916 19404 13972
rect 19460 13916 20188 13972
rect 20244 13916 20254 13972
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 20290 12908 20300 12964
rect 20356 12908 21084 12964
rect 21140 12908 21150 12964
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 41200 11508 42000 11536
rect 40226 11452 40236 11508
rect 40292 11452 42000 11508
rect 41200 11424 42000 11452
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 15474 5180 15484 5236
rect 15540 5180 16716 5236
rect 16772 5180 16782 5236
rect 23538 5180 23548 5236
rect 23604 5180 24780 5236
rect 24836 5180 24846 5236
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 20178 4060 20188 4116
rect 20244 4060 21420 4116
rect 21476 4060 21486 4116
rect 24210 4060 24220 4116
rect 24276 4060 26236 4116
rect 26292 4060 26302 4116
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 20850 3612 20860 3668
rect 20916 3612 22092 3668
rect 22148 3612 22158 3668
rect 24882 3612 24892 3668
rect 24948 3612 29372 3668
rect 29428 3612 29438 3668
rect 16818 3388 16828 3444
rect 16884 3388 18060 3444
rect 18116 3388 18126 3444
rect 22866 3388 22876 3444
rect 22932 3388 25564 3444
rect 25620 3388 25630 3444
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
<< via3 >>
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 23996 22652 24052 22708
rect 23884 22316 23940 22372
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 23996 21308 24052 21364
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 23884 20300 23940 20356
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
<< metal4 >>
rect 4448 38444 4768 38476
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 37660 20128 38476
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19808 34524 20128 36036
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 19808 23548 20128 25060
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 19808 21980 20128 23492
rect 35168 38444 35488 38476
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 35168 22764 35488 24276
rect 23996 22708 24052 22718
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 23884 22372 23940 22382
rect 23884 20356 23940 22316
rect 23996 21364 24052 22652
rect 23996 21298 24052 21308
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 23884 20290 23940 20300
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _103_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 20944 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _104_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 22512 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _105_
timestamp 1698175906
transform -1 0 16576 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _106_
timestamp 1698175906
transform 1 0 14672 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _107_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 16800 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _108_
timestamp 1698175906
transform -1 0 19824 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _109_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 19824 0 -1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _110_
timestamp 1698175906
transform 1 0 17136 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _111_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 16128 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _112_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 18592 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _113_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 17024 0 -1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _114_
timestamp 1698175906
transform -1 0 15568 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _115_
timestamp 1698175906
transform -1 0 16912 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _116_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17248 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _117_
timestamp 1698175906
transform -1 0 16688 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _118_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 15344 0 -1 23520
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _119_
timestamp 1698175906
transform -1 0 14112 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _120_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17360 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _121_
timestamp 1698175906
transform 1 0 17808 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _122_
timestamp 1698175906
transform 1 0 19824 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _123_
timestamp 1698175906
transform 1 0 21168 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _124_
timestamp 1698175906
transform -1 0 19936 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _125_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18480 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _126_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 17248 0 1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _127_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 19152 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _128_
timestamp 1698175906
transform -1 0 17920 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _129_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18256 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _130_
timestamp 1698175906
transform 1 0 20944 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _131_
timestamp 1698175906
transform -1 0 21840 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _132_
timestamp 1698175906
transform 1 0 18928 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _133_
timestamp 1698175906
transform 1 0 21168 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _134_
timestamp 1698175906
transform 1 0 19824 0 -1 20384
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _135_
timestamp 1698175906
transform -1 0 22400 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _136_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 14672 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _137_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17808 0 1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _138_
timestamp 1698175906
transform 1 0 15344 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _139_
timestamp 1698175906
transform -1 0 24864 0 1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _140_
timestamp 1698175906
transform 1 0 23520 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _141_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 15568 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _142_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 15008 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _143_
timestamp 1698175906
transform -1 0 14560 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _144_
timestamp 1698175906
transform -1 0 20944 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _145_
timestamp 1698175906
transform -1 0 15344 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _146_
timestamp 1698175906
transform 1 0 20160 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _147_
timestamp 1698175906
transform 1 0 14224 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _148_
timestamp 1698175906
transform -1 0 14672 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _149_
timestamp 1698175906
transform -1 0 20496 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _150_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18928 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _151_
timestamp 1698175906
transform 1 0 14560 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _152_
timestamp 1698175906
transform 1 0 24080 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _153_
timestamp 1698175906
transform 1 0 19936 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _154_
timestamp 1698175906
transform 1 0 22400 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _155_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 23184 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _156_
timestamp 1698175906
transform -1 0 22512 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _157_
timestamp 1698175906
transform -1 0 23520 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _158_
timestamp 1698175906
transform 1 0 21168 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _159_
timestamp 1698175906
transform 1 0 22736 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _160_
timestamp 1698175906
transform -1 0 24304 0 1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _161_
timestamp 1698175906
transform -1 0 24752 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _162_
timestamp 1698175906
transform 1 0 22288 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _163_
timestamp 1698175906
transform 1 0 22512 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _164_
timestamp 1698175906
transform -1 0 15792 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _165_
timestamp 1698175906
transform -1 0 14896 0 -1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _166_
timestamp 1698175906
transform 1 0 11648 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _167_
timestamp 1698175906
transform -1 0 19264 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _168_
timestamp 1698175906
transform 1 0 23296 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _169_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 20944 0 1 20384
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _170_
timestamp 1698175906
transform 1 0 26096 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _171_
timestamp 1698175906
transform 1 0 18928 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _172_
timestamp 1698175906
transform 1 0 20272 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _173_
timestamp 1698175906
transform 1 0 23520 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _174_
timestamp 1698175906
transform -1 0 25536 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _175_
timestamp 1698175906
transform 1 0 23968 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _176_
timestamp 1698175906
transform 1 0 24304 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _177_
timestamp 1698175906
transform -1 0 26096 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _178_
timestamp 1698175906
transform -1 0 28224 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _179_
timestamp 1698175906
transform 1 0 25088 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _180_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 23632 0 -1 20384
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _181_
timestamp 1698175906
transform 1 0 20048 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _182_
timestamp 1698175906
transform -1 0 19936 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _183_
timestamp 1698175906
transform 1 0 19152 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _184_
timestamp 1698175906
transform -1 0 20496 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _185_
timestamp 1698175906
transform 1 0 19376 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _186_
timestamp 1698175906
transform 1 0 19376 0 -1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _187_
timestamp 1698175906
transform -1 0 22064 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _188_
timestamp 1698175906
transform -1 0 17696 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _189_
timestamp 1698175906
transform -1 0 17696 0 1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _190_
timestamp 1698175906
transform 1 0 20384 0 -1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _191_
timestamp 1698175906
transform -1 0 20944 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _192_
timestamp 1698175906
transform -1 0 26880 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _193_
timestamp 1698175906
transform -1 0 19376 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _194_
timestamp 1698175906
transform 1 0 22176 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _195_
timestamp 1698175906
transform -1 0 26544 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _196_
timestamp 1698175906
transform -1 0 25648 0 1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _197_
timestamp 1698175906
transform -1 0 16464 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _198_
timestamp 1698175906
transform 1 0 17248 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _199_
timestamp 1698175906
transform 1 0 13440 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _200_
timestamp 1698175906
transform 1 0 15120 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _201_
timestamp 1698175906
transform -1 0 15344 0 1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _202_
timestamp 1698175906
transform -1 0 24752 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _203_
timestamp 1698175906
transform 1 0 22288 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _204_
timestamp 1698175906
transform -1 0 23408 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _205_
timestamp 1698175906
transform -1 0 23520 0 -1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _206_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 16800 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _207_
timestamp 1698175906
transform 1 0 13440 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _208_
timestamp 1698175906
transform 1 0 10752 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _209_
timestamp 1698175906
transform 1 0 9856 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _210_
timestamp 1698175906
transform 1 0 17808 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _211_
timestamp 1698175906
transform 1 0 23072 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _212_
timestamp 1698175906
transform 1 0 13328 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _213_
timestamp 1698175906
transform -1 0 14224 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _214_
timestamp 1698175906
transform 1 0 17920 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _215_
timestamp 1698175906
transform 1 0 22736 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _216_
timestamp 1698175906
transform 1 0 25536 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _217_
timestamp 1698175906
transform 1 0 21616 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _218_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 13104 0 1 18816
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _219_
timestamp 1698175906
transform 1 0 25536 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _220_
timestamp 1698175906
transform 1 0 25760 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _221_
timestamp 1698175906
transform 1 0 25536 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _222_
timestamp 1698175906
transform 1 0 17696 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _223_
timestamp 1698175906
transform 1 0 16800 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _224_
timestamp 1698175906
transform 1 0 13776 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _225_
timestamp 1698175906
transform -1 0 21504 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _226_
timestamp 1698175906
transform 1 0 25536 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _227_
timestamp 1698175906
transform -1 0 15792 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _228_
timestamp 1698175906
transform 1 0 22288 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _231_
timestamp 1698175906
transform -1 0 24416 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _232_
timestamp 1698175906
transform -1 0 14000 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _233_
timestamp 1698175906
transform 1 0 27328 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _234_
timestamp 1698175906
transform 1 0 23744 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _235_
timestamp 1698175906
transform -1 0 12992 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__147__B dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 15344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__162__A2
timestamp 1698175906
transform 1 0 22064 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__181__B
timestamp 1698175906
transform 1 0 21168 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__197__A2
timestamp 1698175906
transform 1 0 16688 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__206__CLK
timestamp 1698175906
transform 1 0 17472 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__207__CLK
timestamp 1698175906
transform 1 0 16912 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__208__CLK
timestamp 1698175906
transform 1 0 14336 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__209__CLK
timestamp 1698175906
transform 1 0 13104 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__210__CLK
timestamp 1698175906
transform 1 0 17584 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__211__CLK
timestamp 1698175906
transform 1 0 26544 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__212__CLK
timestamp 1698175906
transform 1 0 16576 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__213__CLK
timestamp 1698175906
transform 1 0 14224 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__214__CLK
timestamp 1698175906
transform -1 0 17920 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__215__CLK
timestamp 1698175906
transform 1 0 26208 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__216__CLK
timestamp 1698175906
transform 1 0 25312 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__217__CLK
timestamp 1698175906
transform 1 0 25312 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__218__CLK
timestamp 1698175906
transform 1 0 13104 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__219__CLK
timestamp 1698175906
transform 1 0 25312 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__220__CLK
timestamp 1698175906
transform 1 0 25536 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__221__CLK
timestamp 1698175906
transform 1 0 25312 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__222__CLK
timestamp 1698175906
transform 1 0 17472 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__223__CLK
timestamp 1698175906
transform 1 0 20048 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__224__CLK
timestamp 1698175906
transform -1 0 17248 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__225__CLK
timestamp 1698175906
transform -1 0 21952 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__226__CLK
timestamp 1698175906
transform 1 0 25312 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__227__CLK
timestamp 1698175906
transform 1 0 15792 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__228__CLK
timestamp 1698175906
transform -1 0 25760 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1698175906
transform 1 0 17808 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18032 0 -1 21952
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1698175906
transform -1 0 20944 0 1 18816
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1698175906
transform 1 0 21504 0 1 20384
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1568 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698175906
transform 1 0 5376 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698175906
transform 1 0 9184 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698175906
transform 1 0 12992 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_138 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 16800 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_165 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19824 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_169
timestamp 1698175906
transform 1 0 20272 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_172 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 20608 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_174
timestamp 1698175906
transform 1 0 20832 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_201
timestamp 1698175906
transform 1 0 23856 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_203
timestamp 1698175906
transform 1 0 24080 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_232
timestamp 1698175906
transform 1 0 27328 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_236
timestamp 1698175906
transform 1 0 27776 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_266
timestamp 1698175906
transform 1 0 31136 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_270
timestamp 1698175906
transform 1 0 31584 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_274
timestamp 1698175906
transform 1 0 32032 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_308
timestamp 1698175906
transform 1 0 35840 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_342
timestamp 1698175906
transform 1 0 39648 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_346
timestamp 1698175906
transform 1 0 40096 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_348
timestamp 1698175906
transform 1 0 40320 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1568 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698175906
transform 1 0 8736 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698175906
transform 1 0 9408 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698175906
transform 1 0 16576 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_142 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17248 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_158 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19040 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_166
timestamp 1698175906
transform 1 0 19936 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_168
timestamp 1698175906
transform 1 0 20160 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_195
timestamp 1698175906
transform 1 0 23184 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_203
timestamp 1698175906
transform 1 0 24080 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_207
timestamp 1698175906
transform 1 0 24528 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_209
timestamp 1698175906
transform 1 0 24752 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_238
timestamp 1698175906
transform 1 0 28000 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_270
timestamp 1698175906
transform 1 0 31584 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_278
timestamp 1698175906
transform 1 0 32480 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_282
timestamp 1698175906
transform 1 0 32928 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_346
timestamp 1698175906
transform 1 0 40096 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_348
timestamp 1698175906
transform 1 0 40320 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698175906
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698175906
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698175906
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698175906
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_107
timestamp 1698175906
transform 1 0 13328 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_123
timestamp 1698175906
transform 1 0 15120 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_153
timestamp 1698175906
transform 1 0 18480 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_169
timestamp 1698175906
transform 1 0 20272 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_173
timestamp 1698175906
transform 1 0 20720 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_177
timestamp 1698175906
transform 1 0 21168 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_193
timestamp 1698175906
transform 1 0 22960 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_197
timestamp 1698175906
transform 1 0 23408 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_225
timestamp 1698175906
transform 1 0 26544 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_241
timestamp 1698175906
transform 1 0 28336 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698175906
transform 1 0 29008 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698175906
transform 1 0 36176 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_317
timestamp 1698175906
transform 1 0 36848 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698175906
transform 1 0 1568 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698175906
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698175906
transform 1 0 9408 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698175906
transform 1 0 16576 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_142
timestamp 1698175906
transform 1 0 17248 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_206
timestamp 1698175906
transform 1 0 24416 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_212
timestamp 1698175906
transform 1 0 25088 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_276
timestamp 1698175906
transform 1 0 32256 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_282
timestamp 1698175906
transform 1 0 32928 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_346
timestamp 1698175906
transform 1 0 40096 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_348
timestamp 1698175906
transform 1 0 40320 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698175906
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698175906
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698175906
transform 1 0 5488 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698175906
transform 1 0 12656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_107
timestamp 1698175906
transform 1 0 13328 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698175906
transform 1 0 20496 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_177
timestamp 1698175906
transform 1 0 21168 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_241
timestamp 1698175906
transform 1 0 28336 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698175906
transform 1 0 29008 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698175906
transform 1 0 36176 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_317
timestamp 1698175906
transform 1 0 36848 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698175906
transform 1 0 1568 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698175906
transform 1 0 8736 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698175906
transform 1 0 9408 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698175906
transform 1 0 16576 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_142
timestamp 1698175906
transform 1 0 17248 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_206
timestamp 1698175906
transform 1 0 24416 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_212
timestamp 1698175906
transform 1 0 25088 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698175906
transform 1 0 32256 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_282
timestamp 1698175906
transform 1 0 32928 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_346
timestamp 1698175906
transform 1 0 40096 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_348
timestamp 1698175906
transform 1 0 40320 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698175906
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698175906
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698175906
transform 1 0 5488 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698175906
transform 1 0 12656 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_107
timestamp 1698175906
transform 1 0 13328 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_171
timestamp 1698175906
transform 1 0 20496 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_177
timestamp 1698175906
transform 1 0 21168 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_241
timestamp 1698175906
transform 1 0 28336 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_247
timestamp 1698175906
transform 1 0 29008 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_311
timestamp 1698175906
transform 1 0 36176 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_317
timestamp 1698175906
transform 1 0 36848 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698175906
transform 1 0 1568 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698175906
transform 1 0 8736 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_72
timestamp 1698175906
transform 1 0 9408 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698175906
transform 1 0 16576 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_142
timestamp 1698175906
transform 1 0 17248 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_206
timestamp 1698175906
transform 1 0 24416 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_212
timestamp 1698175906
transform 1 0 25088 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_276
timestamp 1698175906
transform 1 0 32256 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_282
timestamp 1698175906
transform 1 0 32928 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_346
timestamp 1698175906
transform 1 0 40096 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_348
timestamp 1698175906
transform 1 0 40320 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698175906
transform 1 0 1568 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698175906
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_37
timestamp 1698175906
transform 1 0 5488 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_101
timestamp 1698175906
transform 1 0 12656 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_107
timestamp 1698175906
transform 1 0 13328 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_171
timestamp 1698175906
transform 1 0 20496 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_177
timestamp 1698175906
transform 1 0 21168 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_241
timestamp 1698175906
transform 1 0 28336 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_247
timestamp 1698175906
transform 1 0 29008 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_311
timestamp 1698175906
transform 1 0 36176 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_317
timestamp 1698175906
transform 1 0 36848 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698175906
transform 1 0 1568 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698175906
transform 1 0 8736 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_72
timestamp 1698175906
transform 1 0 9408 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_136
timestamp 1698175906
transform 1 0 16576 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_142
timestamp 1698175906
transform 1 0 17248 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_206
timestamp 1698175906
transform 1 0 24416 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_212
timestamp 1698175906
transform 1 0 25088 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_276
timestamp 1698175906
transform 1 0 32256 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_282
timestamp 1698175906
transform 1 0 32928 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_346
timestamp 1698175906
transform 1 0 40096 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_348
timestamp 1698175906
transform 1 0 40320 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698175906
transform 1 0 1568 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698175906
transform 1 0 5152 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_37
timestamp 1698175906
transform 1 0 5488 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698175906
transform 1 0 12656 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_107
timestamp 1698175906
transform 1 0 13328 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_171
timestamp 1698175906
transform 1 0 20496 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_177
timestamp 1698175906
transform 1 0 21168 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_241
timestamp 1698175906
transform 1 0 28336 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_247
timestamp 1698175906
transform 1 0 29008 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_311
timestamp 1698175906
transform 1 0 36176 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_317
timestamp 1698175906
transform 1 0 36848 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2
timestamp 1698175906
transform 1 0 1568 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698175906
transform 1 0 8736 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_72
timestamp 1698175906
transform 1 0 9408 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698175906
transform 1 0 16576 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_142
timestamp 1698175906
transform 1 0 17248 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_206
timestamp 1698175906
transform 1 0 24416 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_212
timestamp 1698175906
transform 1 0 25088 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_276
timestamp 1698175906
transform 1 0 32256 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_11_282
timestamp 1698175906
transform 1 0 32928 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_314
timestamp 1698175906
transform 1 0 36512 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_330
timestamp 1698175906
transform 1 0 38304 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_338
timestamp 1698175906
transform 1 0 39200 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_342
timestamp 1698175906
transform 1 0 39648 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_344
timestamp 1698175906
transform 1 0 39872 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698175906
transform 1 0 1568 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698175906
transform 1 0 5152 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_37
timestamp 1698175906
transform 1 0 5488 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698175906
transform 1 0 12656 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_107
timestamp 1698175906
transform 1 0 13328 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_139
timestamp 1698175906
transform 1 0 16912 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_142
timestamp 1698175906
transform 1 0 17248 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_148
timestamp 1698175906
transform 1 0 17920 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_164
timestamp 1698175906
transform 1 0 19712 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_166
timestamp 1698175906
transform 1 0 19936 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_171
timestamp 1698175906
transform 1 0 20496 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_177
timestamp 1698175906
transform 1 0 21168 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_193
timestamp 1698175906
transform 1 0 22960 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_197
timestamp 1698175906
transform 1 0 23408 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_199
timestamp 1698175906
transform 1 0 23632 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_206
timestamp 1698175906
transform 1 0 24416 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_238
timestamp 1698175906
transform 1 0 28000 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_242
timestamp 1698175906
transform 1 0 28448 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_244
timestamp 1698175906
transform 1 0 28672 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_247
timestamp 1698175906
transform 1 0 29008 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_311
timestamp 1698175906
transform 1 0 36176 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_317
timestamp 1698175906
transform 1 0 36848 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_2
timestamp 1698175906
transform 1 0 1568 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_66
timestamp 1698175906
transform 1 0 8736 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_72
timestamp 1698175906
transform 1 0 9408 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_104
timestamp 1698175906
transform 1 0 12992 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_108
timestamp 1698175906
transform 1 0 13440 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_110
timestamp 1698175906
transform 1 0 13664 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_146
timestamp 1698175906
transform 1 0 17696 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_177
timestamp 1698175906
transform 1 0 21168 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_212
timestamp 1698175906
transform 1 0 25088 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_216
timestamp 1698175906
transform 1 0 25536 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_282
timestamp 1698175906
transform 1 0 32928 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_346
timestamp 1698175906
transform 1 0 40096 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_348
timestamp 1698175906
transform 1 0 40320 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698175906
transform 1 0 1568 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698175906
transform 1 0 5152 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_37
timestamp 1698175906
transform 1 0 5488 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_101
timestamp 1698175906
transform 1 0 12656 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_177
timestamp 1698175906
transform 1 0 21168 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_192
timestamp 1698175906
transform 1 0 22848 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_206
timestamp 1698175906
transform 1 0 24416 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_238
timestamp 1698175906
transform 1 0 28000 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_242
timestamp 1698175906
transform 1 0 28448 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_244
timestamp 1698175906
transform 1 0 28672 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_247
timestamp 1698175906
transform 1 0 29008 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_311
timestamp 1698175906
transform 1 0 36176 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_317
timestamp 1698175906
transform 1 0 36848 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_2
timestamp 1698175906
transform 1 0 1568 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_66
timestamp 1698175906
transform 1 0 8736 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_72
timestamp 1698175906
transform 1 0 9408 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_104
timestamp 1698175906
transform 1 0 12992 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_112
timestamp 1698175906
transform 1 0 13888 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_118
timestamp 1698175906
transform 1 0 14560 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_132
timestamp 1698175906
transform 1 0 16128 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_138
timestamp 1698175906
transform 1 0 16800 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_142
timestamp 1698175906
transform 1 0 17248 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_146
timestamp 1698175906
transform 1 0 17696 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_154
timestamp 1698175906
transform 1 0 18592 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_156
timestamp 1698175906
transform 1 0 18816 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_175
timestamp 1698175906
transform 1 0 20944 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_179
timestamp 1698175906
transform 1 0 21392 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_187
timestamp 1698175906
transform 1 0 22288 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_197
timestamp 1698175906
transform 1 0 23408 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_205
timestamp 1698175906
transform 1 0 24304 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_209
timestamp 1698175906
transform 1 0 24752 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_212
timestamp 1698175906
transform 1 0 25088 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_276
timestamp 1698175906
transform 1 0 32256 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_282
timestamp 1698175906
transform 1 0 32928 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_346
timestamp 1698175906
transform 1 0 40096 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_348
timestamp 1698175906
transform 1 0 40320 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_2
timestamp 1698175906
transform 1 0 1568 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698175906
transform 1 0 5152 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_37
timestamp 1698175906
transform 1 0 5488 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_101
timestamp 1698175906
transform 1 0 12656 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_107
timestamp 1698175906
transform 1 0 13328 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_117
timestamp 1698175906
transform 1 0 14448 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_125
timestamp 1698175906
transform 1 0 15344 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_129
timestamp 1698175906
transform 1 0 15792 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_136
timestamp 1698175906
transform 1 0 16576 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_144
timestamp 1698175906
transform 1 0 17472 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_148
timestamp 1698175906
transform 1 0 17920 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_150
timestamp 1698175906
transform 1 0 18144 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_156
timestamp 1698175906
transform 1 0 18816 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_166
timestamp 1698175906
transform 1 0 19936 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_174
timestamp 1698175906
transform 1 0 20832 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_177
timestamp 1698175906
transform 1 0 21168 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_185
timestamp 1698175906
transform 1 0 22064 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_189
timestamp 1698175906
transform 1 0 22512 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_220
timestamp 1698175906
transform 1 0 25984 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_224
timestamp 1698175906
transform 1 0 26432 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_240
timestamp 1698175906
transform 1 0 28224 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_244
timestamp 1698175906
transform 1 0 28672 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_247
timestamp 1698175906
transform 1 0 29008 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_311
timestamp 1698175906
transform 1 0 36176 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_317
timestamp 1698175906
transform 1 0 36848 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_2
timestamp 1698175906
transform 1 0 1568 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_66
timestamp 1698175906
transform 1 0 8736 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_72
timestamp 1698175906
transform 1 0 9408 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_80
timestamp 1698175906
transform 1 0 10304 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_84
timestamp 1698175906
transform 1 0 10752 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_123
timestamp 1698175906
transform 1 0 15120 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_127
timestamp 1698175906
transform 1 0 15568 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_135
timestamp 1698175906
transform 1 0 16464 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_139
timestamp 1698175906
transform 1 0 16912 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_142
timestamp 1698175906
transform 1 0 17248 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_144
timestamp 1698175906
transform 1 0 17472 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_176
timestamp 1698175906
transform 1 0 21056 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_192
timestamp 1698175906
transform 1 0 22848 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_194
timestamp 1698175906
transform 1 0 23072 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_209
timestamp 1698175906
transform 1 0 24752 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_212
timestamp 1698175906
transform 1 0 25088 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_276
timestamp 1698175906
transform 1 0 32256 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_282
timestamp 1698175906
transform 1 0 32928 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_346
timestamp 1698175906
transform 1 0 40096 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_348
timestamp 1698175906
transform 1 0 40320 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_28
timestamp 1698175906
transform 1 0 4480 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_32
timestamp 1698175906
transform 1 0 4928 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698175906
transform 1 0 5152 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_37
timestamp 1698175906
transform 1 0 5488 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_101
timestamp 1698175906
transform 1 0 12656 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_107
timestamp 1698175906
transform 1 0 13328 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_111
timestamp 1698175906
transform 1 0 13776 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_119
timestamp 1698175906
transform 1 0 14672 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_135
timestamp 1698175906
transform 1 0 16464 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_139
timestamp 1698175906
transform 1 0 16912 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_141
timestamp 1698175906
transform 1 0 17136 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_148
timestamp 1698175906
transform 1 0 17920 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_156
timestamp 1698175906
transform 1 0 18816 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_189
timestamp 1698175906
transform 1 0 22512 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_193
timestamp 1698175906
transform 1 0 22960 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_223
timestamp 1698175906
transform 1 0 26320 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_227
timestamp 1698175906
transform 1 0 26768 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_243
timestamp 1698175906
transform 1 0 28560 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_247
timestamp 1698175906
transform 1 0 29008 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_311
timestamp 1698175906
transform 1 0 36176 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_317
timestamp 1698175906
transform 1 0 36848 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_28
timestamp 1698175906
transform 1 0 4480 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_60
timestamp 1698175906
transform 1 0 8064 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_68
timestamp 1698175906
transform 1 0 8960 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_72
timestamp 1698175906
transform 1 0 9408 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_88
timestamp 1698175906
transform 1 0 11200 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_96
timestamp 1698175906
transform 1 0 12096 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_104
timestamp 1698175906
transform 1 0 12992 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_108
timestamp 1698175906
transform 1 0 13440 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_138
timestamp 1698175906
transform 1 0 16800 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_142
timestamp 1698175906
transform 1 0 17248 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_146
timestamp 1698175906
transform 1 0 17696 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_154
timestamp 1698175906
transform 1 0 18592 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_156
timestamp 1698175906
transform 1 0 18816 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_165
timestamp 1698175906
transform 1 0 19824 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_181
timestamp 1698175906
transform 1 0 21616 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_197
timestamp 1698175906
transform 1 0 23408 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_206
timestamp 1698175906
transform 1 0 24416 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_212
timestamp 1698175906
transform 1 0 25088 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_228
timestamp 1698175906
transform 1 0 26880 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_240
timestamp 1698175906
transform 1 0 28224 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_272
timestamp 1698175906
transform 1 0 31808 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_282
timestamp 1698175906
transform 1 0 32928 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_314
timestamp 1698175906
transform 1 0 36512 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_322
timestamp 1698175906
transform 1 0 37408 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_28
timestamp 1698175906
transform 1 0 4480 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_32
timestamp 1698175906
transform 1 0 4928 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698175906
transform 1 0 5152 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_37
timestamp 1698175906
transform 1 0 5488 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_69
timestamp 1698175906
transform 1 0 9072 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_73
timestamp 1698175906
transform 1 0 9520 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_113
timestamp 1698175906
transform 1 0 14000 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_117
timestamp 1698175906
transform 1 0 14448 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_177
timestamp 1698175906
transform 1 0 21168 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_181
timestamp 1698175906
transform 1 0 21616 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_188
timestamp 1698175906
transform 1 0 22400 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_196
timestamp 1698175906
transform 1 0 23296 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_200
timestamp 1698175906
transform 1 0 23744 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_210
timestamp 1698175906
transform 1 0 24864 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_247
timestamp 1698175906
transform 1 0 29008 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_311
timestamp 1698175906
transform 1 0 36176 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_317
timestamp 1698175906
transform 1 0 36848 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_28
timestamp 1698175906
transform 1 0 4480 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_60
timestamp 1698175906
transform 1 0 8064 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_68
timestamp 1698175906
transform 1 0 8960 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_72
timestamp 1698175906
transform 1 0 9408 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_88
timestamp 1698175906
transform 1 0 11200 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_96
timestamp 1698175906
transform 1 0 12096 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_104
timestamp 1698175906
transform 1 0 12992 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_107
timestamp 1698175906
transform 1 0 13328 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_129
timestamp 1698175906
transform 1 0 15792 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_142
timestamp 1698175906
transform 1 0 17248 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_150
timestamp 1698175906
transform 1 0 18144 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_154
timestamp 1698175906
transform 1 0 18592 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_185
timestamp 1698175906
transform 1 0 22064 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_196
timestamp 1698175906
transform 1 0 23296 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_198
timestamp 1698175906
transform 1 0 23520 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_212
timestamp 1698175906
transform 1 0 25088 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_245
timestamp 1698175906
transform 1 0 28784 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_277
timestamp 1698175906
transform 1 0 32368 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_279
timestamp 1698175906
transform 1 0 32592 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_282
timestamp 1698175906
transform 1 0 32928 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_314
timestamp 1698175906
transform 1 0 36512 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_322
timestamp 1698175906
transform 1 0 37408 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_28
timestamp 1698175906
transform 1 0 4480 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_32
timestamp 1698175906
transform 1 0 4928 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698175906
transform 1 0 5152 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_37
timestamp 1698175906
transform 1 0 5488 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_101
timestamp 1698175906
transform 1 0 12656 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_107
timestamp 1698175906
transform 1 0 13328 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_115
timestamp 1698175906
transform 1 0 14224 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_117
timestamp 1698175906
transform 1 0 14448 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_124
timestamp 1698175906
transform 1 0 15232 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_132
timestamp 1698175906
transform 1 0 16128 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_136
timestamp 1698175906
transform 1 0 16576 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_146
timestamp 1698175906
transform 1 0 17696 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_177
timestamp 1698175906
transform 1 0 21168 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_179
timestamp 1698175906
transform 1 0 21392 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_230
timestamp 1698175906
transform 1 0 27104 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_238
timestamp 1698175906
transform 1 0 28000 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_242
timestamp 1698175906
transform 1 0 28448 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_244
timestamp 1698175906
transform 1 0 28672 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_247
timestamp 1698175906
transform 1 0 29008 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_311
timestamp 1698175906
transform 1 0 36176 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_317
timestamp 1698175906
transform 1 0 36848 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_2
timestamp 1698175906
transform 1 0 1568 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_66
timestamp 1698175906
transform 1 0 8736 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_72
timestamp 1698175906
transform 1 0 9408 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_104
timestamp 1698175906
transform 1 0 12992 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_107
timestamp 1698175906
transform 1 0 13328 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_111
timestamp 1698175906
transform 1 0 13776 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_137
timestamp 1698175906
transform 1 0 16688 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_139
timestamp 1698175906
transform 1 0 16912 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_142
timestamp 1698175906
transform 1 0 17248 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_146
timestamp 1698175906
transform 1 0 17696 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_209
timestamp 1698175906
transform 1 0 24752 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_225
timestamp 1698175906
transform 1 0 26544 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_257
timestamp 1698175906
transform 1 0 30128 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_273
timestamp 1698175906
transform 1 0 31920 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_277
timestamp 1698175906
transform 1 0 32368 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_279
timestamp 1698175906
transform 1 0 32592 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_282
timestamp 1698175906
transform 1 0 32928 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_314
timestamp 1698175906
transform 1 0 36512 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_322
timestamp 1698175906
transform 1 0 37408 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_2
timestamp 1698175906
transform 1 0 1568 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698175906
transform 1 0 5152 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_37
timestamp 1698175906
transform 1 0 5488 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_69
timestamp 1698175906
transform 1 0 9072 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_73
timestamp 1698175906
transform 1 0 9520 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_75
timestamp 1698175906
transform 1 0 9744 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_107
timestamp 1698175906
transform 1 0 13328 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_114
timestamp 1698175906
transform 1 0 14112 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_118
timestamp 1698175906
transform 1 0 14560 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_126
timestamp 1698175906
transform 1 0 15456 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_128
timestamp 1698175906
transform 1 0 15680 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_146
timestamp 1698175906
transform 1 0 17696 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_173
timestamp 1698175906
transform 1 0 20720 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_185
timestamp 1698175906
transform 1 0 22064 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_187
timestamp 1698175906
transform 1 0 22288 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_229
timestamp 1698175906
transform 1 0 26992 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_247
timestamp 1698175906
transform 1 0 29008 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_311
timestamp 1698175906
transform 1 0 36176 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_317
timestamp 1698175906
transform 1 0 36848 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_2
timestamp 1698175906
transform 1 0 1568 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_66
timestamp 1698175906
transform 1 0 8736 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_72
timestamp 1698175906
transform 1 0 9408 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_80
timestamp 1698175906
transform 1 0 10304 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_125
timestamp 1698175906
transform 1 0 15344 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_129
timestamp 1698175906
transform 1 0 15792 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_131
timestamp 1698175906
transform 1 0 16016 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_138
timestamp 1698175906
transform 1 0 16800 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_142
timestamp 1698175906
transform 1 0 17248 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_159
timestamp 1698175906
transform 1 0 19152 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_172
timestamp 1698175906
transform 1 0 20608 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_176
timestamp 1698175906
transform 1 0 21056 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_183
timestamp 1698175906
transform 1 0 21840 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_191
timestamp 1698175906
transform 1 0 22736 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_198
timestamp 1698175906
transform 1 0 23520 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_212
timestamp 1698175906
transform 1 0 25088 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_216
timestamp 1698175906
transform 1 0 25536 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_247
timestamp 1698175906
transform 1 0 29008 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_279
timestamp 1698175906
transform 1 0 32592 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_282
timestamp 1698175906
transform 1 0 32928 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_314
timestamp 1698175906
transform 1 0 36512 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_322
timestamp 1698175906
transform 1 0 37408 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_2
timestamp 1698175906
transform 1 0 1568 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698175906
transform 1 0 5152 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_37
timestamp 1698175906
transform 1 0 5488 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_101
timestamp 1698175906
transform 1 0 12656 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_107
timestamp 1698175906
transform 1 0 13328 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_114
timestamp 1698175906
transform 1 0 14112 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_146
timestamp 1698175906
transform 1 0 17696 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_160
timestamp 1698175906
transform 1 0 19264 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_167
timestamp 1698175906
transform 1 0 20048 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_174
timestamp 1698175906
transform 1 0 20832 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_177
timestamp 1698175906
transform 1 0 21168 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_193
timestamp 1698175906
transform 1 0 22960 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_195
timestamp 1698175906
transform 1 0 23184 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_202
timestamp 1698175906
transform 1 0 23968 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_206
timestamp 1698175906
transform 1 0 24416 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_247
timestamp 1698175906
transform 1 0 29008 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_311
timestamp 1698175906
transform 1 0 36176 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_317
timestamp 1698175906
transform 1 0 36848 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_321
timestamp 1698175906
transform 1 0 37296 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_2
timestamp 1698175906
transform 1 0 1568 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_66
timestamp 1698175906
transform 1 0 8736 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_72
timestamp 1698175906
transform 1 0 9408 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_104
timestamp 1698175906
transform 1 0 12992 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_120
timestamp 1698175906
transform 1 0 14784 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_122
timestamp 1698175906
transform 1 0 15008 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_129
timestamp 1698175906
transform 1 0 15792 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_139
timestamp 1698175906
transform 1 0 16912 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_150
timestamp 1698175906
transform 1 0 18144 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_154
timestamp 1698175906
transform 1 0 18592 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_156
timestamp 1698175906
transform 1 0 18816 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_161
timestamp 1698175906
transform 1 0 19376 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_177
timestamp 1698175906
transform 1 0 21168 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_185
timestamp 1698175906
transform 1 0 22064 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_192
timestamp 1698175906
transform 1 0 22848 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_208
timestamp 1698175906
transform 1 0 24640 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_212
timestamp 1698175906
transform 1 0 25088 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_218
timestamp 1698175906
transform 1 0 25760 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_250
timestamp 1698175906
transform 1 0 29344 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_266
timestamp 1698175906
transform 1 0 31136 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_274
timestamp 1698175906
transform 1 0 32032 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_278
timestamp 1698175906
transform 1 0 32480 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_282
timestamp 1698175906
transform 1 0 32928 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_346
timestamp 1698175906
transform 1 0 40096 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_348
timestamp 1698175906
transform 1 0 40320 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_2
timestamp 1698175906
transform 1 0 1568 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698175906
transform 1 0 5152 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_37
timestamp 1698175906
transform 1 0 5488 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_101
timestamp 1698175906
transform 1 0 12656 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_107
timestamp 1698175906
transform 1 0 13328 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_137
timestamp 1698175906
transform 1 0 16688 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_149
timestamp 1698175906
transform 1 0 18032 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_157
timestamp 1698175906
transform 1 0 18928 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_171
timestamp 1698175906
transform 1 0 20496 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_177
timestamp 1698175906
transform 1 0 21168 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_181
timestamp 1698175906
transform 1 0 21616 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_197
timestamp 1698175906
transform 1 0 23408 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_205
timestamp 1698175906
transform 1 0 24304 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_207
timestamp 1698175906
transform 1 0 24528 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_217
timestamp 1698175906
transform 1 0 25648 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_233
timestamp 1698175906
transform 1 0 27440 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_241
timestamp 1698175906
transform 1 0 28336 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_247
timestamp 1698175906
transform 1 0 29008 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_311
timestamp 1698175906
transform 1 0 36176 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_317
timestamp 1698175906
transform 1 0 36848 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_2
timestamp 1698175906
transform 1 0 1568 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_66
timestamp 1698175906
transform 1 0 8736 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_72
timestamp 1698175906
transform 1 0 9408 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_88
timestamp 1698175906
transform 1 0 11200 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_96
timestamp 1698175906
transform 1 0 12096 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_129
timestamp 1698175906
transform 1 0 15792 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_135
timestamp 1698175906
transform 1 0 16464 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_139
timestamp 1698175906
transform 1 0 16912 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_142
timestamp 1698175906
transform 1 0 17248 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_150
timestamp 1698175906
transform 1 0 18144 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_154
timestamp 1698175906
transform 1 0 18592 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_179
timestamp 1698175906
transform 1 0 21392 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_187
timestamp 1698175906
transform 1 0 22288 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_209
timestamp 1698175906
transform 1 0 24752 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_212
timestamp 1698175906
transform 1 0 25088 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_216
timestamp 1698175906
transform 1 0 25536 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_228
timestamp 1698175906
transform 1 0 26880 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_238
timestamp 1698175906
transform 1 0 28000 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_270
timestamp 1698175906
transform 1 0 31584 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_278
timestamp 1698175906
transform 1 0 32480 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_282
timestamp 1698175906
transform 1 0 32928 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_314
timestamp 1698175906
transform 1 0 36512 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_322
timestamp 1698175906
transform 1 0 37408 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_28
timestamp 1698175906
transform 1 0 4480 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_32
timestamp 1698175906
transform 1 0 4928 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698175906
transform 1 0 5152 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_37
timestamp 1698175906
transform 1 0 5488 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_101
timestamp 1698175906
transform 1 0 12656 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_107
timestamp 1698175906
transform 1 0 13328 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_115
timestamp 1698175906
transform 1 0 14224 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_125
timestamp 1698175906
transform 1 0 15344 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_131
timestamp 1698175906
transform 1 0 16016 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_135
timestamp 1698175906
transform 1 0 16464 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_137
timestamp 1698175906
transform 1 0 16688 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_185
timestamp 1698175906
transform 1 0 22064 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_247
timestamp 1698175906
transform 1 0 29008 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_311
timestamp 1698175906
transform 1 0 36176 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_317
timestamp 1698175906
transform 1 0 36848 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_321
timestamp 1698175906
transform 1 0 37296 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_2
timestamp 1698175906
transform 1 0 1568 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_66
timestamp 1698175906
transform 1 0 8736 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_72
timestamp 1698175906
transform 1 0 9408 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_136
timestamp 1698175906
transform 1 0 16576 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_142
timestamp 1698175906
transform 1 0 17248 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_150
timestamp 1698175906
transform 1 0 18144 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_180
timestamp 1698175906
transform 1 0 21504 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_184
timestamp 1698175906
transform 1 0 21952 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_200
timestamp 1698175906
transform 1 0 23744 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_208
timestamp 1698175906
transform 1 0 24640 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_212
timestamp 1698175906
transform 1 0 25088 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_218
timestamp 1698175906
transform 1 0 25760 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_250
timestamp 1698175906
transform 1 0 29344 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_266
timestamp 1698175906
transform 1 0 31136 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_274
timestamp 1698175906
transform 1 0 32032 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_278
timestamp 1698175906
transform 1 0 32480 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_282
timestamp 1698175906
transform 1 0 32928 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_346
timestamp 1698175906
transform 1 0 40096 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_348
timestamp 1698175906
transform 1 0 40320 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_2
timestamp 1698175906
transform 1 0 1568 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698175906
transform 1 0 5152 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_37
timestamp 1698175906
transform 1 0 5488 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_101
timestamp 1698175906
transform 1 0 12656 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_107
timestamp 1698175906
transform 1 0 13328 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_139
timestamp 1698175906
transform 1 0 16912 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_155
timestamp 1698175906
transform 1 0 18704 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_163
timestamp 1698175906
transform 1 0 19600 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_169
timestamp 1698175906
transform 1 0 20272 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_173
timestamp 1698175906
transform 1 0 20720 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_177
timestamp 1698175906
transform 1 0 21168 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_241
timestamp 1698175906
transform 1 0 28336 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_247
timestamp 1698175906
transform 1 0 29008 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_311
timestamp 1698175906
transform 1 0 36176 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_317
timestamp 1698175906
transform 1 0 36848 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_2
timestamp 1698175906
transform 1 0 1568 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_66
timestamp 1698175906
transform 1 0 8736 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_72
timestamp 1698175906
transform 1 0 9408 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_136
timestamp 1698175906
transform 1 0 16576 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_142
timestamp 1698175906
transform 1 0 17248 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_206
timestamp 1698175906
transform 1 0 24416 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_212
timestamp 1698175906
transform 1 0 25088 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_276
timestamp 1698175906
transform 1 0 32256 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_282
timestamp 1698175906
transform 1 0 32928 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_346
timestamp 1698175906
transform 1 0 40096 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_348
timestamp 1698175906
transform 1 0 40320 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698175906
transform 1 0 1568 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698175906
transform 1 0 5152 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_37
timestamp 1698175906
transform 1 0 5488 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_101
timestamp 1698175906
transform 1 0 12656 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_107
timestamp 1698175906
transform 1 0 13328 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_171
timestamp 1698175906
transform 1 0 20496 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_177
timestamp 1698175906
transform 1 0 21168 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_241
timestamp 1698175906
transform 1 0 28336 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_247
timestamp 1698175906
transform 1 0 29008 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_311
timestamp 1698175906
transform 1 0 36176 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_317
timestamp 1698175906
transform 1 0 36848 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2
timestamp 1698175906
transform 1 0 1568 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_66
timestamp 1698175906
transform 1 0 8736 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_72
timestamp 1698175906
transform 1 0 9408 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_136
timestamp 1698175906
transform 1 0 16576 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_142
timestamp 1698175906
transform 1 0 17248 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_206
timestamp 1698175906
transform 1 0 24416 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_212
timestamp 1698175906
transform 1 0 25088 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_276
timestamp 1698175906
transform 1 0 32256 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_282
timestamp 1698175906
transform 1 0 32928 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_346
timestamp 1698175906
transform 1 0 40096 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_348
timestamp 1698175906
transform 1 0 40320 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_2
timestamp 1698175906
transform 1 0 1568 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698175906
transform 1 0 5152 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_37
timestamp 1698175906
transform 1 0 5488 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_101
timestamp 1698175906
transform 1 0 12656 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_107
timestamp 1698175906
transform 1 0 13328 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_171
timestamp 1698175906
transform 1 0 20496 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_177
timestamp 1698175906
transform 1 0 21168 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_241
timestamp 1698175906
transform 1 0 28336 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_247
timestamp 1698175906
transform 1 0 29008 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_311
timestamp 1698175906
transform 1 0 36176 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_317
timestamp 1698175906
transform 1 0 36848 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2
timestamp 1698175906
transform 1 0 1568 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_66
timestamp 1698175906
transform 1 0 8736 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_72
timestamp 1698175906
transform 1 0 9408 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_136
timestamp 1698175906
transform 1 0 16576 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_142
timestamp 1698175906
transform 1 0 17248 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_206
timestamp 1698175906
transform 1 0 24416 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_212
timestamp 1698175906
transform 1 0 25088 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_276
timestamp 1698175906
transform 1 0 32256 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_282
timestamp 1698175906
transform 1 0 32928 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_346
timestamp 1698175906
transform 1 0 40096 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_348
timestamp 1698175906
transform 1 0 40320 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698175906
transform 1 0 1568 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698175906
transform 1 0 5152 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_37
timestamp 1698175906
transform 1 0 5488 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_101
timestamp 1698175906
transform 1 0 12656 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_107
timestamp 1698175906
transform 1 0 13328 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_171
timestamp 1698175906
transform 1 0 20496 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_177
timestamp 1698175906
transform 1 0 21168 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_241
timestamp 1698175906
transform 1 0 28336 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_247
timestamp 1698175906
transform 1 0 29008 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_311
timestamp 1698175906
transform 1 0 36176 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_317
timestamp 1698175906
transform 1 0 36848 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_2
timestamp 1698175906
transform 1 0 1568 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_66
timestamp 1698175906
transform 1 0 8736 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_72
timestamp 1698175906
transform 1 0 9408 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_136
timestamp 1698175906
transform 1 0 16576 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_142
timestamp 1698175906
transform 1 0 17248 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_206
timestamp 1698175906
transform 1 0 24416 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_212
timestamp 1698175906
transform 1 0 25088 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_276
timestamp 1698175906
transform 1 0 32256 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_282
timestamp 1698175906
transform 1 0 32928 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_346
timestamp 1698175906
transform 1 0 40096 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_348
timestamp 1698175906
transform 1 0 40320 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698175906
transform 1 0 1568 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698175906
transform 1 0 5152 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_37
timestamp 1698175906
transform 1 0 5488 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_101
timestamp 1698175906
transform 1 0 12656 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_107
timestamp 1698175906
transform 1 0 13328 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_171
timestamp 1698175906
transform 1 0 20496 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_177
timestamp 1698175906
transform 1 0 21168 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_241
timestamp 1698175906
transform 1 0 28336 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_247
timestamp 1698175906
transform 1 0 29008 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_311
timestamp 1698175906
transform 1 0 36176 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_317
timestamp 1698175906
transform 1 0 36848 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2
timestamp 1698175906
transform 1 0 1568 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1698175906
transform 1 0 8736 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_72
timestamp 1698175906
transform 1 0 9408 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_136
timestamp 1698175906
transform 1 0 16576 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_142
timestamp 1698175906
transform 1 0 17248 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_206
timestamp 1698175906
transform 1 0 24416 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_212
timestamp 1698175906
transform 1 0 25088 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_276
timestamp 1698175906
transform 1 0 32256 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_282
timestamp 1698175906
transform 1 0 32928 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_346
timestamp 1698175906
transform 1 0 40096 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_348
timestamp 1698175906
transform 1 0 40320 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_2
timestamp 1698175906
transform 1 0 1568 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698175906
transform 1 0 5152 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_37
timestamp 1698175906
transform 1 0 5488 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_101
timestamp 1698175906
transform 1 0 12656 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_107
timestamp 1698175906
transform 1 0 13328 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_171
timestamp 1698175906
transform 1 0 20496 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_177
timestamp 1698175906
transform 1 0 21168 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_241
timestamp 1698175906
transform 1 0 28336 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_247
timestamp 1698175906
transform 1 0 29008 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_311
timestamp 1698175906
transform 1 0 36176 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_317
timestamp 1698175906
transform 1 0 36848 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_2
timestamp 1698175906
transform 1 0 1568 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_66
timestamp 1698175906
transform 1 0 8736 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_72
timestamp 1698175906
transform 1 0 9408 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_136
timestamp 1698175906
transform 1 0 16576 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_142
timestamp 1698175906
transform 1 0 17248 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_158
timestamp 1698175906
transform 1 0 19040 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_162
timestamp 1698175906
transform 1 0 19488 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_189
timestamp 1698175906
transform 1 0 22512 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_205
timestamp 1698175906
transform 1 0 24304 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_209
timestamp 1698175906
transform 1 0 24752 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_212
timestamp 1698175906
transform 1 0 25088 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_276
timestamp 1698175906
transform 1 0 32256 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_282
timestamp 1698175906
transform 1 0 32928 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_346
timestamp 1698175906
transform 1 0 40096 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_348
timestamp 1698175906
transform 1 0 40320 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_2
timestamp 1698175906
transform 1 0 1568 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_36
timestamp 1698175906
transform 1 0 5376 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_70
timestamp 1698175906
transform 1 0 9184 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_104
timestamp 1698175906
transform 1 0 12992 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_138
timestamp 1698175906
transform 1 0 16800 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_172
timestamp 1698175906
transform 1 0 20608 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_174
timestamp 1698175906
transform 1 0 20832 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_201
timestamp 1698175906
transform 1 0 23856 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_203
timestamp 1698175906
transform 1 0 24080 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_206
timestamp 1698175906
transform 1 0 24416 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_210
timestamp 1698175906
transform 1 0 24864 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_237
timestamp 1698175906
transform 1 0 27888 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_240
timestamp 1698175906
transform 1 0 28224 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_244
timestamp 1698175906
transform 1 0 28672 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_246
timestamp 1698175906
transform 1 0 28896 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_251
timestamp 1698175906
transform 1 0 29456 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_267
timestamp 1698175906
transform 1 0 31248 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_271
timestamp 1698175906
transform 1 0 31696 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_274
timestamp 1698175906
transform 1 0 32032 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_308
timestamp 1698175906
transform 1 0 35840 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_342
timestamp 1698175906
transform 1 0 39648 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_346
timestamp 1698175906
transform 1 0 40096 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_348
timestamp 1698175906
transform 1 0 40320 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita40_25 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 29456 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita40_26
timestamp 1698175906
transform 1 0 39984 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 4480 0 1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output2
timestamp 1698175906
transform 1 0 37520 0 1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output3
timestamp 1698175906
transform 1 0 37520 0 -1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output4
timestamp 1698175906
transform 1 0 24976 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output5
timestamp 1698175906
transform 1 0 23632 0 1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output6
timestamp 1698175906
transform -1 0 4480 0 1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output7
timestamp 1698175906
transform 1 0 24416 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output8
timestamp 1698175906
transform -1 0 4480 0 1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output9
timestamp 1698175906
transform 1 0 37520 0 -1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output10
timestamp 1698175906
transform 1 0 20944 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output11
timestamp 1698175906
transform 1 0 37520 0 -1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output12
timestamp 1698175906
transform 1 0 37520 0 1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output13
timestamp 1698175906
transform 1 0 25088 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output14
timestamp 1698175906
transform 1 0 19600 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output15
timestamp 1698175906
transform 1 0 16912 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output16
timestamp 1698175906
transform 1 0 37520 0 -1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output17
timestamp 1698175906
transform 1 0 28224 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output18
timestamp 1698175906
transform 1 0 20944 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output19
timestamp 1698175906
transform -1 0 4480 0 1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output20
timestamp 1698175906
transform 1 0 15568 0 1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output21
timestamp 1698175906
transform 1 0 37520 0 -1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output22
timestamp 1698175906
transform 1 0 20272 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output23
timestamp 1698175906
transform -1 0 4480 0 -1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output24
timestamp 1698175906
transform -1 0 4480 0 -1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_45 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698175906
transform -1 0 40656 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_46
timestamp 1698175906
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698175906
transform -1 0 40656 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_47
timestamp 1698175906
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698175906
transform -1 0 40656 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_48
timestamp 1698175906
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698175906
transform -1 0 40656 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_49
timestamp 1698175906
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698175906
transform -1 0 40656 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_50
timestamp 1698175906
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698175906
transform -1 0 40656 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_51
timestamp 1698175906
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698175906
transform -1 0 40656 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_52
timestamp 1698175906
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698175906
transform -1 0 40656 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_53
timestamp 1698175906
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698175906
transform -1 0 40656 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_54
timestamp 1698175906
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698175906
transform -1 0 40656 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_55
timestamp 1698175906
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698175906
transform -1 0 40656 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_56
timestamp 1698175906
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698175906
transform -1 0 40656 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_57
timestamp 1698175906
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698175906
transform -1 0 40656 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_58
timestamp 1698175906
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698175906
transform -1 0 40656 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_59
timestamp 1698175906
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698175906
transform -1 0 40656 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_60
timestamp 1698175906
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698175906
transform -1 0 40656 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_61
timestamp 1698175906
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698175906
transform -1 0 40656 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_62
timestamp 1698175906
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698175906
transform -1 0 40656 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_63
timestamp 1698175906
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698175906
transform -1 0 40656 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_64
timestamp 1698175906
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698175906
transform -1 0 40656 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_65
timestamp 1698175906
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698175906
transform -1 0 40656 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_66
timestamp 1698175906
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698175906
transform -1 0 40656 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_67
timestamp 1698175906
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698175906
transform -1 0 40656 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_68
timestamp 1698175906
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698175906
transform -1 0 40656 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_69
timestamp 1698175906
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698175906
transform -1 0 40656 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_70
timestamp 1698175906
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698175906
transform -1 0 40656 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_71
timestamp 1698175906
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698175906
transform -1 0 40656 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_72
timestamp 1698175906
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698175906
transform -1 0 40656 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_73
timestamp 1698175906
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698175906
transform -1 0 40656 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_74
timestamp 1698175906
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698175906
transform -1 0 40656 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_75
timestamp 1698175906
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698175906
transform -1 0 40656 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_76
timestamp 1698175906
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698175906
transform -1 0 40656 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_77
timestamp 1698175906
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698175906
transform -1 0 40656 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_78
timestamp 1698175906
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698175906
transform -1 0 40656 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_79
timestamp 1698175906
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698175906
transform -1 0 40656 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_80
timestamp 1698175906
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698175906
transform -1 0 40656 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_81
timestamp 1698175906
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698175906
transform -1 0 40656 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_82
timestamp 1698175906
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698175906
transform -1 0 40656 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_83
timestamp 1698175906
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698175906
transform -1 0 40656 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_84
timestamp 1698175906
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698175906
transform -1 0 40656 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_85
timestamp 1698175906
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698175906
transform -1 0 40656 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_86
timestamp 1698175906
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698175906
transform -1 0 40656 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_87
timestamp 1698175906
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698175906
transform -1 0 40656 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_88
timestamp 1698175906
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698175906
transform -1 0 40656 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_89
timestamp 1698175906
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698175906
transform -1 0 40656 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_90 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_91
timestamp 1698175906
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_92
timestamp 1698175906
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_93
timestamp 1698175906
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_94
timestamp 1698175906
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_95
timestamp 1698175906
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_96
timestamp 1698175906
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_97
timestamp 1698175906
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_98
timestamp 1698175906
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_99
timestamp 1698175906
transform 1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_100
timestamp 1698175906
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_101
timestamp 1698175906
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_102
timestamp 1698175906
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_103
timestamp 1698175906
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_104
timestamp 1698175906
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_105
timestamp 1698175906
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_106
timestamp 1698175906
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_107
timestamp 1698175906
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_108
timestamp 1698175906
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_109
timestamp 1698175906
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_110
timestamp 1698175906
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_111
timestamp 1698175906
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_112
timestamp 1698175906
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_113
timestamp 1698175906
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_114
timestamp 1698175906
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_115
timestamp 1698175906
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_116
timestamp 1698175906
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_117
timestamp 1698175906
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_118
timestamp 1698175906
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_119
timestamp 1698175906
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_120
timestamp 1698175906
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_121
timestamp 1698175906
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_122
timestamp 1698175906
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_123
timestamp 1698175906
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_124
timestamp 1698175906
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_125
timestamp 1698175906
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_126
timestamp 1698175906
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_127
timestamp 1698175906
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_128
timestamp 1698175906
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_129
timestamp 1698175906
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_130
timestamp 1698175906
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_131
timestamp 1698175906
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_132
timestamp 1698175906
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_133
timestamp 1698175906
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_134
timestamp 1698175906
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_135
timestamp 1698175906
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_136
timestamp 1698175906
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_137
timestamp 1698175906
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_138
timestamp 1698175906
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_139
timestamp 1698175906
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_140
timestamp 1698175906
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_141
timestamp 1698175906
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_142
timestamp 1698175906
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_143
timestamp 1698175906
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_144
timestamp 1698175906
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_145
timestamp 1698175906
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_146
timestamp 1698175906
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_147
timestamp 1698175906
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_148
timestamp 1698175906
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_149
timestamp 1698175906
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_150
timestamp 1698175906
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_151
timestamp 1698175906
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_152
timestamp 1698175906
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_153
timestamp 1698175906
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_154
timestamp 1698175906
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_155
timestamp 1698175906
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_156
timestamp 1698175906
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_157
timestamp 1698175906
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_158
timestamp 1698175906
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_159
timestamp 1698175906
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_160
timestamp 1698175906
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_161
timestamp 1698175906
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_162
timestamp 1698175906
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_163
timestamp 1698175906
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_164
timestamp 1698175906
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_165
timestamp 1698175906
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_166
timestamp 1698175906
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_167
timestamp 1698175906
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_168
timestamp 1698175906
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_169
timestamp 1698175906
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_170
timestamp 1698175906
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_171
timestamp 1698175906
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_172
timestamp 1698175906
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_173
timestamp 1698175906
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_174
timestamp 1698175906
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_175
timestamp 1698175906
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_176
timestamp 1698175906
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_177
timestamp 1698175906
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_178
timestamp 1698175906
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_179
timestamp 1698175906
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_180
timestamp 1698175906
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_181
timestamp 1698175906
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_182
timestamp 1698175906
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_183
timestamp 1698175906
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_184
timestamp 1698175906
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_185
timestamp 1698175906
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_186
timestamp 1698175906
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_187
timestamp 1698175906
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_188
timestamp 1698175906
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_189
timestamp 1698175906
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_190
timestamp 1698175906
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_191
timestamp 1698175906
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_192
timestamp 1698175906
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_193
timestamp 1698175906
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_194
timestamp 1698175906
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_195
timestamp 1698175906
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_196
timestamp 1698175906
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_197
timestamp 1698175906
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_198
timestamp 1698175906
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_199
timestamp 1698175906
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_200
timestamp 1698175906
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_201
timestamp 1698175906
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_202
timestamp 1698175906
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_203
timestamp 1698175906
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_204
timestamp 1698175906
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_205
timestamp 1698175906
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_206
timestamp 1698175906
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_207
timestamp 1698175906
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_208
timestamp 1698175906
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_209
timestamp 1698175906
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_210
timestamp 1698175906
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_211
timestamp 1698175906
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_212
timestamp 1698175906
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_213
timestamp 1698175906
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_214
timestamp 1698175906
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_215
timestamp 1698175906
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_216
timestamp 1698175906
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_217
timestamp 1698175906
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_218
timestamp 1698175906
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_219
timestamp 1698175906
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_220
timestamp 1698175906
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_221
timestamp 1698175906
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_222
timestamp 1698175906
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_223
timestamp 1698175906
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_224
timestamp 1698175906
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_225
timestamp 1698175906
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_226
timestamp 1698175906
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_227
timestamp 1698175906
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_228
timestamp 1698175906
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_229
timestamp 1698175906
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_230
timestamp 1698175906
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_231
timestamp 1698175906
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_232
timestamp 1698175906
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_233
timestamp 1698175906
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_234
timestamp 1698175906
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_235
timestamp 1698175906
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_236
timestamp 1698175906
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_237
timestamp 1698175906
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_238
timestamp 1698175906
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_239
timestamp 1698175906
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_240
timestamp 1698175906
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_241
timestamp 1698175906
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_242
timestamp 1698175906
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_243
timestamp 1698175906
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_244
timestamp 1698175906
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_245
timestamp 1698175906
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_246
timestamp 1698175906
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_247
timestamp 1698175906
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_248
timestamp 1698175906
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_249
timestamp 1698175906
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_250
timestamp 1698175906
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_251
timestamp 1698175906
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_252
timestamp 1698175906
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_253
timestamp 1698175906
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_254
timestamp 1698175906
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_255
timestamp 1698175906
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_256
timestamp 1698175906
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_257
timestamp 1698175906
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_258
timestamp 1698175906
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_259
timestamp 1698175906
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_260
timestamp 1698175906
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_261
timestamp 1698175906
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_262
timestamp 1698175906
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_263
timestamp 1698175906
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_264
timestamp 1698175906
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_265
timestamp 1698175906
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_266
timestamp 1698175906
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_267
timestamp 1698175906
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_268
timestamp 1698175906
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_269
timestamp 1698175906
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_270
timestamp 1698175906
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_271
timestamp 1698175906
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_272
timestamp 1698175906
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_273
timestamp 1698175906
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_274
timestamp 1698175906
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_275
timestamp 1698175906
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_276
timestamp 1698175906
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_277
timestamp 1698175906
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_278
timestamp 1698175906
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_279
timestamp 1698175906
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_280
timestamp 1698175906
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_281
timestamp 1698175906
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_282
timestamp 1698175906
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_283
timestamp 1698175906
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_284
timestamp 1698175906
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_285
timestamp 1698175906
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_286
timestamp 1698175906
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_287
timestamp 1698175906
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_288
timestamp 1698175906
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_289
timestamp 1698175906
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_290
timestamp 1698175906
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_291
timestamp 1698175906
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_292
timestamp 1698175906
transform 1 0 32704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_293
timestamp 1698175906
transform 1 0 5152 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_294
timestamp 1698175906
transform 1 0 8960 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_295
timestamp 1698175906
transform 1 0 12768 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_296
timestamp 1698175906
transform 1 0 16576 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_297
timestamp 1698175906
transform 1 0 20384 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_298
timestamp 1698175906
transform 1 0 24192 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_299
timestamp 1698175906
transform 1 0 28000 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_300
timestamp 1698175906
transform 1 0 31808 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_301
timestamp 1698175906
transform 1 0 35616 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_302
timestamp 1698175906
transform 1 0 39424 0 1 37632
box -86 -86 310 870
<< labels >>
flabel metal3 s 0 27552 800 27664 0 FreeSans 448 0 0 0 clk
port 0 nsew signal input
flabel metal2 s 28896 41200 29008 42000 0 FreeSans 448 90 0 0 segm[0]
port 1 nsew signal tristate
flabel metal3 s 0 26208 800 26320 0 FreeSans 448 0 0 0 segm[10]
port 2 nsew signal tristate
flabel metal3 s 41200 23520 42000 23632 0 FreeSans 448 0 0 0 segm[11]
port 3 nsew signal tristate
flabel metal3 s 41200 22848 42000 22960 0 FreeSans 448 0 0 0 segm[12]
port 4 nsew signal tristate
flabel metal2 s 24864 41200 24976 42000 0 FreeSans 448 90 0 0 segm[13]
port 5 nsew signal tristate
flabel metal2 s 23520 0 23632 800 0 FreeSans 448 90 0 0 segm[1]
port 6 nsew signal tristate
flabel metal3 s 0 18816 800 18928 0 FreeSans 448 0 0 0 segm[2]
port 7 nsew signal tristate
flabel metal3 s 41200 11424 42000 11536 0 FreeSans 448 0 0 0 segm[3]
port 8 nsew signal tristate
flabel metal2 s 22848 0 22960 800 0 FreeSans 448 90 0 0 segm[4]
port 9 nsew signal tristate
flabel metal3 s 0 20160 800 20272 0 FreeSans 448 0 0 0 segm[5]
port 10 nsew signal tristate
flabel metal3 s 41200 19488 42000 19600 0 FreeSans 448 0 0 0 segm[6]
port 11 nsew signal tristate
flabel metal2 s 20832 41200 20944 42000 0 FreeSans 448 90 0 0 segm[7]
port 12 nsew signal tristate
flabel metal3 s 41200 26880 42000 26992 0 FreeSans 448 0 0 0 segm[8]
port 13 nsew signal tristate
flabel metal3 s 41200 26208 42000 26320 0 FreeSans 448 0 0 0 segm[9]
port 14 nsew signal tristate
flabel metal2 s 24192 0 24304 800 0 FreeSans 448 90 0 0 sel[0]
port 15 nsew signal tristate
flabel metal2 s 19488 41200 19600 42000 0 FreeSans 448 90 0 0 sel[10]
port 16 nsew signal tristate
flabel metal2 s 16800 0 16912 800 0 FreeSans 448 90 0 0 sel[11]
port 17 nsew signal tristate
flabel metal3 s 41200 20832 42000 20944 0 FreeSans 448 0 0 0 sel[1]
port 18 nsew signal tristate
flabel metal2 s 24864 0 24976 800 0 FreeSans 448 90 0 0 sel[2]
port 19 nsew signal tristate
flabel metal2 s 20832 0 20944 800 0 FreeSans 448 90 0 0 sel[3]
port 20 nsew signal tristate
flabel metal3 s 0 16800 800 16912 0 FreeSans 448 0 0 0 sel[4]
port 21 nsew signal tristate
flabel metal2 s 15456 0 15568 800 0 FreeSans 448 90 0 0 sel[5]
port 22 nsew signal tristate
flabel metal3 s 41200 18144 42000 18256 0 FreeSans 448 0 0 0 sel[6]
port 23 nsew signal tristate
flabel metal2 s 20160 0 20272 800 0 FreeSans 448 90 0 0 sel[7]
port 24 nsew signal tristate
flabel metal3 s 0 18144 800 18256 0 FreeSans 448 0 0 0 sel[8]
port 25 nsew signal tristate
flabel metal3 s 0 19488 800 19600 0 FreeSans 448 0 0 0 sel[9]
port 26 nsew signal tristate
flabel metal4 s 4448 3076 4768 38476 0 FreeSans 1280 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 35168 3076 35488 38476 0 FreeSans 1280 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 19808 3076 20128 38476 0 FreeSans 1280 90 0 0 vss
port 28 nsew ground bidirectional
rlabel metal1 21000 38416 21000 38416 0 vdd
rlabel metal1 21000 37632 21000 37632 0 vss
rlabel metal2 24472 20776 24472 20776 0 _000_
rlabel metal2 22624 13832 22624 13832 0 _001_
rlabel metal2 12152 19544 12152 19544 0 _002_
rlabel metal3 25872 23800 25872 23800 0 _003_
rlabel metal2 25816 22512 25816 22512 0 _004_
rlabel metal2 26488 19600 26488 19600 0 _005_
rlabel metal2 19040 16184 19040 16184 0 _006_
rlabel metal3 19768 27048 19768 27048 0 _007_
rlabel metal2 14728 14056 14728 14056 0 _008_
rlabel metal2 20608 27160 20608 27160 0 _009_
rlabel metal3 25816 26936 25816 26936 0 _010_
rlabel metal2 14840 26600 14840 26600 0 _011_
rlabel metal2 23128 26936 23128 26936 0 _012_
rlabel metal2 15288 18032 15288 18032 0 _013_
rlabel metal2 14392 24472 14392 24472 0 _014_
rlabel via2 13608 23016 13608 23016 0 _015_
rlabel metal2 10808 22512 10808 22512 0 _016_
rlabel metal2 18760 17024 18760 17024 0 _017_
rlabel metal2 23968 17752 23968 17752 0 _018_
rlabel metal2 14280 14840 14280 14840 0 _019_
rlabel metal2 13272 17192 13272 17192 0 _020_
rlabel metal2 19040 13832 19040 13832 0 _021_
rlabel metal2 23688 16240 23688 16240 0 _022_
rlabel metal2 24024 21224 24024 21224 0 _023_
rlabel metal2 23632 22344 23632 22344 0 _024_
rlabel metal3 22568 22344 22568 22344 0 _025_
rlabel metal2 23016 17584 23016 17584 0 _026_
rlabel metal2 23800 21840 23800 21840 0 _027_
rlabel metal2 22568 15008 22568 15008 0 _028_
rlabel metal3 14952 20104 14952 20104 0 _029_
rlabel metal3 13104 19880 13104 19880 0 _030_
rlabel metal3 21224 24024 21224 24024 0 _031_
rlabel metal2 25144 24640 25144 24640 0 _032_
rlabel metal2 24584 22568 24584 22568 0 _033_
rlabel metal2 26264 22456 26264 22456 0 _034_
rlabel metal2 20328 25144 20328 25144 0 _035_
rlabel metal2 22680 25984 22680 25984 0 _036_
rlabel metal2 22008 26992 22008 26992 0 _037_
rlabel metal3 25032 22344 25032 22344 0 _038_
rlabel metal2 24696 22176 24696 22176 0 _039_
rlabel metal2 24808 18928 24808 18928 0 _040_
rlabel metal2 24248 20720 24248 20720 0 _041_
rlabel metal2 20328 15736 20328 15736 0 _042_
rlabel metal3 20048 25368 20048 25368 0 _043_
rlabel metal3 20608 26264 20608 26264 0 _044_
rlabel metal2 19768 25928 19768 25928 0 _045_
rlabel metal3 20832 26936 20832 26936 0 _046_
rlabel metal2 17360 13944 17360 13944 0 _047_
rlabel metal3 20552 26712 20552 26712 0 _048_
rlabel metal2 25032 25760 25032 25760 0 _049_
rlabel metal2 14728 26768 14728 26768 0 _050_
rlabel metal2 22680 20832 22680 20832 0 _051_
rlabel metal2 26040 21896 26040 21896 0 _052_
rlabel metal2 14616 26656 14616 26656 0 _053_
rlabel metal2 14952 26264 14952 26264 0 _054_
rlabel metal2 13944 24304 13944 24304 0 _055_
rlabel metal2 15288 26936 15288 26936 0 _056_
rlabel metal3 23688 26264 23688 26264 0 _057_
rlabel metal2 22792 25088 22792 25088 0 _058_
rlabel metal2 23184 25592 23184 25592 0 _059_
rlabel metal2 20664 18144 20664 18144 0 _060_
rlabel metal3 21112 15512 21112 15512 0 _061_
rlabel metal2 15064 16464 15064 16464 0 _062_
rlabel metal2 19824 23128 19824 23128 0 _063_
rlabel metal2 19656 20384 19656 20384 0 _064_
rlabel metal2 19880 24192 19880 24192 0 _065_
rlabel metal2 17416 24976 17416 24976 0 _066_
rlabel metal2 18200 23576 18200 23576 0 _067_
rlabel metal2 18424 23576 18424 23576 0 _068_
rlabel metal2 16856 19936 16856 19936 0 _069_
rlabel metal2 15512 17864 15512 17864 0 _070_
rlabel metal2 14840 22736 14840 22736 0 _071_
rlabel metal3 17024 22120 17024 22120 0 _072_
rlabel metal2 13944 22680 13944 22680 0 _073_
rlabel metal3 19824 22904 19824 22904 0 _074_
rlabel metal2 18368 20552 18368 20552 0 _075_
rlabel metal2 20552 20048 20552 20048 0 _076_
rlabel metal2 21392 22232 21392 22232 0 _077_
rlabel metal2 19432 22008 19432 22008 0 _078_
rlabel metal2 19152 23128 19152 23128 0 _079_
rlabel metal3 18872 15064 18872 15064 0 _080_
rlabel metal3 16576 15176 16576 15176 0 _081_
rlabel metal2 18536 16968 18536 16968 0 _082_
rlabel metal2 23128 22736 23128 22736 0 _083_
rlabel metal2 19656 17696 19656 17696 0 _084_
rlabel metal2 24024 20440 24024 20440 0 _085_
rlabel metal2 22456 25032 22456 25032 0 _086_
rlabel metal3 21504 15288 21504 15288 0 _087_
rlabel metal2 14168 21952 14168 21952 0 _088_
rlabel metal2 23688 23128 23688 23128 0 _089_
rlabel metal2 24584 19376 24584 19376 0 _090_
rlabel metal2 24304 18536 24304 18536 0 _091_
rlabel metal2 15848 16352 15848 16352 0 _092_
rlabel metal3 14840 15176 14840 15176 0 _093_
rlabel metal2 13944 19488 13944 19488 0 _094_
rlabel metal2 14280 18424 14280 18424 0 _095_
rlabel metal3 21672 14616 21672 14616 0 _096_
rlabel metal2 14504 17304 14504 17304 0 _097_
rlabel metal2 20216 13552 20216 13552 0 _098_
rlabel metal2 14728 19880 14728 19880 0 _099_
rlabel metal3 23968 16744 23968 16744 0 _100_
rlabel metal2 23352 22512 23352 22512 0 _101_
rlabel metal2 22792 21728 22792 21728 0 _102_
rlabel metal3 2478 27608 2478 27608 0 clk
rlabel metal2 21672 21112 21672 21112 0 clknet_0_clk
rlabel metal2 10920 22736 10920 22736 0 clknet_1_0__leaf_clk
rlabel metal2 21616 27832 21616 27832 0 clknet_1_1__leaf_clk
rlabel metal2 16520 25536 16520 25536 0 dut40.count\[0\]
rlabel metal3 14168 23016 14168 23016 0 dut40.count\[1\]
rlabel metal2 14392 21616 14392 21616 0 dut40.count\[2\]
rlabel metal3 20440 17640 20440 17640 0 dut40.count\[3\]
rlabel metal2 12712 26600 12712 26600 0 net1
rlabel metal2 20720 26936 20720 26936 0 net10
rlabel metal3 29876 26376 29876 26376 0 net11
rlabel metal2 27608 26376 27608 26376 0 net12
rlabel metal3 24864 14280 24864 14280 0 net13
rlabel metal2 19880 27608 19880 27608 0 net14
rlabel metal2 17080 5964 17080 5964 0 net15
rlabel metal2 28616 20720 28616 20720 0 net16
rlabel metal2 28616 9856 28616 9856 0 net17
rlabel metal2 21056 13608 21056 13608 0 net18
rlabel metal2 11144 17192 11144 17192 0 net19
rlabel metal2 28616 23184 28616 23184 0 net2
rlabel metal2 15736 6748 15736 6748 0 net20
rlabel metal2 37688 18088 37688 18088 0 net21
rlabel metal2 20440 6356 20440 6356 0 net22
rlabel metal3 6356 18424 6356 18424 0 net23
rlabel metal2 12488 19320 12488 19320 0 net24
rlabel metal2 29064 37912 29064 37912 0 net25
rlabel metal2 40264 11872 40264 11872 0 net26
rlabel metal2 28840 23072 28840 23072 0 net3
rlabel metal2 25368 32592 25368 32592 0 net4
rlabel metal2 23800 6748 23800 6748 0 net5
rlabel metal2 13496 19152 13496 19152 0 net6
rlabel metal2 24584 5964 24584 5964 0 net7
rlabel metal2 4200 20048 4200 20048 0 net8
rlabel metal2 28056 18872 28056 18872 0 net9
rlabel metal3 1358 26264 1358 26264 0 segm[10]
rlabel metal2 40040 23800 40040 23800 0 segm[11]
rlabel metal3 40642 22904 40642 22904 0 segm[12]
rlabel metal2 24920 39746 24920 39746 0 segm[13]
rlabel metal2 23576 2982 23576 2982 0 segm[1]
rlabel metal3 1358 18872 1358 18872 0 segm[2]
rlabel metal2 22904 2086 22904 2086 0 segm[4]
rlabel metal3 1358 20216 1358 20216 0 segm[5]
rlabel metal2 40040 19656 40040 19656 0 segm[6]
rlabel metal2 20888 39746 20888 39746 0 segm[7]
rlabel metal2 39928 26488 39928 26488 0 segm[8]
rlabel metal2 40040 26712 40040 26712 0 segm[9]
rlabel metal2 24248 2422 24248 2422 0 sel[0]
rlabel metal2 19544 39354 19544 39354 0 sel[10]
rlabel metal2 16856 2086 16856 2086 0 sel[11]
rlabel metal2 40040 21112 40040 21112 0 sel[1]
rlabel metal2 24920 2198 24920 2198 0 sel[2]
rlabel metal2 20888 2198 20888 2198 0 sel[3]
rlabel metal3 1358 16856 1358 16856 0 sel[4]
rlabel metal2 15512 2982 15512 2982 0 sel[5]
rlabel metal3 40642 18200 40642 18200 0 sel[6]
rlabel metal2 20216 2422 20216 2422 0 sel[7]
rlabel metal3 1358 18200 1358 18200 0 sel[8]
rlabel metal3 1358 19544 1358 19544 0 sel[9]
<< properties >>
string FIXED_BBOX 0 0 42000 42000
<< end >>
