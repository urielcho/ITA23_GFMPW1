magic
tech gf180mcuD
magscale 1 10
timestamp 1699642131
<< metal1 >>
rect 1344 38442 40656 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 40656 38442
rect 1344 38356 40656 38390
rect 25566 38274 25618 38286
rect 25566 38210 25618 38222
rect 18162 38110 18174 38162
rect 18226 38110 18238 38162
rect 22194 38110 22206 38162
rect 22258 38110 22270 38162
rect 19730 37998 19742 38050
rect 19794 37998 19806 38050
rect 23762 37998 23774 38050
rect 23826 37998 23838 38050
rect 24546 37998 24558 38050
rect 24610 37998 24622 38050
rect 1344 37658 40656 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 40656 37658
rect 1344 37572 40656 37606
rect 22094 37490 22146 37502
rect 22094 37426 22146 37438
rect 21074 37214 21086 37266
rect 21138 37214 21150 37266
rect 1344 36874 40656 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 40656 36874
rect 1344 36788 40656 36822
rect 1344 36090 40656 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 40656 36090
rect 1344 36004 40656 36038
rect 1344 35306 40656 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 40656 35306
rect 1344 35220 40656 35254
rect 1344 34522 40656 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 40656 34522
rect 1344 34436 40656 34470
rect 1344 33738 40656 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 40656 33738
rect 1344 33652 40656 33686
rect 1344 32954 40656 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 40656 32954
rect 1344 32868 40656 32902
rect 1344 32170 40656 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 40656 32170
rect 1344 32084 40656 32118
rect 1344 31386 40656 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 40656 31386
rect 1344 31300 40656 31334
rect 1344 30602 40656 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 40656 30602
rect 1344 30516 40656 30550
rect 1344 29818 40656 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 40656 29818
rect 1344 29732 40656 29766
rect 1344 29034 40656 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 40656 29034
rect 1344 28948 40656 28982
rect 20738 28702 20750 28754
rect 20802 28702 20814 28754
rect 17826 28590 17838 28642
rect 17890 28590 17902 28642
rect 18610 28478 18622 28530
rect 18674 28478 18686 28530
rect 21422 28418 21474 28430
rect 21422 28354 21474 28366
rect 1344 28250 40656 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 40656 28250
rect 1344 28164 40656 28198
rect 19182 28082 19234 28094
rect 19182 28018 19234 28030
rect 20078 28082 20130 28094
rect 20078 28018 20130 28030
rect 23774 28082 23826 28094
rect 24098 28030 24110 28082
rect 24162 28030 24174 28082
rect 23774 28018 23826 28030
rect 19854 27970 19906 27982
rect 19854 27906 19906 27918
rect 19070 27858 19122 27870
rect 14354 27806 14366 27858
rect 14418 27806 14430 27858
rect 19070 27794 19122 27806
rect 19294 27858 19346 27870
rect 19294 27794 19346 27806
rect 19742 27858 19794 27870
rect 19742 27794 19794 27806
rect 20190 27858 20242 27870
rect 24670 27858 24722 27870
rect 20626 27806 20638 27858
rect 20690 27806 20702 27858
rect 20190 27794 20242 27806
rect 24670 27794 24722 27806
rect 14814 27746 14866 27758
rect 11442 27694 11454 27746
rect 11506 27694 11518 27746
rect 13570 27694 13582 27746
rect 13634 27694 13646 27746
rect 21298 27694 21310 27746
rect 21362 27694 21374 27746
rect 23426 27694 23438 27746
rect 23490 27694 23502 27746
rect 14814 27682 14866 27694
rect 1344 27466 40656 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 40656 27466
rect 1344 27380 40656 27414
rect 13918 27298 13970 27310
rect 13918 27234 13970 27246
rect 22318 27298 22370 27310
rect 22318 27234 22370 27246
rect 1934 27186 1986 27198
rect 21422 27186 21474 27198
rect 19842 27134 19854 27186
rect 19906 27134 19918 27186
rect 1934 27122 1986 27134
rect 21422 27122 21474 27134
rect 40238 27186 40290 27198
rect 40238 27122 40290 27134
rect 20190 27074 20242 27086
rect 4274 27022 4286 27074
rect 4338 27022 4350 27074
rect 17042 27022 17054 27074
rect 17106 27022 17118 27074
rect 20190 27010 20242 27022
rect 20750 27074 20802 27086
rect 20750 27010 20802 27022
rect 21982 27074 22034 27086
rect 21982 27010 22034 27022
rect 22206 27074 22258 27086
rect 22206 27010 22258 27022
rect 13470 26962 13522 26974
rect 13470 26898 13522 26910
rect 14030 26962 14082 26974
rect 21310 26962 21362 26974
rect 17714 26910 17726 26962
rect 17778 26910 17790 26962
rect 14030 26898 14082 26910
rect 21310 26898 21362 26910
rect 22318 26962 22370 26974
rect 22318 26898 22370 26910
rect 13582 26850 13634 26862
rect 13582 26786 13634 26798
rect 14926 26850 14978 26862
rect 14926 26786 14978 26798
rect 21534 26850 21586 26862
rect 21534 26786 21586 26798
rect 1344 26682 40656 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 40656 26682
rect 1344 26596 40656 26630
rect 15374 26514 15426 26526
rect 15374 26450 15426 26462
rect 18734 26514 18786 26526
rect 18734 26450 18786 26462
rect 21086 26514 21138 26526
rect 21086 26450 21138 26462
rect 13906 26350 13918 26402
rect 13970 26350 13982 26402
rect 15262 26290 15314 26302
rect 4274 26238 4286 26290
rect 4338 26238 4350 26290
rect 14690 26238 14702 26290
rect 14754 26238 14766 26290
rect 15026 26238 15038 26290
rect 15090 26238 15102 26290
rect 15262 26226 15314 26238
rect 15486 26290 15538 26302
rect 18622 26290 18674 26302
rect 20638 26290 20690 26302
rect 15698 26238 15710 26290
rect 15762 26238 15774 26290
rect 20178 26238 20190 26290
rect 20242 26238 20254 26290
rect 15486 26226 15538 26238
rect 18622 26226 18674 26238
rect 20638 26226 20690 26238
rect 2034 26126 2046 26178
rect 2098 26126 2110 26178
rect 11778 26126 11790 26178
rect 11842 26126 11854 26178
rect 1344 25898 40656 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 40656 25898
rect 1344 25812 40656 25846
rect 14254 25618 14306 25630
rect 19742 25618 19794 25630
rect 18274 25566 18286 25618
rect 18338 25566 18350 25618
rect 14254 25554 14306 25566
rect 19742 25554 19794 25566
rect 14030 25506 14082 25518
rect 14030 25442 14082 25454
rect 14366 25506 14418 25518
rect 19070 25506 19122 25518
rect 14578 25454 14590 25506
rect 14642 25454 14654 25506
rect 15474 25454 15486 25506
rect 15538 25454 15550 25506
rect 21410 25454 21422 25506
rect 21474 25454 21486 25506
rect 14366 25442 14418 25454
rect 19070 25442 19122 25454
rect 18622 25394 18674 25406
rect 16146 25342 16158 25394
rect 16210 25342 16222 25394
rect 21634 25342 21646 25394
rect 21698 25342 21710 25394
rect 18622 25330 18674 25342
rect 14142 25282 14194 25294
rect 14142 25218 14194 25230
rect 18846 25282 18898 25294
rect 18846 25218 18898 25230
rect 18958 25282 19010 25294
rect 18958 25218 19010 25230
rect 19182 25282 19234 25294
rect 19182 25218 19234 25230
rect 1344 25114 40656 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 40656 25114
rect 1344 25028 40656 25062
rect 17502 24946 17554 24958
rect 17502 24882 17554 24894
rect 17950 24834 18002 24846
rect 18274 24782 18286 24834
rect 18338 24782 18350 24834
rect 17950 24770 18002 24782
rect 17390 24722 17442 24734
rect 17390 24658 17442 24670
rect 17614 24722 17666 24734
rect 25342 24722 25394 24734
rect 18498 24670 18510 24722
rect 18562 24670 18574 24722
rect 24658 24670 24670 24722
rect 24722 24670 24734 24722
rect 37874 24670 37886 24722
rect 37938 24670 37950 24722
rect 17614 24658 17666 24670
rect 25342 24658 25394 24670
rect 21746 24558 21758 24610
rect 21810 24558 21822 24610
rect 23874 24558 23886 24610
rect 23938 24558 23950 24610
rect 40014 24498 40066 24510
rect 40014 24434 40066 24446
rect 1344 24330 40656 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 40656 24330
rect 1344 24244 40656 24278
rect 13470 24162 13522 24174
rect 13470 24098 13522 24110
rect 28142 24162 28194 24174
rect 28142 24098 28194 24110
rect 14254 24050 14306 24062
rect 14254 23986 14306 23998
rect 15374 24050 15426 24062
rect 21422 24050 21474 24062
rect 18834 23998 18846 24050
rect 18898 23998 18910 24050
rect 15374 23986 15426 23998
rect 21422 23986 21474 23998
rect 22654 24050 22706 24062
rect 40014 24050 40066 24062
rect 26338 23998 26350 24050
rect 26402 23998 26414 24050
rect 22654 23986 22706 23998
rect 40014 23986 40066 23998
rect 22542 23938 22594 23950
rect 13794 23886 13806 23938
rect 13858 23886 13870 23938
rect 18610 23886 18622 23938
rect 18674 23886 18686 23938
rect 21634 23886 21646 23938
rect 21698 23886 21710 23938
rect 22542 23874 22594 23886
rect 23214 23938 23266 23950
rect 27358 23938 27410 23950
rect 23538 23886 23550 23938
rect 23602 23886 23614 23938
rect 37650 23886 37662 23938
rect 37714 23886 37726 23938
rect 23214 23874 23266 23886
rect 27358 23874 27410 23886
rect 17726 23826 17778 23838
rect 19854 23826 19906 23838
rect 18050 23774 18062 23826
rect 18114 23774 18126 23826
rect 17726 23762 17778 23774
rect 19854 23762 19906 23774
rect 21310 23826 21362 23838
rect 28030 23826 28082 23838
rect 24210 23774 24222 23826
rect 24274 23774 24286 23826
rect 21310 23762 21362 23774
rect 28030 23762 28082 23774
rect 13582 23714 13634 23726
rect 13582 23650 13634 23662
rect 14142 23714 14194 23726
rect 14142 23650 14194 23662
rect 18510 23714 18562 23726
rect 18510 23650 18562 23662
rect 19742 23714 19794 23726
rect 19742 23650 19794 23662
rect 22766 23714 22818 23726
rect 22766 23650 22818 23662
rect 26686 23714 26738 23726
rect 28142 23714 28194 23726
rect 27010 23662 27022 23714
rect 27074 23662 27086 23714
rect 27682 23662 27694 23714
rect 27746 23662 27758 23714
rect 26686 23650 26738 23662
rect 28142 23650 28194 23662
rect 1344 23546 40656 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 40656 23546
rect 1344 23460 40656 23494
rect 18734 23378 18786 23390
rect 23550 23378 23602 23390
rect 22530 23326 22542 23378
rect 22594 23326 22606 23378
rect 18734 23314 18786 23326
rect 23550 23314 23602 23326
rect 23662 23378 23714 23390
rect 23662 23314 23714 23326
rect 26574 23378 26626 23390
rect 26574 23314 26626 23326
rect 18510 23266 18562 23278
rect 13010 23214 13022 23266
rect 13074 23214 13086 23266
rect 27682 23214 27694 23266
rect 27746 23214 27758 23266
rect 18510 23202 18562 23214
rect 15822 23154 15874 23166
rect 18398 23154 18450 23166
rect 12226 23102 12238 23154
rect 12290 23102 12302 23154
rect 17602 23102 17614 23154
rect 17666 23102 17678 23154
rect 15822 23090 15874 23102
rect 18398 23090 18450 23102
rect 19294 23154 19346 23166
rect 19294 23090 19346 23102
rect 19518 23154 19570 23166
rect 19518 23090 19570 23102
rect 19854 23154 19906 23166
rect 22206 23154 22258 23166
rect 20402 23102 20414 23154
rect 20466 23102 20478 23154
rect 21746 23102 21758 23154
rect 21810 23102 21822 23154
rect 19854 23090 19906 23102
rect 22206 23090 22258 23102
rect 22878 23154 22930 23166
rect 22878 23090 22930 23102
rect 22990 23154 23042 23166
rect 22990 23090 23042 23102
rect 23774 23154 23826 23166
rect 23774 23090 23826 23102
rect 24222 23154 24274 23166
rect 30270 23154 30322 23166
rect 26898 23102 26910 23154
rect 26962 23102 26974 23154
rect 37650 23102 37662 23154
rect 37714 23102 37726 23154
rect 24222 23090 24274 23102
rect 30270 23090 30322 23102
rect 16382 23042 16434 23054
rect 15138 22990 15150 23042
rect 15202 22990 15214 23042
rect 16382 22978 16434 22990
rect 18062 23042 18114 23054
rect 20178 22990 20190 23042
rect 20242 22990 20254 23042
rect 21410 22990 21422 23042
rect 21474 22990 21486 23042
rect 29810 22990 29822 23042
rect 29874 22990 29886 23042
rect 18062 22978 18114 22990
rect 40014 22930 40066 22942
rect 18946 22878 18958 22930
rect 19010 22878 19022 22930
rect 40014 22866 40066 22878
rect 1344 22762 40656 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 40656 22762
rect 1344 22676 40656 22710
rect 19394 22542 19406 22594
rect 19458 22542 19470 22594
rect 28142 22482 28194 22494
rect 24210 22430 24222 22482
rect 24274 22430 24286 22482
rect 28142 22418 28194 22430
rect 28590 22482 28642 22494
rect 28590 22418 28642 22430
rect 40014 22482 40066 22494
rect 40014 22418 40066 22430
rect 13470 22370 13522 22382
rect 13470 22306 13522 22318
rect 13806 22370 13858 22382
rect 16046 22370 16098 22382
rect 21310 22370 21362 22382
rect 15586 22318 15598 22370
rect 15650 22318 15662 22370
rect 16706 22318 16718 22370
rect 16770 22318 16782 22370
rect 17602 22318 17614 22370
rect 17666 22318 17678 22370
rect 18722 22318 18734 22370
rect 18786 22318 18798 22370
rect 19170 22318 19182 22370
rect 19234 22318 19246 22370
rect 19618 22318 19630 22370
rect 19682 22318 19694 22370
rect 20514 22318 20526 22370
rect 20578 22318 20590 22370
rect 13806 22306 13858 22318
rect 16046 22306 16098 22318
rect 21310 22306 21362 22318
rect 21758 22370 21810 22382
rect 21758 22306 21810 22318
rect 22430 22370 22482 22382
rect 22430 22306 22482 22318
rect 22990 22370 23042 22382
rect 22990 22306 23042 22318
rect 23662 22370 23714 22382
rect 23662 22306 23714 22318
rect 29038 22370 29090 22382
rect 29038 22306 29090 22318
rect 29374 22370 29426 22382
rect 37874 22318 37886 22370
rect 37938 22318 37950 22370
rect 29374 22306 29426 22318
rect 14030 22258 14082 22270
rect 22094 22258 22146 22270
rect 16482 22206 16494 22258
rect 16546 22206 16558 22258
rect 18274 22206 18286 22258
rect 18338 22206 18350 22258
rect 19282 22206 19294 22258
rect 19346 22206 19358 22258
rect 14030 22194 14082 22206
rect 22094 22194 22146 22206
rect 24222 22258 24274 22270
rect 24222 22194 24274 22206
rect 29262 22258 29314 22270
rect 29262 22194 29314 22206
rect 13582 22146 13634 22158
rect 23998 22146 24050 22158
rect 17714 22094 17726 22146
rect 17778 22094 17790 22146
rect 13582 22082 13634 22094
rect 23998 22082 24050 22094
rect 1344 21978 40656 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 40656 21978
rect 1344 21892 40656 21926
rect 17726 21810 17778 21822
rect 17378 21758 17390 21810
rect 17442 21758 17454 21810
rect 17726 21746 17778 21758
rect 12338 21646 12350 21698
rect 12402 21646 12414 21698
rect 16382 21586 16434 21598
rect 4274 21534 4286 21586
rect 4338 21534 4350 21586
rect 11554 21534 11566 21586
rect 11618 21534 11630 21586
rect 16258 21534 16270 21586
rect 16322 21534 16334 21586
rect 16382 21522 16434 21534
rect 18510 21586 18562 21598
rect 19394 21534 19406 21586
rect 19458 21534 19470 21586
rect 25330 21534 25342 21586
rect 25394 21534 25406 21586
rect 28578 21534 28590 21586
rect 28642 21534 28654 21586
rect 37650 21534 37662 21586
rect 37714 21534 37726 21586
rect 18510 21522 18562 21534
rect 14926 21474 14978 21486
rect 18734 21474 18786 21486
rect 14466 21422 14478 21474
rect 14530 21422 14542 21474
rect 16146 21422 16158 21474
rect 16210 21422 16222 21474
rect 23314 21422 23326 21474
rect 23378 21422 23390 21474
rect 26002 21422 26014 21474
rect 26066 21422 26078 21474
rect 28130 21422 28142 21474
rect 28194 21422 28206 21474
rect 29250 21422 29262 21474
rect 29314 21422 29326 21474
rect 31378 21422 31390 21474
rect 31442 21422 31454 21474
rect 39890 21422 39902 21474
rect 39954 21422 39966 21474
rect 14926 21410 14978 21422
rect 18734 21410 18786 21422
rect 1934 21362 1986 21374
rect 18174 21362 18226 21374
rect 15698 21310 15710 21362
rect 15762 21310 15774 21362
rect 1934 21298 1986 21310
rect 18174 21298 18226 21310
rect 1344 21194 40656 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 40656 21194
rect 1344 21108 40656 21142
rect 17838 21026 17890 21038
rect 21858 20974 21870 21026
rect 21922 20974 21934 21026
rect 17838 20962 17890 20974
rect 13582 20914 13634 20926
rect 19294 20914 19346 20926
rect 20526 20914 20578 20926
rect 29598 20914 29650 20926
rect 9986 20862 9998 20914
rect 10050 20862 10062 20914
rect 14242 20862 14254 20914
rect 14306 20862 14318 20914
rect 19730 20862 19742 20914
rect 19794 20862 19806 20914
rect 25330 20862 25342 20914
rect 25394 20862 25406 20914
rect 13582 20850 13634 20862
rect 19294 20850 19346 20862
rect 20526 20850 20578 20862
rect 29598 20850 29650 20862
rect 40014 20914 40066 20926
rect 40014 20850 40066 20862
rect 15822 20802 15874 20814
rect 12114 20750 12126 20802
rect 12178 20750 12190 20802
rect 12786 20750 12798 20802
rect 12850 20750 12862 20802
rect 14130 20750 14142 20802
rect 14194 20750 14206 20802
rect 14802 20750 14814 20802
rect 14866 20750 14878 20802
rect 15822 20738 15874 20750
rect 16830 20802 16882 20814
rect 16830 20738 16882 20750
rect 18062 20802 18114 20814
rect 18062 20738 18114 20750
rect 18622 20802 18674 20814
rect 18622 20738 18674 20750
rect 19070 20802 19122 20814
rect 29486 20802 29538 20814
rect 19842 20750 19854 20802
rect 19906 20750 19918 20802
rect 21522 20750 21534 20802
rect 21586 20750 21598 20802
rect 21858 20750 21870 20802
rect 21922 20750 21934 20802
rect 23314 20750 23326 20802
rect 23378 20750 23390 20802
rect 19070 20738 19122 20750
rect 29486 20738 29538 20750
rect 29710 20802 29762 20814
rect 29710 20738 29762 20750
rect 30046 20802 30098 20814
rect 30046 20738 30098 20750
rect 30606 20802 30658 20814
rect 37650 20750 37662 20802
rect 37714 20750 37726 20802
rect 30606 20738 30658 20750
rect 15374 20690 15426 20702
rect 15374 20626 15426 20638
rect 21310 20690 21362 20702
rect 29150 20690 29202 20702
rect 22754 20638 22766 20690
rect 22818 20638 22830 20690
rect 21310 20626 21362 20638
rect 29150 20626 29202 20638
rect 30158 20690 30210 20702
rect 30158 20626 30210 20638
rect 30718 20690 30770 20702
rect 30718 20626 30770 20638
rect 14366 20578 14418 20590
rect 14366 20514 14418 20526
rect 14590 20578 14642 20590
rect 14590 20514 14642 20526
rect 15150 20578 15202 20590
rect 15150 20514 15202 20526
rect 15262 20578 15314 20590
rect 18398 20578 18450 20590
rect 17154 20526 17166 20578
rect 17218 20526 17230 20578
rect 17490 20526 17502 20578
rect 17554 20526 17566 20578
rect 15262 20514 15314 20526
rect 18398 20514 18450 20526
rect 18510 20578 18562 20590
rect 22430 20578 22482 20590
rect 21746 20526 21758 20578
rect 21810 20526 21822 20578
rect 18510 20514 18562 20526
rect 22430 20514 22482 20526
rect 30382 20578 30434 20590
rect 30382 20514 30434 20526
rect 1344 20410 40656 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 40656 20410
rect 1344 20324 40656 20358
rect 24558 20242 24610 20254
rect 24558 20178 24610 20190
rect 23102 20130 23154 20142
rect 15698 20078 15710 20130
rect 15762 20078 15774 20130
rect 19394 20078 19406 20130
rect 19458 20078 19470 20130
rect 23102 20066 23154 20078
rect 23326 20130 23378 20142
rect 23326 20066 23378 20078
rect 24334 20130 24386 20142
rect 24334 20066 24386 20078
rect 24446 20130 24498 20142
rect 24446 20066 24498 20078
rect 24670 20130 24722 20142
rect 24670 20066 24722 20078
rect 25230 20130 25282 20142
rect 25230 20066 25282 20078
rect 26238 20130 26290 20142
rect 26238 20066 26290 20078
rect 26686 20130 26738 20142
rect 26686 20066 26738 20078
rect 26798 20130 26850 20142
rect 26798 20066 26850 20078
rect 22990 20018 23042 20030
rect 25566 20018 25618 20030
rect 15474 19966 15486 20018
rect 15538 19966 15550 20018
rect 22530 19966 22542 20018
rect 22594 19966 22606 20018
rect 23874 19966 23886 20018
rect 23938 19966 23950 20018
rect 22990 19954 23042 19966
rect 25566 19954 25618 19966
rect 25678 20018 25730 20030
rect 25678 19954 25730 19966
rect 26126 20018 26178 20030
rect 26126 19954 26178 19966
rect 26462 20018 26514 20030
rect 27682 19966 27694 20018
rect 27746 19966 27758 20018
rect 37650 19966 37662 20018
rect 37714 19966 37726 20018
rect 26462 19954 26514 19966
rect 14142 19906 14194 19918
rect 14142 19842 14194 19854
rect 25342 19906 25394 19918
rect 25342 19842 25394 19854
rect 27358 19906 27410 19918
rect 28466 19854 28478 19906
rect 28530 19854 28542 19906
rect 30594 19854 30606 19906
rect 30658 19854 30670 19906
rect 27358 19842 27410 19854
rect 40014 19794 40066 19806
rect 40014 19730 40066 19742
rect 1344 19626 40656 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 40656 19626
rect 1344 19540 40656 19574
rect 28366 19458 28418 19470
rect 28366 19394 28418 19406
rect 1934 19346 1986 19358
rect 21746 19294 21758 19346
rect 21810 19294 21822 19346
rect 27234 19294 27246 19346
rect 27298 19294 27310 19346
rect 1934 19282 1986 19294
rect 13470 19234 13522 19246
rect 4274 19182 4286 19234
rect 4338 19182 4350 19234
rect 13470 19170 13522 19182
rect 13806 19234 13858 19246
rect 13806 19170 13858 19182
rect 14814 19234 14866 19246
rect 16942 19234 16994 19246
rect 18846 19234 18898 19246
rect 15026 19182 15038 19234
rect 15090 19182 15102 19234
rect 16258 19182 16270 19234
rect 16322 19182 16334 19234
rect 18274 19182 18286 19234
rect 18338 19182 18350 19234
rect 14814 19170 14866 19182
rect 16942 19170 16994 19182
rect 18846 19170 18898 19182
rect 20302 19234 20354 19246
rect 20302 19170 20354 19182
rect 21198 19234 21250 19246
rect 28478 19234 28530 19246
rect 21522 19182 21534 19234
rect 21586 19182 21598 19234
rect 24322 19182 24334 19234
rect 24386 19182 24398 19234
rect 21198 19170 21250 19182
rect 28478 19170 28530 19182
rect 14030 19122 14082 19134
rect 14030 19058 14082 19070
rect 14366 19122 14418 19134
rect 14366 19058 14418 19070
rect 14702 19122 14754 19134
rect 14702 19058 14754 19070
rect 15934 19122 15986 19134
rect 19966 19122 20018 19134
rect 16594 19070 16606 19122
rect 16658 19070 16670 19122
rect 18498 19070 18510 19122
rect 18562 19070 18574 19122
rect 15934 19058 15986 19070
rect 19966 19058 20018 19070
rect 21758 19122 21810 19134
rect 21758 19058 21810 19070
rect 22430 19122 22482 19134
rect 25106 19070 25118 19122
rect 25170 19070 25182 19122
rect 22430 19058 22482 19070
rect 13582 19010 13634 19022
rect 13582 18946 13634 18958
rect 14590 19010 14642 19022
rect 14590 18946 14642 18958
rect 16046 19010 16098 19022
rect 27694 19010 27746 19022
rect 19170 18958 19182 19010
rect 19234 18958 19246 19010
rect 22082 18958 22094 19010
rect 22146 18958 22158 19010
rect 16046 18946 16098 18958
rect 27694 18946 27746 18958
rect 28366 19010 28418 19022
rect 28366 18946 28418 18958
rect 1344 18842 40656 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 40656 18842
rect 1344 18756 40656 18790
rect 17502 18674 17554 18686
rect 23426 18622 23438 18674
rect 23490 18622 23502 18674
rect 17502 18610 17554 18622
rect 14366 18562 14418 18574
rect 14366 18498 14418 18510
rect 15486 18562 15538 18574
rect 15486 18498 15538 18510
rect 15822 18562 15874 18574
rect 15822 18498 15874 18510
rect 17614 18562 17666 18574
rect 17614 18498 17666 18510
rect 18622 18562 18674 18574
rect 18622 18498 18674 18510
rect 19518 18562 19570 18574
rect 19518 18498 19570 18510
rect 20526 18562 20578 18574
rect 20526 18498 20578 18510
rect 22542 18562 22594 18574
rect 22542 18498 22594 18510
rect 25342 18562 25394 18574
rect 25342 18498 25394 18510
rect 25566 18562 25618 18574
rect 25566 18498 25618 18510
rect 14590 18450 14642 18462
rect 4274 18398 4286 18450
rect 4338 18398 4350 18450
rect 13122 18398 13134 18450
rect 13186 18398 13198 18450
rect 13906 18398 13918 18450
rect 13970 18398 13982 18450
rect 14590 18386 14642 18398
rect 14814 18450 14866 18462
rect 14814 18386 14866 18398
rect 15038 18450 15090 18462
rect 15038 18386 15090 18398
rect 15262 18450 15314 18462
rect 15262 18386 15314 18398
rect 16606 18450 16658 18462
rect 16606 18386 16658 18398
rect 17278 18450 17330 18462
rect 17278 18386 17330 18398
rect 18062 18450 18114 18462
rect 18062 18386 18114 18398
rect 18286 18450 18338 18462
rect 18286 18386 18338 18398
rect 19070 18450 19122 18462
rect 19070 18386 19122 18398
rect 19182 18450 19234 18462
rect 19182 18386 19234 18398
rect 19406 18450 19458 18462
rect 19842 18398 19854 18450
rect 19906 18398 19918 18450
rect 22082 18398 22094 18450
rect 22146 18398 22158 18450
rect 19406 18386 19458 18398
rect 15710 18338 15762 18350
rect 10994 18286 11006 18338
rect 11058 18286 11070 18338
rect 15710 18274 15762 18286
rect 18174 18338 18226 18350
rect 25218 18286 25230 18338
rect 25282 18286 25294 18338
rect 18174 18274 18226 18286
rect 1934 18226 1986 18238
rect 1934 18162 1986 18174
rect 1344 18058 40656 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 40656 18058
rect 1344 17972 40656 18006
rect 22990 17890 23042 17902
rect 22990 17826 23042 17838
rect 23662 17890 23714 17902
rect 23662 17826 23714 17838
rect 21646 17778 21698 17790
rect 13458 17726 13470 17778
rect 13522 17726 13534 17778
rect 15586 17726 15598 17778
rect 15650 17726 15662 17778
rect 21646 17714 21698 17726
rect 22766 17778 22818 17790
rect 40014 17778 40066 17790
rect 27906 17726 27918 17778
rect 27970 17726 27982 17778
rect 22766 17714 22818 17726
rect 40014 17714 40066 17726
rect 16830 17666 16882 17678
rect 16258 17614 16270 17666
rect 16322 17614 16334 17666
rect 16830 17602 16882 17614
rect 16942 17666 16994 17678
rect 16942 17602 16994 17614
rect 17166 17666 17218 17678
rect 17166 17602 17218 17614
rect 17950 17666 18002 17678
rect 21870 17666 21922 17678
rect 19618 17614 19630 17666
rect 19682 17614 19694 17666
rect 20178 17614 20190 17666
rect 20242 17614 20254 17666
rect 20738 17614 20750 17666
rect 20802 17614 20814 17666
rect 17950 17602 18002 17614
rect 21870 17602 21922 17614
rect 22430 17666 22482 17678
rect 22430 17602 22482 17614
rect 23774 17666 23826 17678
rect 27806 17666 27858 17678
rect 23986 17614 23998 17666
rect 24050 17614 24062 17666
rect 23774 17602 23826 17614
rect 27806 17602 27858 17614
rect 29150 17666 29202 17678
rect 37650 17614 37662 17666
rect 37714 17614 37726 17666
rect 29150 17602 29202 17614
rect 17614 17554 17666 17566
rect 21422 17554 21474 17566
rect 27358 17554 27410 17566
rect 19394 17502 19406 17554
rect 19458 17502 19470 17554
rect 19954 17502 19966 17554
rect 20018 17502 20030 17554
rect 22082 17502 22094 17554
rect 22146 17502 22158 17554
rect 17614 17490 17666 17502
rect 21422 17490 21474 17502
rect 27358 17490 27410 17502
rect 27582 17554 27634 17566
rect 27582 17490 27634 17502
rect 27918 17554 27970 17566
rect 27918 17490 27970 17502
rect 29262 17554 29314 17566
rect 29262 17490 29314 17502
rect 17054 17442 17106 17454
rect 17054 17378 17106 17390
rect 17278 17442 17330 17454
rect 17278 17378 17330 17390
rect 17838 17442 17890 17454
rect 21970 17390 21982 17442
rect 22034 17390 22046 17442
rect 23314 17390 23326 17442
rect 23378 17390 23390 17442
rect 17838 17378 17890 17390
rect 1344 17274 40656 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 40656 17274
rect 1344 17188 40656 17222
rect 17502 17106 17554 17118
rect 17502 17042 17554 17054
rect 18734 17106 18786 17118
rect 18734 17042 18786 17054
rect 14690 16942 14702 16994
rect 14754 16942 14766 16994
rect 22082 16942 22094 16994
rect 22146 16942 22158 16994
rect 28018 16942 28030 16994
rect 28082 16942 28094 16994
rect 24670 16882 24722 16894
rect 14018 16830 14030 16882
rect 14082 16830 14094 16882
rect 20290 16830 20302 16882
rect 20354 16830 20366 16882
rect 21410 16830 21422 16882
rect 21474 16830 21486 16882
rect 24670 16818 24722 16830
rect 26910 16882 26962 16894
rect 27234 16830 27246 16882
rect 27298 16830 27310 16882
rect 37650 16830 37662 16882
rect 37714 16830 37726 16882
rect 26910 16818 26962 16830
rect 18846 16770 18898 16782
rect 16818 16718 16830 16770
rect 16882 16718 16894 16770
rect 18846 16706 18898 16718
rect 19070 16770 19122 16782
rect 19070 16706 19122 16718
rect 20078 16770 20130 16782
rect 24210 16718 24222 16770
rect 24274 16718 24286 16770
rect 30146 16718 30158 16770
rect 30210 16718 30222 16770
rect 20078 16706 20130 16718
rect 18734 16658 18786 16670
rect 18734 16594 18786 16606
rect 19294 16658 19346 16670
rect 19294 16594 19346 16606
rect 19742 16658 19794 16670
rect 19742 16594 19794 16606
rect 19854 16658 19906 16670
rect 19854 16594 19906 16606
rect 40014 16658 40066 16670
rect 40014 16594 40066 16606
rect 1344 16490 40656 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 40656 16490
rect 1344 16404 40656 16438
rect 18174 16322 18226 16334
rect 18174 16258 18226 16270
rect 18510 16322 18562 16334
rect 18510 16258 18562 16270
rect 19182 16322 19234 16334
rect 19182 16258 19234 16270
rect 19294 16322 19346 16334
rect 19294 16258 19346 16270
rect 19518 16322 19570 16334
rect 19518 16258 19570 16270
rect 20078 16322 20130 16334
rect 20078 16258 20130 16270
rect 20302 16322 20354 16334
rect 20302 16258 20354 16270
rect 21758 16322 21810 16334
rect 21758 16258 21810 16270
rect 24670 16210 24722 16222
rect 21410 16158 21422 16210
rect 21474 16158 21486 16210
rect 24670 16146 24722 16158
rect 25118 16210 25170 16222
rect 29262 16210 29314 16222
rect 28578 16158 28590 16210
rect 28642 16158 28654 16210
rect 25118 16146 25170 16158
rect 29262 16146 29314 16158
rect 19630 16098 19682 16110
rect 18498 16046 18510 16098
rect 18562 16046 18574 16098
rect 19630 16034 19682 16046
rect 20526 16098 20578 16110
rect 20738 16046 20750 16098
rect 20802 16046 20814 16098
rect 25666 16046 25678 16098
rect 25730 16046 25742 16098
rect 20526 16034 20578 16046
rect 24446 15986 24498 15998
rect 24446 15922 24498 15934
rect 25006 15986 25058 15998
rect 26450 15934 26462 15986
rect 26514 15934 26526 15986
rect 25006 15922 25058 15934
rect 20638 15874 20690 15886
rect 20638 15810 20690 15822
rect 21534 15874 21586 15886
rect 21534 15810 21586 15822
rect 24558 15874 24610 15886
rect 24558 15810 24610 15822
rect 25230 15874 25282 15886
rect 25230 15810 25282 15822
rect 1344 15706 40656 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 40656 15706
rect 1344 15620 40656 15654
rect 26686 15538 26738 15550
rect 26686 15474 26738 15486
rect 17390 15426 17442 15438
rect 17390 15362 17442 15374
rect 17726 15426 17778 15438
rect 20190 15426 20242 15438
rect 18722 15374 18734 15426
rect 18786 15374 18798 15426
rect 17726 15362 17778 15374
rect 20190 15362 20242 15374
rect 20526 15426 20578 15438
rect 20526 15362 20578 15374
rect 26910 15314 26962 15326
rect 18498 15262 18510 15314
rect 18562 15262 18574 15314
rect 26910 15250 26962 15262
rect 27358 15314 27410 15326
rect 27570 15262 27582 15314
rect 27634 15262 27646 15314
rect 27358 15250 27410 15262
rect 26562 15150 26574 15202
rect 26626 15150 26638 15202
rect 27246 15090 27298 15102
rect 27246 15026 27298 15038
rect 1344 14922 40656 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 40656 14922
rect 1344 14836 40656 14870
rect 18946 14702 18958 14754
rect 19010 14751 19022 14754
rect 19282 14751 19294 14754
rect 19010 14705 19294 14751
rect 19010 14702 19022 14705
rect 19282 14702 19294 14705
rect 19346 14702 19358 14754
rect 26910 14642 26962 14654
rect 16594 14590 16606 14642
rect 16658 14590 16670 14642
rect 18722 14590 18734 14642
rect 18786 14590 18798 14642
rect 24210 14590 24222 14642
rect 24274 14590 24286 14642
rect 26338 14590 26350 14642
rect 26402 14590 26414 14642
rect 26910 14578 26962 14590
rect 15922 14478 15934 14530
rect 15986 14478 15998 14530
rect 23538 14478 23550 14530
rect 23602 14478 23614 14530
rect 19182 14306 19234 14318
rect 19182 14242 19234 14254
rect 1344 14138 40656 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 40656 14138
rect 1344 14052 40656 14086
rect 20066 13806 20078 13858
rect 20130 13806 20142 13858
rect 22654 13746 22706 13758
rect 19394 13694 19406 13746
rect 19458 13694 19470 13746
rect 22654 13682 22706 13694
rect 22194 13582 22206 13634
rect 22258 13582 22270 13634
rect 1344 13354 40656 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 40656 13354
rect 1344 13268 40656 13302
rect 1344 12570 40656 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 40656 12570
rect 1344 12484 40656 12518
rect 1344 11786 40656 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 40656 11786
rect 1344 11700 40656 11734
rect 1344 11002 40656 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 40656 11002
rect 1344 10916 40656 10950
rect 1344 10218 40656 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 40656 10218
rect 1344 10132 40656 10166
rect 1344 9434 40656 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 40656 9434
rect 1344 9348 40656 9382
rect 1344 8650 40656 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 40656 8650
rect 1344 8564 40656 8598
rect 1344 7866 40656 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 40656 7866
rect 1344 7780 40656 7814
rect 1344 7082 40656 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 40656 7082
rect 1344 6996 40656 7030
rect 1344 6298 40656 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 40656 6298
rect 1344 6212 40656 6246
rect 1344 5514 40656 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 40656 5514
rect 1344 5428 40656 5462
rect 18734 5234 18786 5246
rect 18734 5170 18786 5182
rect 17714 5070 17726 5122
rect 17778 5070 17790 5122
rect 1344 4730 40656 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 40656 4730
rect 1344 4644 40656 4678
rect 24446 4450 24498 4462
rect 24446 4386 24498 4398
rect 19058 4286 19070 4338
rect 19122 4286 19134 4338
rect 25778 4286 25790 4338
rect 25842 4286 25854 4338
rect 20078 4114 20130 4126
rect 20078 4050 20130 4062
rect 26798 4114 26850 4126
rect 26798 4050 26850 4062
rect 1344 3946 40656 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 40656 3946
rect 1344 3860 40656 3894
rect 25566 3666 25618 3678
rect 18162 3614 18174 3666
rect 18226 3614 18238 3666
rect 25566 3602 25618 3614
rect 19730 3502 19742 3554
rect 19794 3502 19806 3554
rect 21410 3502 21422 3554
rect 21474 3502 21486 3554
rect 24546 3502 24558 3554
rect 24610 3502 24622 3554
rect 22430 3330 22482 3342
rect 22430 3266 22482 3278
rect 1344 3162 40656 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 40656 3162
rect 1344 3076 40656 3110
<< via1 >>
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 25566 38222 25618 38274
rect 18174 38110 18226 38162
rect 22206 38110 22258 38162
rect 19742 37998 19794 38050
rect 23774 37998 23826 38050
rect 24558 37998 24610 38050
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 22094 37438 22146 37490
rect 21086 37214 21138 37266
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 20750 28702 20802 28754
rect 17838 28590 17890 28642
rect 18622 28478 18674 28530
rect 21422 28366 21474 28418
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 19182 28030 19234 28082
rect 20078 28030 20130 28082
rect 23774 28030 23826 28082
rect 24110 28030 24162 28082
rect 19854 27918 19906 27970
rect 14366 27806 14418 27858
rect 19070 27806 19122 27858
rect 19294 27806 19346 27858
rect 19742 27806 19794 27858
rect 20190 27806 20242 27858
rect 20638 27806 20690 27858
rect 24670 27806 24722 27858
rect 11454 27694 11506 27746
rect 13582 27694 13634 27746
rect 14814 27694 14866 27746
rect 21310 27694 21362 27746
rect 23438 27694 23490 27746
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 13918 27246 13970 27298
rect 22318 27246 22370 27298
rect 1934 27134 1986 27186
rect 19854 27134 19906 27186
rect 21422 27134 21474 27186
rect 40238 27134 40290 27186
rect 4286 27022 4338 27074
rect 17054 27022 17106 27074
rect 20190 27022 20242 27074
rect 20750 27022 20802 27074
rect 21982 27022 22034 27074
rect 22206 27022 22258 27074
rect 13470 26910 13522 26962
rect 14030 26910 14082 26962
rect 17726 26910 17778 26962
rect 21310 26910 21362 26962
rect 22318 26910 22370 26962
rect 13582 26798 13634 26850
rect 14926 26798 14978 26850
rect 21534 26798 21586 26850
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 15374 26462 15426 26514
rect 18734 26462 18786 26514
rect 21086 26462 21138 26514
rect 13918 26350 13970 26402
rect 4286 26238 4338 26290
rect 14702 26238 14754 26290
rect 15038 26238 15090 26290
rect 15262 26238 15314 26290
rect 15486 26238 15538 26290
rect 15710 26238 15762 26290
rect 18622 26238 18674 26290
rect 20190 26238 20242 26290
rect 20638 26238 20690 26290
rect 2046 26126 2098 26178
rect 11790 26126 11842 26178
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 14254 25566 14306 25618
rect 18286 25566 18338 25618
rect 19742 25566 19794 25618
rect 14030 25454 14082 25506
rect 14366 25454 14418 25506
rect 14590 25454 14642 25506
rect 15486 25454 15538 25506
rect 19070 25454 19122 25506
rect 21422 25454 21474 25506
rect 16158 25342 16210 25394
rect 18622 25342 18674 25394
rect 21646 25342 21698 25394
rect 14142 25230 14194 25282
rect 18846 25230 18898 25282
rect 18958 25230 19010 25282
rect 19182 25230 19234 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 17502 24894 17554 24946
rect 17950 24782 18002 24834
rect 18286 24782 18338 24834
rect 17390 24670 17442 24722
rect 17614 24670 17666 24722
rect 18510 24670 18562 24722
rect 24670 24670 24722 24722
rect 25342 24670 25394 24722
rect 37886 24670 37938 24722
rect 21758 24558 21810 24610
rect 23886 24558 23938 24610
rect 40014 24446 40066 24498
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 13470 24110 13522 24162
rect 28142 24110 28194 24162
rect 14254 23998 14306 24050
rect 15374 23998 15426 24050
rect 18846 23998 18898 24050
rect 21422 23998 21474 24050
rect 22654 23998 22706 24050
rect 26350 23998 26402 24050
rect 40014 23998 40066 24050
rect 13806 23886 13858 23938
rect 18622 23886 18674 23938
rect 21646 23886 21698 23938
rect 22542 23886 22594 23938
rect 23214 23886 23266 23938
rect 23550 23886 23602 23938
rect 27358 23886 27410 23938
rect 37662 23886 37714 23938
rect 17726 23774 17778 23826
rect 18062 23774 18114 23826
rect 19854 23774 19906 23826
rect 21310 23774 21362 23826
rect 24222 23774 24274 23826
rect 28030 23774 28082 23826
rect 13582 23662 13634 23714
rect 14142 23662 14194 23714
rect 18510 23662 18562 23714
rect 19742 23662 19794 23714
rect 22766 23662 22818 23714
rect 26686 23662 26738 23714
rect 27022 23662 27074 23714
rect 27694 23662 27746 23714
rect 28142 23662 28194 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 18734 23326 18786 23378
rect 22542 23326 22594 23378
rect 23550 23326 23602 23378
rect 23662 23326 23714 23378
rect 26574 23326 26626 23378
rect 13022 23214 13074 23266
rect 18510 23214 18562 23266
rect 27694 23214 27746 23266
rect 12238 23102 12290 23154
rect 15822 23102 15874 23154
rect 17614 23102 17666 23154
rect 18398 23102 18450 23154
rect 19294 23102 19346 23154
rect 19518 23102 19570 23154
rect 19854 23102 19906 23154
rect 20414 23102 20466 23154
rect 21758 23102 21810 23154
rect 22206 23102 22258 23154
rect 22878 23102 22930 23154
rect 22990 23102 23042 23154
rect 23774 23102 23826 23154
rect 24222 23102 24274 23154
rect 26910 23102 26962 23154
rect 30270 23102 30322 23154
rect 37662 23102 37714 23154
rect 15150 22990 15202 23042
rect 16382 22990 16434 23042
rect 18062 22990 18114 23042
rect 20190 22990 20242 23042
rect 21422 22990 21474 23042
rect 29822 22990 29874 23042
rect 18958 22878 19010 22930
rect 40014 22878 40066 22930
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 19406 22542 19458 22594
rect 24222 22430 24274 22482
rect 28142 22430 28194 22482
rect 28590 22430 28642 22482
rect 40014 22430 40066 22482
rect 13470 22318 13522 22370
rect 13806 22318 13858 22370
rect 15598 22318 15650 22370
rect 16046 22318 16098 22370
rect 16718 22318 16770 22370
rect 17614 22318 17666 22370
rect 18734 22318 18786 22370
rect 19182 22318 19234 22370
rect 19630 22318 19682 22370
rect 20526 22318 20578 22370
rect 21310 22318 21362 22370
rect 21758 22318 21810 22370
rect 22430 22318 22482 22370
rect 22990 22318 23042 22370
rect 23662 22318 23714 22370
rect 29038 22318 29090 22370
rect 29374 22318 29426 22370
rect 37886 22318 37938 22370
rect 14030 22206 14082 22258
rect 16494 22206 16546 22258
rect 18286 22206 18338 22258
rect 19294 22206 19346 22258
rect 22094 22206 22146 22258
rect 24222 22206 24274 22258
rect 29262 22206 29314 22258
rect 13582 22094 13634 22146
rect 17726 22094 17778 22146
rect 23998 22094 24050 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 17390 21758 17442 21810
rect 17726 21758 17778 21810
rect 12350 21646 12402 21698
rect 4286 21534 4338 21586
rect 11566 21534 11618 21586
rect 16270 21534 16322 21586
rect 16382 21534 16434 21586
rect 18510 21534 18562 21586
rect 19406 21534 19458 21586
rect 25342 21534 25394 21586
rect 28590 21534 28642 21586
rect 37662 21534 37714 21586
rect 14478 21422 14530 21474
rect 14926 21422 14978 21474
rect 16158 21422 16210 21474
rect 18734 21422 18786 21474
rect 23326 21422 23378 21474
rect 26014 21422 26066 21474
rect 28142 21422 28194 21474
rect 29262 21422 29314 21474
rect 31390 21422 31442 21474
rect 39902 21422 39954 21474
rect 1934 21310 1986 21362
rect 15710 21310 15762 21362
rect 18174 21310 18226 21362
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 17838 20974 17890 21026
rect 21870 20974 21922 21026
rect 9998 20862 10050 20914
rect 13582 20862 13634 20914
rect 14254 20862 14306 20914
rect 19294 20862 19346 20914
rect 19742 20862 19794 20914
rect 20526 20862 20578 20914
rect 25342 20862 25394 20914
rect 29598 20862 29650 20914
rect 40014 20862 40066 20914
rect 12126 20750 12178 20802
rect 12798 20750 12850 20802
rect 14142 20750 14194 20802
rect 14814 20750 14866 20802
rect 15822 20750 15874 20802
rect 16830 20750 16882 20802
rect 18062 20750 18114 20802
rect 18622 20750 18674 20802
rect 19070 20750 19122 20802
rect 19854 20750 19906 20802
rect 21534 20750 21586 20802
rect 21870 20750 21922 20802
rect 23326 20750 23378 20802
rect 29486 20750 29538 20802
rect 29710 20750 29762 20802
rect 30046 20750 30098 20802
rect 30606 20750 30658 20802
rect 37662 20750 37714 20802
rect 15374 20638 15426 20690
rect 21310 20638 21362 20690
rect 22766 20638 22818 20690
rect 29150 20638 29202 20690
rect 30158 20638 30210 20690
rect 30718 20638 30770 20690
rect 14366 20526 14418 20578
rect 14590 20526 14642 20578
rect 15150 20526 15202 20578
rect 15262 20526 15314 20578
rect 17166 20526 17218 20578
rect 17502 20526 17554 20578
rect 18398 20526 18450 20578
rect 18510 20526 18562 20578
rect 21758 20526 21810 20578
rect 22430 20526 22482 20578
rect 30382 20526 30434 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 24558 20190 24610 20242
rect 15710 20078 15762 20130
rect 19406 20078 19458 20130
rect 23102 20078 23154 20130
rect 23326 20078 23378 20130
rect 24334 20078 24386 20130
rect 24446 20078 24498 20130
rect 24670 20078 24722 20130
rect 25230 20078 25282 20130
rect 26238 20078 26290 20130
rect 26686 20078 26738 20130
rect 26798 20078 26850 20130
rect 15486 19966 15538 20018
rect 22542 19966 22594 20018
rect 22990 19966 23042 20018
rect 23886 19966 23938 20018
rect 25566 19966 25618 20018
rect 25678 19966 25730 20018
rect 26126 19966 26178 20018
rect 26462 19966 26514 20018
rect 27694 19966 27746 20018
rect 37662 19966 37714 20018
rect 14142 19854 14194 19906
rect 25342 19854 25394 19906
rect 27358 19854 27410 19906
rect 28478 19854 28530 19906
rect 30606 19854 30658 19906
rect 40014 19742 40066 19794
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 28366 19406 28418 19458
rect 1934 19294 1986 19346
rect 21758 19294 21810 19346
rect 27246 19294 27298 19346
rect 4286 19182 4338 19234
rect 13470 19182 13522 19234
rect 13806 19182 13858 19234
rect 14814 19182 14866 19234
rect 15038 19182 15090 19234
rect 16270 19182 16322 19234
rect 16942 19182 16994 19234
rect 18286 19182 18338 19234
rect 18846 19182 18898 19234
rect 20302 19182 20354 19234
rect 21198 19182 21250 19234
rect 21534 19182 21586 19234
rect 24334 19182 24386 19234
rect 28478 19182 28530 19234
rect 14030 19070 14082 19122
rect 14366 19070 14418 19122
rect 14702 19070 14754 19122
rect 15934 19070 15986 19122
rect 16606 19070 16658 19122
rect 18510 19070 18562 19122
rect 19966 19070 20018 19122
rect 21758 19070 21810 19122
rect 22430 19070 22482 19122
rect 25118 19070 25170 19122
rect 13582 18958 13634 19010
rect 14590 18958 14642 19010
rect 16046 18958 16098 19010
rect 19182 18958 19234 19010
rect 22094 18958 22146 19010
rect 27694 18958 27746 19010
rect 28366 18958 28418 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 17502 18622 17554 18674
rect 23438 18622 23490 18674
rect 14366 18510 14418 18562
rect 15486 18510 15538 18562
rect 15822 18510 15874 18562
rect 17614 18510 17666 18562
rect 18622 18510 18674 18562
rect 19518 18510 19570 18562
rect 20526 18510 20578 18562
rect 22542 18510 22594 18562
rect 25342 18510 25394 18562
rect 25566 18510 25618 18562
rect 4286 18398 4338 18450
rect 13134 18398 13186 18450
rect 13918 18398 13970 18450
rect 14590 18398 14642 18450
rect 14814 18398 14866 18450
rect 15038 18398 15090 18450
rect 15262 18398 15314 18450
rect 16606 18398 16658 18450
rect 17278 18398 17330 18450
rect 18062 18398 18114 18450
rect 18286 18398 18338 18450
rect 19070 18398 19122 18450
rect 19182 18398 19234 18450
rect 19406 18398 19458 18450
rect 19854 18398 19906 18450
rect 22094 18398 22146 18450
rect 11006 18286 11058 18338
rect 15710 18286 15762 18338
rect 18174 18286 18226 18338
rect 25230 18286 25282 18338
rect 1934 18174 1986 18226
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 22990 17838 23042 17890
rect 23662 17838 23714 17890
rect 13470 17726 13522 17778
rect 15598 17726 15650 17778
rect 21646 17726 21698 17778
rect 22766 17726 22818 17778
rect 27918 17726 27970 17778
rect 40014 17726 40066 17778
rect 16270 17614 16322 17666
rect 16830 17614 16882 17666
rect 16942 17614 16994 17666
rect 17166 17614 17218 17666
rect 17950 17614 18002 17666
rect 19630 17614 19682 17666
rect 20190 17614 20242 17666
rect 20750 17614 20802 17666
rect 21870 17614 21922 17666
rect 22430 17614 22482 17666
rect 23774 17614 23826 17666
rect 23998 17614 24050 17666
rect 27806 17614 27858 17666
rect 29150 17614 29202 17666
rect 37662 17614 37714 17666
rect 17614 17502 17666 17554
rect 19406 17502 19458 17554
rect 19966 17502 20018 17554
rect 21422 17502 21474 17554
rect 22094 17502 22146 17554
rect 27358 17502 27410 17554
rect 27582 17502 27634 17554
rect 27918 17502 27970 17554
rect 29262 17502 29314 17554
rect 17054 17390 17106 17442
rect 17278 17390 17330 17442
rect 17838 17390 17890 17442
rect 21982 17390 22034 17442
rect 23326 17390 23378 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 17502 17054 17554 17106
rect 18734 17054 18786 17106
rect 14702 16942 14754 16994
rect 22094 16942 22146 16994
rect 28030 16942 28082 16994
rect 14030 16830 14082 16882
rect 20302 16830 20354 16882
rect 21422 16830 21474 16882
rect 24670 16830 24722 16882
rect 26910 16830 26962 16882
rect 27246 16830 27298 16882
rect 37662 16830 37714 16882
rect 16830 16718 16882 16770
rect 18846 16718 18898 16770
rect 19070 16718 19122 16770
rect 20078 16718 20130 16770
rect 24222 16718 24274 16770
rect 30158 16718 30210 16770
rect 18734 16606 18786 16658
rect 19294 16606 19346 16658
rect 19742 16606 19794 16658
rect 19854 16606 19906 16658
rect 40014 16606 40066 16658
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 18174 16270 18226 16322
rect 18510 16270 18562 16322
rect 19182 16270 19234 16322
rect 19294 16270 19346 16322
rect 19518 16270 19570 16322
rect 20078 16270 20130 16322
rect 20302 16270 20354 16322
rect 21758 16270 21810 16322
rect 21422 16158 21474 16210
rect 24670 16158 24722 16210
rect 25118 16158 25170 16210
rect 28590 16158 28642 16210
rect 29262 16158 29314 16210
rect 18510 16046 18562 16098
rect 19630 16046 19682 16098
rect 20526 16046 20578 16098
rect 20750 16046 20802 16098
rect 25678 16046 25730 16098
rect 24446 15934 24498 15986
rect 25006 15934 25058 15986
rect 26462 15934 26514 15986
rect 20638 15822 20690 15874
rect 21534 15822 21586 15874
rect 24558 15822 24610 15874
rect 25230 15822 25282 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 26686 15486 26738 15538
rect 17390 15374 17442 15426
rect 17726 15374 17778 15426
rect 18734 15374 18786 15426
rect 20190 15374 20242 15426
rect 20526 15374 20578 15426
rect 18510 15262 18562 15314
rect 26910 15262 26962 15314
rect 27358 15262 27410 15314
rect 27582 15262 27634 15314
rect 26574 15150 26626 15202
rect 27246 15038 27298 15090
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 18958 14702 19010 14754
rect 19294 14702 19346 14754
rect 16606 14590 16658 14642
rect 18734 14590 18786 14642
rect 24222 14590 24274 14642
rect 26350 14590 26402 14642
rect 26910 14590 26962 14642
rect 15934 14478 15986 14530
rect 23550 14478 23602 14530
rect 19182 14254 19234 14306
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 20078 13806 20130 13858
rect 19406 13694 19458 13746
rect 22654 13694 22706 13746
rect 22206 13582 22258 13634
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 18734 5182 18786 5234
rect 17726 5070 17778 5122
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 24446 4398 24498 4450
rect 19070 4286 19122 4338
rect 25790 4286 25842 4338
rect 20078 4062 20130 4114
rect 26798 4062 26850 4114
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 18174 3614 18226 3666
rect 25566 3614 25618 3666
rect 19742 3502 19794 3554
rect 21422 3502 21474 3554
rect 24558 3502 24610 3554
rect 22430 3278 22482 3330
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
<< metal2 >>
rect 18144 41200 18256 42000
rect 20832 41200 20944 42000
rect 22176 41200 22288 42000
rect 22848 41200 22960 42000
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 18172 38162 18228 41200
rect 18172 38110 18174 38162
rect 18226 38110 18228 38162
rect 18172 38098 18228 38110
rect 19740 38052 19796 38062
rect 19404 38050 19796 38052
rect 19404 37998 19742 38050
rect 19794 37998 19796 38050
rect 19404 37996 19796 37998
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 17836 28642 17892 28654
rect 17836 28590 17838 28642
rect 17890 28590 17892 28642
rect 14364 27858 14420 27870
rect 14364 27806 14366 27858
rect 14418 27806 14420 27858
rect 11452 27746 11508 27758
rect 11452 27694 11454 27746
rect 11506 27694 11508 27746
rect 4172 27636 4228 27646
rect 1932 27186 1988 27198
rect 1932 27134 1934 27186
rect 1986 27134 1988 27186
rect 1932 26292 1988 27134
rect 1932 26226 1988 26236
rect 2044 26964 2100 26974
rect 2044 26178 2100 26908
rect 2044 26126 2046 26178
rect 2098 26126 2100 26178
rect 2044 26114 2100 26126
rect 4172 21700 4228 27580
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 4284 27076 4340 27086
rect 4284 26982 4340 27020
rect 11452 26964 11508 27694
rect 13580 27748 13636 27758
rect 14364 27748 14420 27806
rect 14812 27748 14868 27758
rect 13580 27746 13972 27748
rect 13580 27694 13582 27746
rect 13634 27694 13972 27746
rect 13580 27692 13972 27694
rect 14364 27746 14868 27748
rect 14364 27694 14814 27746
rect 14866 27694 14868 27746
rect 14364 27692 14868 27694
rect 13580 27682 13636 27692
rect 13916 27298 13972 27692
rect 13916 27246 13918 27298
rect 13970 27246 13972 27298
rect 13916 27234 13972 27246
rect 11452 26898 11508 26908
rect 13468 26962 13524 26974
rect 13468 26910 13470 26962
rect 13522 26910 13524 26962
rect 13468 26740 13524 26910
rect 14028 26964 14084 26974
rect 14364 26964 14420 26974
rect 14028 26962 14308 26964
rect 14028 26910 14030 26962
rect 14082 26910 14308 26962
rect 14028 26908 14308 26910
rect 14028 26898 14084 26908
rect 13580 26852 13636 26862
rect 13580 26850 13860 26852
rect 13580 26798 13582 26850
rect 13634 26798 13860 26850
rect 13580 26796 13860 26798
rect 13580 26786 13636 26796
rect 13468 26674 13524 26684
rect 13804 26404 13860 26796
rect 13916 26404 13972 26414
rect 13804 26402 13972 26404
rect 13804 26350 13918 26402
rect 13970 26350 13972 26402
rect 13804 26348 13972 26350
rect 13916 26338 13972 26348
rect 4284 26292 4340 26302
rect 4284 26198 4340 26236
rect 11788 26292 11844 26302
rect 11788 26178 11844 26236
rect 11788 26126 11790 26178
rect 11842 26126 11844 26178
rect 11788 26114 11844 26126
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 14252 25618 14308 26908
rect 14252 25566 14254 25618
rect 14306 25566 14308 25618
rect 14252 25554 14308 25566
rect 14028 25506 14084 25518
rect 14028 25454 14030 25506
rect 14082 25454 14084 25506
rect 14028 25396 14084 25454
rect 14364 25506 14420 26908
rect 14812 26852 14868 27692
rect 17052 27074 17108 27086
rect 17052 27022 17054 27074
rect 17106 27022 17108 27074
rect 14924 26852 14980 26862
rect 14812 26850 14980 26852
rect 14812 26798 14926 26850
rect 14978 26798 14980 26850
rect 14812 26796 14980 26798
rect 14700 26292 14756 26302
rect 14812 26292 14868 26796
rect 14924 26516 14980 26796
rect 17052 26852 17108 27022
rect 17724 26964 17780 26974
rect 17724 26870 17780 26908
rect 17052 26786 17108 26796
rect 17836 26852 17892 28590
rect 18620 28532 18676 28542
rect 18620 28530 19236 28532
rect 18620 28478 18622 28530
rect 18674 28478 19236 28530
rect 18620 28476 19236 28478
rect 18620 28466 18676 28476
rect 19180 28082 19236 28476
rect 19180 28030 19182 28082
rect 19234 28030 19236 28082
rect 19180 28018 19236 28030
rect 18732 27860 18788 27870
rect 19068 27860 19124 27870
rect 14924 26450 14980 26460
rect 15372 26740 15428 26750
rect 15372 26514 15428 26684
rect 15372 26462 15374 26514
rect 15426 26462 15428 26514
rect 15372 26450 15428 26462
rect 15596 26516 15652 26526
rect 14700 26290 14868 26292
rect 14700 26238 14702 26290
rect 14754 26238 14868 26290
rect 14700 26236 14868 26238
rect 15036 26290 15092 26302
rect 15036 26238 15038 26290
rect 15090 26238 15092 26290
rect 14700 26226 14756 26236
rect 14364 25454 14366 25506
rect 14418 25454 14420 25506
rect 14364 25442 14420 25454
rect 14588 25732 14644 25742
rect 14588 25506 14644 25676
rect 15036 25732 15092 26238
rect 15260 26292 15316 26302
rect 15484 26292 15540 26302
rect 15260 26198 15316 26236
rect 15372 26290 15540 26292
rect 15372 26238 15486 26290
rect 15538 26238 15540 26290
rect 15372 26236 15540 26238
rect 15036 25666 15092 25676
rect 14588 25454 14590 25506
rect 14642 25454 14644 25506
rect 14588 25442 14644 25454
rect 13804 25340 14028 25396
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 13468 24164 13524 24174
rect 13524 24108 13748 24164
rect 13468 24070 13524 24108
rect 13580 23714 13636 23726
rect 13580 23662 13582 23714
rect 13634 23662 13636 23714
rect 13580 23604 13636 23662
rect 13020 23548 13636 23604
rect 13020 23266 13076 23548
rect 13020 23214 13022 23266
rect 13074 23214 13076 23266
rect 13020 23202 13076 23214
rect 12236 23154 12292 23166
rect 12236 23102 12238 23154
rect 12290 23102 12292 23154
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 4172 21634 4228 21644
rect 4284 21588 4340 21598
rect 4284 21494 4340 21532
rect 9996 21588 10052 21598
rect 1932 21362 1988 21374
rect 1932 21310 1934 21362
rect 1986 21310 1988 21362
rect 1932 20916 1988 21310
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 1932 20850 1988 20860
rect 9996 20914 10052 21532
rect 11564 21588 11620 21598
rect 11564 21494 11620 21532
rect 12236 21588 12292 23102
rect 13692 22932 13748 24108
rect 13804 23938 13860 25340
rect 14028 25330 14084 25340
rect 15372 25396 15428 26236
rect 15484 26226 15540 26236
rect 15372 25330 15428 25340
rect 15484 25620 15540 25630
rect 15596 25620 15652 26460
rect 15540 25564 15652 25620
rect 15708 26290 15764 26302
rect 15708 26238 15710 26290
rect 15762 26238 15764 26290
rect 15484 25506 15540 25564
rect 15484 25454 15486 25506
rect 15538 25454 15540 25506
rect 13804 23886 13806 23938
rect 13858 23886 13860 23938
rect 13804 23874 13860 23886
rect 14140 25282 14196 25294
rect 14140 25230 14142 25282
rect 14194 25230 14196 25282
rect 14140 23940 14196 25230
rect 14252 24052 14308 24062
rect 14252 23958 14308 23996
rect 15372 24052 15428 24062
rect 15484 24052 15540 25454
rect 15372 24050 15540 24052
rect 15372 23998 15374 24050
rect 15426 23998 15540 24050
rect 15372 23996 15540 23998
rect 15708 24052 15764 26238
rect 17836 25620 17892 26796
rect 18620 27076 18676 27086
rect 18620 26292 18676 27020
rect 18732 26964 18788 27804
rect 18732 26514 18788 26908
rect 18956 27858 19124 27860
rect 18956 27806 19070 27858
rect 19122 27806 19124 27858
rect 18956 27804 19124 27806
rect 18956 26964 19012 27804
rect 19068 27794 19124 27804
rect 19292 27860 19348 27870
rect 19292 27766 19348 27804
rect 19404 27636 19460 37996
rect 19740 37986 19796 37996
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 20860 37492 20916 41200
rect 22204 38162 22260 41200
rect 22876 38276 22932 41200
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 22876 38210 22932 38220
rect 25564 38276 25620 38286
rect 25564 38182 25620 38220
rect 22204 38110 22206 38162
rect 22258 38110 22260 38162
rect 22204 38098 22260 38110
rect 23772 38050 23828 38062
rect 23772 37998 23774 38050
rect 23826 37998 23828 38050
rect 20860 37426 20916 37436
rect 22092 37492 22148 37502
rect 22092 37398 22148 37436
rect 21084 37266 21140 37278
rect 21084 37214 21086 37266
rect 21138 37214 21140 37266
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 21084 31948 21140 37214
rect 20748 31892 21140 31948
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 20748 28756 20804 31892
rect 20188 28754 20804 28756
rect 20188 28702 20750 28754
rect 20802 28702 20804 28754
rect 20188 28700 20804 28702
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 20076 28084 20132 28094
rect 20188 28084 20244 28700
rect 20748 28690 20804 28700
rect 21420 28420 21476 28430
rect 20076 28082 20244 28084
rect 20076 28030 20078 28082
rect 20130 28030 20244 28082
rect 20076 28028 20244 28030
rect 21084 28418 21476 28420
rect 21084 28366 21422 28418
rect 21474 28366 21476 28418
rect 21084 28364 21476 28366
rect 20076 28018 20132 28028
rect 19852 27970 19908 27982
rect 19852 27918 19854 27970
rect 19906 27918 19908 27970
rect 19740 27860 19796 27870
rect 19852 27860 19908 27918
rect 19740 27858 19908 27860
rect 19740 27806 19742 27858
rect 19794 27806 19908 27858
rect 19740 27804 19908 27806
rect 20188 27860 20244 27870
rect 20636 27860 20692 27870
rect 20188 27858 20356 27860
rect 20188 27806 20190 27858
rect 20242 27806 20356 27858
rect 20188 27804 20356 27806
rect 19740 27794 19796 27804
rect 20188 27794 20244 27804
rect 18956 26898 19012 26908
rect 19068 27580 19460 27636
rect 18732 26462 18734 26514
rect 18786 26462 18788 26514
rect 18732 26450 18788 26462
rect 18508 26290 18676 26292
rect 18508 26238 18622 26290
rect 18674 26238 18676 26290
rect 18508 26236 18676 26238
rect 17836 25554 17892 25564
rect 18284 25732 18340 25742
rect 18284 25618 18340 25676
rect 18284 25566 18286 25618
rect 18338 25566 18340 25618
rect 18284 25554 18340 25566
rect 16156 25394 16212 25406
rect 16156 25342 16158 25394
rect 16210 25342 16212 25394
rect 16156 24948 16212 25342
rect 16156 24882 16212 24892
rect 16492 25396 16548 25406
rect 15372 23986 15428 23996
rect 15708 23986 15764 23996
rect 16492 24724 16548 25340
rect 17948 25284 18004 25294
rect 17500 24948 17556 24958
rect 17500 24854 17556 24892
rect 15596 23940 15652 23950
rect 14140 23874 14196 23884
rect 15484 23884 15596 23940
rect 14140 23716 14196 23726
rect 13468 22876 13748 22932
rect 13804 23714 14196 23716
rect 13804 23662 14142 23714
rect 14194 23662 14196 23714
rect 13804 23660 14196 23662
rect 13468 22370 13524 22876
rect 13468 22318 13470 22370
rect 13522 22318 13524 22370
rect 13468 22306 13524 22318
rect 13804 22370 13860 23660
rect 14140 23650 14196 23660
rect 15148 23042 15204 23054
rect 15148 22990 15150 23042
rect 15202 22990 15204 23042
rect 14812 22932 14868 22942
rect 13804 22318 13806 22370
rect 13858 22318 13860 22370
rect 13804 22306 13860 22318
rect 14476 22372 14532 22382
rect 14028 22258 14084 22270
rect 14028 22206 14030 22258
rect 14082 22206 14084 22258
rect 12348 22148 12404 22158
rect 12348 21698 12404 22092
rect 13580 22148 13636 22158
rect 13580 22054 13636 22092
rect 14028 22148 14084 22206
rect 14028 22082 14084 22092
rect 12348 21646 12350 21698
rect 12402 21646 12404 21698
rect 12348 21634 12404 21646
rect 12236 21522 12292 21532
rect 12796 21588 12852 21598
rect 9996 20862 9998 20914
rect 10050 20862 10052 20914
rect 9996 20692 10052 20862
rect 12796 20916 12852 21532
rect 14476 21474 14532 22316
rect 14476 21422 14478 21474
rect 14530 21422 14532 21474
rect 14476 21410 14532 21422
rect 14252 21364 14308 21374
rect 14140 21308 14252 21364
rect 12124 20804 12180 20814
rect 12124 20710 12180 20748
rect 12796 20802 12852 20860
rect 12796 20750 12798 20802
rect 12850 20750 12852 20802
rect 12796 20738 12852 20750
rect 13580 20916 13636 20926
rect 9996 20626 10052 20636
rect 13468 20244 13524 20254
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 1932 19346 1988 19358
rect 1932 19294 1934 19346
rect 1986 19294 1988 19346
rect 1932 18900 1988 19294
rect 4284 19236 4340 19246
rect 4284 19142 4340 19180
rect 13468 19234 13524 20188
rect 13580 19908 13636 20860
rect 14140 20802 14196 21308
rect 14252 21298 14308 21308
rect 14140 20750 14142 20802
rect 14194 20750 14196 20802
rect 14140 20244 14196 20750
rect 14252 20914 14308 20926
rect 14252 20862 14254 20914
rect 14306 20862 14308 20914
rect 14252 20804 14308 20862
rect 14252 20738 14308 20748
rect 14812 20802 14868 22876
rect 15148 22820 15204 22990
rect 15148 22754 15204 22764
rect 15148 22148 15204 22158
rect 14924 21474 14980 21486
rect 14924 21422 14926 21474
rect 14978 21422 14980 21474
rect 14924 20916 14980 21422
rect 14924 20850 14980 20860
rect 14812 20750 14814 20802
rect 14866 20750 14868 20802
rect 14812 20738 14868 20750
rect 14364 20578 14420 20590
rect 14364 20526 14366 20578
rect 14418 20526 14420 20578
rect 14364 20188 14420 20526
rect 14588 20580 14644 20590
rect 14588 20486 14644 20524
rect 15148 20578 15204 22092
rect 15372 20692 15428 20702
rect 15372 20598 15428 20636
rect 15148 20526 15150 20578
rect 15202 20526 15204 20578
rect 14140 20132 14308 20188
rect 14364 20132 14868 20188
rect 14140 19908 14196 19918
rect 13580 19906 14196 19908
rect 13580 19854 14142 19906
rect 14194 19854 14196 19906
rect 13580 19852 14196 19854
rect 13468 19182 13470 19234
rect 13522 19182 13524 19234
rect 13468 19170 13524 19182
rect 13804 19236 13860 19246
rect 13804 19142 13860 19180
rect 14028 19124 14084 19134
rect 14028 19030 14084 19068
rect 13580 19012 13636 19022
rect 13132 19010 13636 19012
rect 13132 18958 13582 19010
rect 13634 18958 13636 19010
rect 13132 18956 13636 18958
rect 1932 18834 1988 18844
rect 11004 18900 11060 18910
rect 4284 18450 4340 18462
rect 4284 18398 4286 18450
rect 4338 18398 4340 18450
rect 4284 18340 4340 18398
rect 4284 18274 4340 18284
rect 11004 18338 11060 18844
rect 13132 18450 13188 18956
rect 13580 18946 13636 18956
rect 13132 18398 13134 18450
rect 13186 18398 13188 18450
rect 13132 18386 13188 18398
rect 13916 18452 13972 18462
rect 14140 18452 14196 19852
rect 14252 18564 14308 20132
rect 14812 19236 14868 20132
rect 14812 19142 14868 19180
rect 15036 19348 15092 19358
rect 15036 19234 15092 19292
rect 15036 19182 15038 19234
rect 15090 19182 15092 19234
rect 15036 19170 15092 19182
rect 14364 19122 14420 19134
rect 14364 19070 14366 19122
rect 14418 19070 14420 19122
rect 14364 18900 14420 19070
rect 14700 19124 14756 19134
rect 14700 19030 14756 19068
rect 14364 18834 14420 18844
rect 14588 19010 14644 19022
rect 14588 18958 14590 19010
rect 14642 18958 14644 19010
rect 14588 18676 14644 18958
rect 14588 18620 14980 18676
rect 14364 18564 14420 18574
rect 14252 18562 14420 18564
rect 14252 18510 14366 18562
rect 14418 18510 14420 18562
rect 14252 18508 14420 18510
rect 14924 18564 14980 18620
rect 15036 18564 15092 18574
rect 14924 18508 15036 18564
rect 14364 18498 14420 18508
rect 13916 18450 14196 18452
rect 13916 18398 13918 18450
rect 13970 18398 14196 18450
rect 13916 18396 14196 18398
rect 13916 18386 13972 18396
rect 11004 18286 11006 18338
rect 11058 18286 11060 18338
rect 11004 18274 11060 18286
rect 13468 18340 13524 18350
rect 1932 18228 1988 18238
rect 1932 18134 1988 18172
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 13468 17778 13524 18284
rect 13468 17726 13470 17778
rect 13522 17726 13524 17778
rect 13468 17714 13524 17726
rect 14140 18340 14196 18396
rect 14588 18452 14644 18462
rect 14588 18358 14644 18396
rect 14812 18452 14868 18462
rect 14812 18358 14868 18396
rect 15036 18450 15092 18508
rect 15036 18398 15038 18450
rect 15090 18398 15092 18450
rect 15036 18386 15092 18398
rect 14028 16884 14084 16894
rect 14140 16884 14196 18284
rect 15148 17892 15204 20526
rect 15260 20580 15316 20590
rect 15484 20580 15540 23884
rect 15596 23874 15652 23884
rect 16268 23492 16324 23502
rect 15820 23156 15876 23166
rect 15596 23154 15876 23156
rect 15596 23102 15822 23154
rect 15874 23102 15876 23154
rect 15596 23100 15876 23102
rect 15596 22372 15652 23100
rect 15820 23090 15876 23100
rect 15596 22278 15652 22316
rect 16044 22372 16100 22382
rect 16156 22372 16212 22382
rect 16044 22370 16156 22372
rect 16044 22318 16046 22370
rect 16098 22318 16156 22370
rect 16044 22316 16156 22318
rect 16044 22306 16100 22316
rect 16156 21474 16212 22316
rect 16268 21586 16324 23436
rect 16380 23042 16436 23054
rect 16380 22990 16382 23042
rect 16434 22990 16436 23042
rect 16380 21924 16436 22990
rect 16492 22258 16548 24668
rect 17388 24836 17444 24846
rect 17388 24724 17444 24780
rect 17948 24834 18004 25228
rect 18508 24948 18564 26236
rect 18620 26226 18676 26236
rect 19068 25732 19124 27580
rect 19852 27188 19908 27198
rect 20300 27188 20356 27804
rect 20636 27766 20692 27804
rect 19852 27186 20244 27188
rect 19852 27134 19854 27186
rect 19906 27134 20244 27186
rect 19852 27132 20244 27134
rect 19852 27122 19908 27132
rect 20188 27074 20244 27132
rect 20188 27022 20190 27074
rect 20242 27022 20244 27074
rect 19404 26964 19460 26974
rect 19068 25506 19124 25676
rect 19068 25454 19070 25506
rect 19122 25454 19124 25506
rect 19068 25442 19124 25454
rect 19292 26852 19460 26908
rect 18396 24892 18564 24948
rect 18620 25394 18676 25406
rect 18620 25342 18622 25394
rect 18674 25342 18676 25394
rect 17948 24782 17950 24834
rect 18002 24782 18004 24834
rect 17948 24770 18004 24782
rect 18284 24836 18340 24846
rect 18284 24742 18340 24780
rect 17612 24724 17668 24734
rect 17388 24722 17556 24724
rect 17388 24670 17390 24722
rect 17442 24670 17556 24722
rect 17388 24668 17556 24670
rect 17388 24658 17444 24668
rect 17500 24052 17556 24668
rect 17612 24630 17668 24668
rect 18396 24612 18452 24892
rect 18620 24836 18676 25342
rect 18620 24770 18676 24780
rect 18844 25282 18900 25294
rect 18844 25230 18846 25282
rect 18898 25230 18900 25282
rect 17388 23268 17444 23278
rect 16492 22206 16494 22258
rect 16546 22206 16548 22258
rect 16492 22194 16548 22206
rect 16716 22370 16772 22382
rect 16716 22318 16718 22370
rect 16770 22318 16772 22370
rect 16380 21858 16436 21868
rect 16492 22036 16548 22046
rect 16268 21534 16270 21586
rect 16322 21534 16324 21586
rect 16268 21522 16324 21534
rect 16380 21588 16436 21598
rect 16492 21588 16548 21980
rect 16380 21586 16548 21588
rect 16380 21534 16382 21586
rect 16434 21534 16548 21586
rect 16380 21532 16548 21534
rect 16156 21422 16158 21474
rect 16210 21422 16212 21474
rect 16156 21410 16212 21422
rect 15708 21364 15764 21374
rect 15708 21270 15764 21308
rect 15820 20916 15876 20926
rect 15820 20802 15876 20860
rect 15820 20750 15822 20802
rect 15874 20750 15876 20802
rect 15820 20738 15876 20750
rect 15484 20524 15764 20580
rect 15260 20486 15316 20524
rect 15708 20130 15764 20524
rect 15708 20078 15710 20130
rect 15762 20078 15764 20130
rect 15484 20018 15540 20030
rect 15484 19966 15486 20018
rect 15538 19966 15540 20018
rect 15484 19796 15540 19966
rect 15484 19730 15540 19740
rect 15484 19236 15540 19246
rect 15484 18562 15540 19180
rect 15484 18510 15486 18562
rect 15538 18510 15540 18562
rect 15484 18498 15540 18510
rect 15708 18564 15764 20078
rect 16268 19236 16324 19246
rect 16380 19236 16436 21532
rect 16716 21028 16772 22318
rect 16716 20962 16772 20972
rect 16828 21924 16884 21934
rect 16828 20802 16884 21868
rect 17388 21812 17444 23212
rect 16828 20750 16830 20802
rect 16882 20750 16884 20802
rect 16828 20738 16884 20750
rect 16940 21810 17444 21812
rect 16940 21758 17390 21810
rect 17442 21758 17444 21810
rect 16940 21756 17444 21758
rect 16268 19234 16436 19236
rect 16268 19182 16270 19234
rect 16322 19182 16436 19234
rect 16268 19180 16436 19182
rect 16604 19236 16660 19246
rect 16268 19170 16324 19180
rect 15932 19122 15988 19134
rect 15932 19070 15934 19122
rect 15986 19070 15988 19122
rect 15820 18564 15876 18574
rect 15708 18562 15876 18564
rect 15708 18510 15822 18562
rect 15874 18510 15876 18562
rect 15708 18508 15876 18510
rect 15260 18452 15316 18462
rect 15260 18358 15316 18396
rect 15708 18340 15764 18350
rect 15148 17826 15204 17836
rect 15596 18338 15764 18340
rect 15596 18286 15710 18338
rect 15762 18286 15764 18338
rect 15596 18284 15764 18286
rect 15596 17778 15652 18284
rect 15708 18274 15764 18284
rect 15596 17726 15598 17778
rect 15650 17726 15652 17778
rect 15596 17714 15652 17726
rect 14700 17444 14756 17454
rect 14700 16994 14756 17388
rect 15820 17332 15876 18508
rect 15932 17892 15988 19070
rect 16604 19122 16660 19180
rect 16940 19236 16996 21756
rect 17388 21746 17444 21756
rect 17500 21588 17556 23996
rect 18284 24556 18452 24612
rect 18508 24722 18564 24734
rect 18508 24670 18510 24722
rect 18562 24670 18564 24722
rect 17724 23826 17780 23838
rect 17724 23774 17726 23826
rect 17778 23774 17780 23826
rect 17612 23156 17668 23166
rect 17724 23156 17780 23774
rect 18060 23826 18116 23838
rect 18060 23774 18062 23826
rect 18114 23774 18116 23826
rect 18060 23716 18116 23774
rect 18060 23650 18116 23660
rect 17612 23154 17780 23156
rect 17612 23102 17614 23154
rect 17666 23102 17780 23154
rect 17612 23100 17780 23102
rect 17612 22820 17668 23100
rect 17612 22754 17668 22764
rect 18060 23042 18116 23054
rect 18060 22990 18062 23042
rect 18114 22990 18116 23042
rect 17612 22484 17668 22494
rect 17612 22370 17668 22428
rect 17612 22318 17614 22370
rect 17666 22318 17668 22370
rect 17612 21924 17668 22318
rect 17724 22148 17780 22158
rect 17724 22054 17780 22092
rect 17612 21858 17668 21868
rect 17724 21812 17780 21822
rect 17724 21718 17780 21756
rect 18060 21812 18116 22990
rect 18284 22260 18340 24556
rect 18508 24500 18564 24670
rect 18844 24500 18900 25230
rect 18956 25284 19012 25294
rect 18956 25190 19012 25228
rect 19180 25284 19236 25294
rect 19180 25190 19236 25228
rect 18284 22166 18340 22204
rect 18396 24444 18900 24500
rect 18956 24836 19012 24846
rect 18396 23156 18452 24444
rect 18508 24164 18564 24174
rect 18508 23714 18564 24108
rect 18844 24052 18900 24062
rect 18956 24052 19012 24780
rect 18844 24050 19012 24052
rect 18844 23998 18846 24050
rect 18898 23998 19012 24050
rect 18844 23996 19012 23998
rect 18508 23662 18510 23714
rect 18562 23662 18564 23714
rect 18508 23650 18564 23662
rect 18620 23940 18676 23950
rect 18620 23492 18676 23884
rect 18620 23426 18676 23436
rect 18844 23716 18900 23996
rect 18732 23380 18788 23390
rect 18732 23286 18788 23324
rect 18508 23268 18564 23278
rect 18508 23174 18564 23212
rect 18060 21746 18116 21756
rect 18396 21588 18452 23100
rect 17388 21532 17556 21588
rect 18060 21532 18452 21588
rect 18508 22820 18564 22830
rect 18508 21586 18564 22764
rect 18844 22596 18900 23660
rect 19068 23716 19124 23726
rect 18956 22932 19012 22942
rect 18956 22838 19012 22876
rect 18844 22530 18900 22540
rect 18508 21534 18510 21586
rect 18562 21534 18564 21586
rect 17164 20578 17220 20590
rect 17164 20526 17166 20578
rect 17218 20526 17220 20578
rect 17164 20244 17220 20526
rect 17388 20356 17444 21532
rect 17836 21028 17892 21038
rect 18060 21028 18116 21532
rect 18508 21522 18564 21534
rect 18620 22372 18676 22382
rect 17836 21026 18116 21028
rect 17836 20974 17838 21026
rect 17890 20974 18116 21026
rect 17836 20972 18116 20974
rect 18172 21362 18228 21374
rect 18172 21310 18174 21362
rect 18226 21310 18228 21362
rect 17836 20962 17892 20972
rect 18060 20802 18116 20814
rect 18060 20750 18062 20802
rect 18114 20750 18116 20802
rect 17500 20580 17556 20590
rect 18060 20580 18116 20750
rect 18172 20580 18228 21310
rect 18620 20802 18676 22316
rect 18732 22370 18788 22382
rect 18732 22318 18734 22370
rect 18786 22318 18788 22370
rect 18732 21812 18788 22318
rect 18732 21746 18788 21756
rect 18844 22260 18900 22270
rect 18732 21476 18788 21486
rect 18844 21476 18900 22204
rect 18788 21420 18900 21476
rect 18732 21382 18788 21420
rect 19068 21140 19124 23660
rect 19292 23380 19348 26852
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 20188 26290 20244 27022
rect 20188 26238 20190 26290
rect 20242 26238 20244 26290
rect 20188 26226 20244 26238
rect 20300 25844 20356 27132
rect 20748 27076 20804 27086
rect 20748 26982 20804 27020
rect 21084 26514 21140 28364
rect 21420 28354 21476 28364
rect 23772 28084 23828 37998
rect 24556 38050 24612 38062
rect 24556 37998 24558 38050
rect 24610 37998 24612 38050
rect 24556 31948 24612 37998
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 23436 28082 23828 28084
rect 23436 28030 23774 28082
rect 23826 28030 23828 28082
rect 23436 28028 23828 28030
rect 21308 27746 21364 27758
rect 21308 27694 21310 27746
rect 21362 27694 21364 27746
rect 21308 27188 21364 27694
rect 23436 27746 23492 28028
rect 23772 28018 23828 28028
rect 24108 31892 24612 31948
rect 24108 28082 24164 31892
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 24108 28030 24110 28082
rect 24162 28030 24164 28082
rect 24108 28018 24164 28030
rect 23436 27694 23438 27746
rect 23490 27694 23492 27746
rect 22316 27300 22372 27310
rect 21980 27298 22372 27300
rect 21980 27246 22318 27298
rect 22370 27246 22372 27298
rect 21980 27244 22372 27246
rect 21420 27188 21476 27198
rect 21308 27186 21476 27188
rect 21308 27134 21422 27186
rect 21474 27134 21476 27186
rect 21308 27132 21476 27134
rect 21420 27122 21476 27132
rect 21980 27074 22036 27244
rect 22316 27234 22372 27244
rect 21980 27022 21982 27074
rect 22034 27022 22036 27074
rect 21980 27010 22036 27022
rect 22204 27076 22260 27086
rect 22204 26982 22260 27020
rect 21308 26964 21364 26974
rect 21308 26870 21364 26908
rect 22316 26964 22372 26974
rect 22316 26870 22372 26908
rect 23436 26964 23492 27694
rect 23436 26898 23492 26908
rect 24668 27860 24724 27870
rect 21084 26462 21086 26514
rect 21138 26462 21140 26514
rect 20300 25778 20356 25788
rect 20636 26292 20692 26302
rect 19740 25620 19796 25630
rect 19628 25564 19740 25620
rect 19292 23154 19348 23324
rect 19516 23828 19572 23838
rect 19516 23156 19572 23772
rect 19292 23102 19294 23154
rect 19346 23102 19348 23154
rect 19292 23090 19348 23102
rect 19404 23154 19572 23156
rect 19404 23102 19518 23154
rect 19570 23102 19572 23154
rect 19404 23100 19572 23102
rect 19404 22594 19460 23100
rect 19516 23090 19572 23100
rect 19628 22596 19684 25564
rect 19740 25526 19796 25564
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 19852 23826 19908 23838
rect 19852 23774 19854 23826
rect 19906 23774 19908 23826
rect 19740 23716 19796 23754
rect 19852 23716 19908 23774
rect 19852 23660 20244 23716
rect 19740 23650 19796 23660
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 19852 23156 19908 23166
rect 19852 23062 19908 23100
rect 19404 22542 19406 22594
rect 19458 22542 19460 22594
rect 19404 22530 19460 22542
rect 19516 22540 19684 22596
rect 20188 23042 20244 23660
rect 20188 22990 20190 23042
rect 20242 22990 20244 23042
rect 19180 22372 19236 22382
rect 19180 22278 19236 22316
rect 19292 22258 19348 22270
rect 19292 22206 19294 22258
rect 19346 22206 19348 22258
rect 19292 22036 19348 22206
rect 19292 21970 19348 21980
rect 19404 21700 19460 21710
rect 19404 21586 19460 21644
rect 19404 21534 19406 21586
rect 19458 21534 19460 21586
rect 19404 21522 19460 21534
rect 19516 21364 19572 22540
rect 20076 22484 20132 22494
rect 20188 22484 20244 22990
rect 20412 23154 20468 23166
rect 20412 23102 20414 23154
rect 20466 23102 20468 23154
rect 20412 23044 20468 23102
rect 20412 22978 20468 22988
rect 20132 22428 20244 22484
rect 20076 22418 20132 22428
rect 19628 22370 19684 22382
rect 19628 22318 19630 22370
rect 19682 22318 19684 22370
rect 19628 21812 19684 22318
rect 20524 22372 20580 22382
rect 20636 22372 20692 26236
rect 21084 25620 21140 26462
rect 21532 26850 21588 26862
rect 21532 26798 21534 26850
rect 21586 26798 21588 26850
rect 21532 26292 21588 26798
rect 21532 26226 21588 26236
rect 21084 25554 21140 25564
rect 21644 25844 21700 25854
rect 21420 25506 21476 25518
rect 21420 25454 21422 25506
rect 21474 25454 21476 25506
rect 21420 25284 21476 25454
rect 21644 25394 21700 25788
rect 21644 25342 21646 25394
rect 21698 25342 21700 25394
rect 21644 25330 21700 25342
rect 21420 24052 21476 25228
rect 23548 24724 23604 24734
rect 21756 24612 21812 24622
rect 21420 23958 21476 23996
rect 21532 24610 21812 24612
rect 21532 24558 21758 24610
rect 21810 24558 21812 24610
rect 21532 24556 21812 24558
rect 21308 23826 21364 23838
rect 21308 23774 21310 23826
rect 21362 23774 21364 23826
rect 21308 23716 21364 23774
rect 21308 23650 21364 23660
rect 21420 23042 21476 23054
rect 21420 22990 21422 23042
rect 21474 22990 21476 23042
rect 20524 22370 20692 22372
rect 20524 22318 20526 22370
rect 20578 22318 20692 22370
rect 20524 22316 20692 22318
rect 20524 22306 20580 22316
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 19684 21756 19796 21812
rect 19628 21718 19684 21756
rect 18620 20750 18622 20802
rect 18674 20750 18676 20802
rect 18620 20738 18676 20750
rect 18956 21084 19124 21140
rect 19404 21308 19572 21364
rect 18396 20580 18452 20590
rect 17500 20578 17780 20580
rect 17500 20526 17502 20578
rect 17554 20526 17780 20578
rect 17500 20524 17780 20526
rect 18060 20578 18452 20580
rect 18060 20526 18398 20578
rect 18450 20526 18452 20578
rect 18060 20524 18452 20526
rect 17500 20514 17556 20524
rect 17388 20300 17668 20356
rect 17164 20178 17220 20188
rect 16940 19234 17108 19236
rect 16940 19182 16942 19234
rect 16994 19182 17108 19234
rect 16940 19180 17108 19182
rect 16940 19170 16996 19180
rect 16604 19070 16606 19122
rect 16658 19070 16660 19122
rect 16604 19058 16660 19070
rect 16044 19010 16100 19022
rect 16044 18958 16046 19010
rect 16098 18958 16100 19010
rect 16044 18564 16100 18958
rect 16044 18498 16100 18508
rect 16940 18564 16996 18574
rect 16604 18452 16660 18462
rect 16660 18396 16772 18452
rect 16604 18358 16660 18396
rect 15932 17826 15988 17836
rect 16268 18340 16324 18350
rect 16268 17666 16324 18284
rect 16268 17614 16270 17666
rect 16322 17614 16324 17666
rect 16268 17602 16324 17614
rect 15820 17266 15876 17276
rect 14700 16942 14702 16994
rect 14754 16942 14756 16994
rect 14700 16930 14756 16942
rect 14028 16882 14196 16884
rect 14028 16830 14030 16882
rect 14082 16830 14196 16882
rect 14028 16828 14196 16830
rect 14028 16818 14084 16828
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 16604 15428 16660 15438
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 16604 14642 16660 15372
rect 16604 14590 16606 14642
rect 16658 14590 16660 14642
rect 16604 14578 16660 14590
rect 15932 14530 15988 14542
rect 15932 14478 15934 14530
rect 15986 14478 15988 14530
rect 15932 14308 15988 14478
rect 16044 14308 16100 14318
rect 15932 14252 16044 14308
rect 16044 14242 16100 14252
rect 16716 14308 16772 18396
rect 16828 17666 16884 17678
rect 16828 17614 16830 17666
rect 16882 17614 16884 17666
rect 16828 17556 16884 17614
rect 16940 17666 16996 18508
rect 17052 18340 17108 19180
rect 17500 18900 17556 18910
rect 17500 18674 17556 18844
rect 17500 18622 17502 18674
rect 17554 18622 17556 18674
rect 17500 18610 17556 18622
rect 17612 18562 17668 20300
rect 17612 18510 17614 18562
rect 17666 18510 17668 18562
rect 17612 18498 17668 18510
rect 17052 18274 17108 18284
rect 17276 18450 17332 18462
rect 17276 18398 17278 18450
rect 17330 18398 17332 18450
rect 16940 17614 16942 17666
rect 16994 17614 16996 17666
rect 16940 17602 16996 17614
rect 17164 17668 17220 17678
rect 17276 17668 17332 18398
rect 17164 17666 17332 17668
rect 17164 17614 17166 17666
rect 17218 17614 17332 17666
rect 17164 17612 17332 17614
rect 17500 18452 17556 18462
rect 17164 17602 17220 17612
rect 16828 17490 16884 17500
rect 17052 17444 17108 17454
rect 17052 17350 17108 17388
rect 17276 17444 17332 17454
rect 17276 17350 17332 17388
rect 17500 17106 17556 18396
rect 17724 18228 17780 20524
rect 17724 18162 17780 18172
rect 18060 20244 18116 20254
rect 18060 18450 18116 20188
rect 18284 20020 18340 20030
rect 18284 19234 18340 19964
rect 18284 19182 18286 19234
rect 18338 19182 18340 19234
rect 18284 19012 18340 19182
rect 18396 19236 18452 20524
rect 18508 20580 18564 20590
rect 18508 20486 18564 20524
rect 18396 19170 18452 19180
rect 18508 20356 18564 20366
rect 18508 19122 18564 20300
rect 18956 20020 19012 21084
rect 19292 21028 19348 21038
rect 19292 20914 19348 20972
rect 19292 20862 19294 20914
rect 19346 20862 19348 20914
rect 19068 20802 19124 20814
rect 19068 20750 19070 20802
rect 19122 20750 19124 20802
rect 19068 20244 19124 20750
rect 19292 20468 19348 20862
rect 19292 20402 19348 20412
rect 19068 20178 19124 20188
rect 19404 20132 19460 21308
rect 19740 20914 19796 21756
rect 20524 21700 20580 21710
rect 19740 20862 19742 20914
rect 19794 20862 19796 20914
rect 19740 20850 19796 20862
rect 20412 21476 20468 21486
rect 19852 20804 19908 20814
rect 19852 20710 19908 20748
rect 19628 20692 19684 20702
rect 18956 19954 19012 19964
rect 19292 20130 19460 20132
rect 19292 20078 19406 20130
rect 19458 20078 19460 20130
rect 19292 20076 19460 20078
rect 18732 19348 18788 19358
rect 18508 19070 18510 19122
rect 18562 19070 18564 19122
rect 18508 19058 18564 19070
rect 18620 19292 18732 19348
rect 18284 18946 18340 18956
rect 18620 18564 18676 19292
rect 18732 19282 18788 19292
rect 18844 19236 18900 19246
rect 18844 19142 18900 19180
rect 19180 19010 19236 19022
rect 19180 18958 19182 19010
rect 19234 18958 19236 19010
rect 19180 18900 19236 18958
rect 19180 18834 19236 18844
rect 19292 18676 19348 20076
rect 19404 20066 19460 20076
rect 19516 20636 19628 20692
rect 19516 20356 19572 20636
rect 19628 20626 19684 20636
rect 19404 19796 19460 19806
rect 19404 18788 19460 19740
rect 19404 18722 19460 18732
rect 19292 18610 19348 18620
rect 18620 18470 18676 18508
rect 19068 18564 19124 18574
rect 18060 18398 18062 18450
rect 18114 18398 18116 18450
rect 17948 17668 18004 17678
rect 18060 17668 18116 18398
rect 18284 18450 18340 18462
rect 18284 18398 18286 18450
rect 18338 18398 18340 18450
rect 17948 17666 18116 17668
rect 17948 17614 17950 17666
rect 18002 17614 18116 17666
rect 17948 17612 18116 17614
rect 18172 18338 18228 18350
rect 18172 18286 18174 18338
rect 18226 18286 18228 18338
rect 17948 17602 18004 17612
rect 17612 17556 17668 17566
rect 17612 17462 17668 17500
rect 17500 17054 17502 17106
rect 17554 17054 17556 17106
rect 17500 17042 17556 17054
rect 17836 17442 17892 17454
rect 17836 17390 17838 17442
rect 17890 17390 17892 17442
rect 16828 16772 16884 16782
rect 17836 16772 17892 17390
rect 16828 16770 17892 16772
rect 16828 16718 16830 16770
rect 16882 16718 17892 16770
rect 16828 16716 17892 16718
rect 16828 16706 16884 16716
rect 17724 16548 17780 16558
rect 17388 15428 17444 15438
rect 17388 15334 17444 15372
rect 17724 15426 17780 16492
rect 17724 15374 17726 15426
rect 17778 15374 17780 15426
rect 17724 15362 17780 15374
rect 16716 14242 16772 14252
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 17836 8428 17892 16716
rect 18172 17444 18228 18286
rect 18284 18340 18340 18398
rect 19068 18450 19124 18508
rect 19516 18562 19572 20300
rect 19516 18510 19518 18562
rect 19570 18510 19572 18562
rect 19068 18398 19070 18450
rect 19122 18398 19124 18450
rect 19068 18386 19124 18398
rect 19180 18450 19236 18462
rect 19404 18452 19460 18462
rect 19180 18398 19182 18450
rect 19234 18398 19236 18450
rect 18284 18274 18340 18284
rect 19180 18340 19236 18398
rect 19180 18274 19236 18284
rect 19292 18450 19460 18452
rect 19292 18398 19406 18450
rect 19458 18398 19460 18450
rect 19292 18396 19460 18398
rect 18172 16322 18228 17388
rect 18844 18228 18900 18238
rect 18844 17668 18900 18172
rect 19292 18004 19348 18396
rect 19404 18386 19460 18396
rect 19292 17938 19348 17948
rect 19404 18228 19460 18238
rect 18732 17106 18788 17118
rect 18732 17054 18734 17106
rect 18786 17054 18788 17106
rect 18732 16884 18788 17054
rect 18732 16818 18788 16828
rect 18844 16770 18900 17612
rect 19404 17554 19460 18172
rect 19404 17502 19406 17554
rect 19458 17502 19460 17554
rect 19404 17490 19460 17502
rect 19180 17444 19236 17454
rect 18844 16718 18846 16770
rect 18898 16718 18900 16770
rect 18844 16706 18900 16718
rect 19068 17332 19124 17342
rect 19068 17108 19124 17276
rect 19068 16770 19124 17052
rect 19068 16718 19070 16770
rect 19122 16718 19124 16770
rect 19068 16706 19124 16718
rect 18732 16660 18788 16670
rect 18172 16270 18174 16322
rect 18226 16270 18228 16322
rect 18172 16258 18228 16270
rect 18508 16658 18788 16660
rect 18508 16606 18734 16658
rect 18786 16606 18788 16658
rect 18508 16604 18788 16606
rect 18508 16322 18564 16604
rect 18732 16594 18788 16604
rect 18508 16270 18510 16322
rect 18562 16270 18564 16322
rect 18508 16258 18564 16270
rect 19180 16322 19236 17388
rect 19292 16660 19348 16670
rect 19292 16566 19348 16604
rect 19516 16548 19572 18510
rect 19628 20468 19684 20478
rect 19628 19124 19684 20412
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 20300 20244 20356 20254
rect 19628 17666 19684 19068
rect 19964 19348 20020 19358
rect 19964 19124 20020 19292
rect 20300 19236 20356 20188
rect 20300 19142 20356 19180
rect 19964 19122 20244 19124
rect 19964 19070 19966 19122
rect 20018 19070 20244 19122
rect 19964 19068 20244 19070
rect 19964 19058 20020 19068
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 19628 17614 19630 17666
rect 19682 17614 19684 17666
rect 19628 17602 19684 17614
rect 19740 18564 19796 18574
rect 19740 17444 19796 18508
rect 19852 18452 19908 18462
rect 19852 18358 19908 18396
rect 20188 17892 20244 19068
rect 20412 18564 20468 21420
rect 20524 20914 20580 21644
rect 20524 20862 20526 20914
rect 20578 20862 20580 20914
rect 20524 20850 20580 20862
rect 20636 20804 20692 22316
rect 21308 22372 21364 22382
rect 21420 22372 21476 22990
rect 21532 23044 21588 24556
rect 21756 24546 21812 24556
rect 22652 24612 22708 24622
rect 22540 24164 22596 24174
rect 21644 23940 21700 23950
rect 21644 23938 21812 23940
rect 21644 23886 21646 23938
rect 21698 23886 21812 23938
rect 21644 23884 21812 23886
rect 21644 23874 21700 23884
rect 21756 23156 21812 23884
rect 22540 23938 22596 24108
rect 22652 24050 22708 24556
rect 22652 23998 22654 24050
rect 22706 23998 22708 24050
rect 22652 23986 22708 23998
rect 23436 24164 23492 24174
rect 22540 23886 22542 23938
rect 22594 23886 22596 23938
rect 22540 23874 22596 23886
rect 23212 23938 23268 23950
rect 23212 23886 23214 23938
rect 23266 23886 23268 23938
rect 23212 23828 23268 23886
rect 23212 23762 23268 23772
rect 22764 23716 22820 23726
rect 22652 23714 22820 23716
rect 22652 23662 22766 23714
rect 22818 23662 22820 23714
rect 22652 23660 22820 23662
rect 23436 23716 23492 24108
rect 23548 23938 23604 24668
rect 24668 24724 24724 27804
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 40236 27186 40292 27198
rect 40236 27134 40238 27186
rect 40290 27134 40292 27186
rect 40236 26292 40292 27134
rect 40236 26226 40292 26236
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 24668 24630 24724 24668
rect 25340 24724 25396 24734
rect 23884 24612 23940 24622
rect 23884 24518 23940 24556
rect 23548 23886 23550 23938
rect 23602 23886 23604 23938
rect 23548 23874 23604 23886
rect 24220 23828 24276 23838
rect 23660 23826 24276 23828
rect 23660 23774 24222 23826
rect 24274 23774 24276 23826
rect 23660 23772 24276 23774
rect 23436 23660 23604 23716
rect 22540 23380 22596 23390
rect 22652 23380 22708 23660
rect 22764 23650 22820 23660
rect 22540 23378 22708 23380
rect 22540 23326 22542 23378
rect 22594 23326 22708 23378
rect 22540 23324 22708 23326
rect 22540 23314 22596 23324
rect 22204 23156 22260 23166
rect 21756 23154 22204 23156
rect 21756 23102 21758 23154
rect 21810 23102 22204 23154
rect 21756 23100 22204 23102
rect 21644 23044 21700 23054
rect 21532 22988 21644 23044
rect 21644 22978 21700 22988
rect 21420 22316 21588 22372
rect 21308 22278 21364 22316
rect 21532 22148 21588 22316
rect 21756 22370 21812 23100
rect 22204 23062 22260 23100
rect 21756 22318 21758 22370
rect 21810 22318 21812 22370
rect 21756 22306 21812 22318
rect 22428 22370 22484 22382
rect 22428 22318 22430 22370
rect 22482 22318 22484 22370
rect 22092 22258 22148 22270
rect 22092 22206 22094 22258
rect 22146 22206 22148 22258
rect 21588 22092 21700 22148
rect 21532 22082 21588 22092
rect 20636 20738 20692 20748
rect 21532 20804 21588 20814
rect 21532 20710 21588 20748
rect 21308 20692 21364 20702
rect 21308 20598 21364 20636
rect 21532 20356 21588 20366
rect 21196 19234 21252 19246
rect 21196 19182 21198 19234
rect 21250 19182 21252 19234
rect 21196 19124 21252 19182
rect 21532 19234 21588 20300
rect 21532 19182 21534 19234
rect 21586 19182 21588 19234
rect 21532 19170 21588 19182
rect 21644 19124 21700 22092
rect 21868 21028 21924 21038
rect 21868 21026 22036 21028
rect 21868 20974 21870 21026
rect 21922 20974 22036 21026
rect 21868 20972 22036 20974
rect 21868 20962 21924 20972
rect 21868 20804 21924 20814
rect 21868 20710 21924 20748
rect 21756 20580 21812 20590
rect 21756 20486 21812 20524
rect 21868 20020 21924 20030
rect 21756 19460 21812 19470
rect 21756 19346 21812 19404
rect 21756 19294 21758 19346
rect 21810 19294 21812 19346
rect 21756 19282 21812 19294
rect 21756 19124 21812 19134
rect 21644 19122 21812 19124
rect 21644 19070 21758 19122
rect 21810 19070 21812 19122
rect 21644 19068 21812 19070
rect 21196 19058 21252 19068
rect 21756 19058 21812 19068
rect 20748 18676 20804 18686
rect 20524 18564 20580 18574
rect 20412 18562 20580 18564
rect 20412 18510 20526 18562
rect 20578 18510 20580 18562
rect 20412 18508 20580 18510
rect 20524 18498 20580 18508
rect 20188 17836 20356 17892
rect 20188 17668 20244 17678
rect 20188 17574 20244 17612
rect 19964 17556 20020 17566
rect 19964 17462 20020 17500
rect 19740 17378 19796 17388
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 20300 17108 20356 17836
rect 20748 17666 20804 18620
rect 21644 18564 21700 18574
rect 21644 18452 21700 18508
rect 21868 18452 21924 19964
rect 21980 18676 22036 20972
rect 22092 20132 22148 22206
rect 22092 19796 22148 20076
rect 22428 20578 22484 22318
rect 22428 20526 22430 20578
rect 22482 20526 22484 20578
rect 22428 19796 22484 20526
rect 22540 20804 22596 20814
rect 22540 20018 22596 20748
rect 22540 19966 22542 20018
rect 22594 19966 22596 20018
rect 22540 19954 22596 19966
rect 22540 19796 22596 19806
rect 22428 19740 22540 19796
rect 22092 19730 22148 19740
rect 22540 19730 22596 19740
rect 22428 19124 22484 19134
rect 22428 19122 22596 19124
rect 22428 19070 22430 19122
rect 22482 19070 22596 19122
rect 22428 19068 22596 19070
rect 22428 19058 22484 19068
rect 22092 19010 22148 19022
rect 22092 18958 22094 19010
rect 22146 18958 22148 19010
rect 22092 18900 22148 18958
rect 22540 19012 22596 19068
rect 22092 18844 22484 18900
rect 21980 18610 22036 18620
rect 21644 18396 21924 18452
rect 22092 18564 22148 18574
rect 22092 18450 22148 18508
rect 22428 18452 22484 18844
rect 22540 18562 22596 18956
rect 22540 18510 22542 18562
rect 22594 18510 22596 18562
rect 22540 18498 22596 18510
rect 22092 18398 22094 18450
rect 22146 18398 22148 18450
rect 21644 17778 21700 18396
rect 22092 18386 22148 18398
rect 22316 18396 22428 18452
rect 21644 17726 21646 17778
rect 21698 17726 21700 17778
rect 21644 17714 21700 17726
rect 20748 17614 20750 17666
rect 20802 17614 20804 17666
rect 20748 17602 20804 17614
rect 21868 17668 21924 17678
rect 21868 17574 21924 17612
rect 20188 17052 20356 17108
rect 21420 17554 21476 17566
rect 21420 17502 21422 17554
rect 21474 17502 21476 17554
rect 21420 17108 21476 17502
rect 22092 17556 22148 17566
rect 22092 17462 22148 17500
rect 20076 16772 20132 16782
rect 20188 16772 20244 17052
rect 21420 17042 21476 17052
rect 21756 17444 21812 17454
rect 20300 16884 20356 16894
rect 21420 16884 21476 16894
rect 20300 16882 20468 16884
rect 20300 16830 20302 16882
rect 20354 16830 20468 16882
rect 20300 16828 20468 16830
rect 20300 16818 20356 16828
rect 19964 16770 20244 16772
rect 19964 16718 20078 16770
rect 20130 16718 20244 16770
rect 19964 16716 20244 16718
rect 19740 16660 19796 16670
rect 19740 16566 19796 16604
rect 19852 16658 19908 16670
rect 19852 16606 19854 16658
rect 19906 16606 19908 16658
rect 19404 16492 19572 16548
rect 19852 16548 19908 16606
rect 19404 16436 19460 16492
rect 19852 16482 19908 16492
rect 19180 16270 19182 16322
rect 19234 16270 19236 16322
rect 19180 16258 19236 16270
rect 19292 16324 19348 16334
rect 19404 16324 19460 16380
rect 19292 16322 19460 16324
rect 19292 16270 19294 16322
rect 19346 16270 19460 16322
rect 19292 16268 19460 16270
rect 19516 16324 19572 16334
rect 19964 16324 20020 16716
rect 20076 16706 20132 16716
rect 20300 16660 20356 16670
rect 20188 16548 20244 16558
rect 19516 16322 20020 16324
rect 19516 16270 19518 16322
rect 19570 16270 20020 16322
rect 19516 16268 20020 16270
rect 20076 16492 20188 16548
rect 20076 16322 20132 16492
rect 20188 16482 20244 16492
rect 20076 16270 20078 16322
rect 20130 16270 20132 16322
rect 19292 16258 19348 16268
rect 19516 16258 19572 16268
rect 20076 16258 20132 16270
rect 20300 16322 20356 16604
rect 20412 16436 20468 16828
rect 21420 16790 21476 16828
rect 20412 16370 20468 16380
rect 20300 16270 20302 16322
rect 20354 16270 20356 16322
rect 20300 16258 20356 16270
rect 21756 16322 21812 17388
rect 21980 17442 22036 17454
rect 21980 17390 21982 17442
rect 22034 17390 22036 17442
rect 21980 16996 22036 17390
rect 22092 16996 22148 17006
rect 21980 16994 22148 16996
rect 21980 16942 22094 16994
rect 22146 16942 22148 16994
rect 21980 16940 22148 16942
rect 22092 16930 22148 16940
rect 22316 16996 22372 18396
rect 22428 18386 22484 18396
rect 22652 17780 22708 23324
rect 23548 23378 23604 23660
rect 23548 23326 23550 23378
rect 23602 23326 23604 23378
rect 23548 23314 23604 23326
rect 23660 23378 23716 23772
rect 24220 23762 24276 23772
rect 23660 23326 23662 23378
rect 23714 23326 23716 23378
rect 23660 23314 23716 23326
rect 22876 23156 22932 23166
rect 22876 23062 22932 23100
rect 22988 23154 23044 23166
rect 22988 23102 22990 23154
rect 23042 23102 23044 23154
rect 22988 23044 23044 23102
rect 23772 23156 23828 23166
rect 23772 23154 23940 23156
rect 23772 23102 23774 23154
rect 23826 23102 23940 23154
rect 23772 23100 23940 23102
rect 23772 23090 23828 23100
rect 22988 22370 23044 22988
rect 22988 22318 22990 22370
rect 23042 22318 23044 22370
rect 22988 22306 23044 22318
rect 23660 22370 23716 22382
rect 23660 22318 23662 22370
rect 23714 22318 23716 22370
rect 23324 21474 23380 21486
rect 23324 21422 23326 21474
rect 23378 21422 23380 21474
rect 22764 20916 22820 20926
rect 22764 20690 22820 20860
rect 23324 20804 23380 21422
rect 23324 20710 23380 20748
rect 22764 20638 22766 20690
rect 22818 20638 22820 20690
rect 22764 20626 22820 20638
rect 23660 20356 23716 22318
rect 23660 20290 23716 20300
rect 23100 20132 23156 20142
rect 23100 20038 23156 20076
rect 23324 20132 23380 20142
rect 23884 20132 23940 23100
rect 24220 23154 24276 23166
rect 24220 23102 24222 23154
rect 24274 23102 24276 23154
rect 24220 22482 24276 23102
rect 24220 22430 24222 22482
rect 24274 22430 24276 22482
rect 24220 22418 24276 22430
rect 24220 22260 24276 22270
rect 24220 22166 24276 22204
rect 23996 22146 24052 22158
rect 23996 22094 23998 22146
rect 24050 22094 24052 22146
rect 23996 20916 24052 22094
rect 25340 21586 25396 24668
rect 26572 24724 26628 24734
rect 26348 24050 26404 24062
rect 26348 23998 26350 24050
rect 26402 23998 26404 24050
rect 26348 23604 26404 23998
rect 26348 22260 26404 23548
rect 26572 23380 26628 24668
rect 37884 24722 37940 24734
rect 37884 24670 37886 24722
rect 37938 24670 37940 24722
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 28140 24164 28196 24174
rect 27804 24162 28196 24164
rect 27804 24110 28142 24162
rect 28194 24110 28196 24162
rect 27804 24108 28196 24110
rect 27356 24052 27412 24062
rect 27356 23938 27412 23996
rect 27356 23886 27358 23938
rect 27410 23886 27412 23938
rect 27356 23874 27412 23886
rect 26684 23714 26740 23726
rect 26684 23662 26686 23714
rect 26738 23662 26740 23714
rect 26684 23604 26740 23662
rect 27020 23716 27076 23726
rect 27020 23622 27076 23660
rect 27692 23714 27748 23726
rect 27692 23662 27694 23714
rect 27746 23662 27748 23714
rect 26684 23538 26740 23548
rect 27692 23492 27748 23662
rect 27692 23426 27748 23436
rect 26572 23378 26964 23380
rect 26572 23326 26574 23378
rect 26626 23326 26964 23378
rect 26572 23324 26964 23326
rect 26572 23314 26628 23324
rect 26908 23156 26964 23324
rect 27692 23268 27748 23278
rect 27804 23268 27860 24108
rect 28140 24098 28196 24108
rect 37660 23940 37716 23950
rect 37660 23846 37716 23884
rect 28028 23828 28084 23838
rect 28028 23734 28084 23772
rect 28140 23714 28196 23726
rect 28140 23662 28142 23714
rect 28194 23662 28196 23714
rect 28140 23380 28196 23662
rect 37884 23604 37940 24670
rect 40012 24498 40068 24510
rect 40012 24446 40014 24498
rect 40066 24446 40068 24498
rect 40012 24276 40068 24446
rect 40012 24210 40068 24220
rect 37884 23538 37940 23548
rect 40012 24050 40068 24062
rect 40012 23998 40014 24050
rect 40066 23998 40068 24050
rect 40012 23604 40068 23998
rect 40012 23538 40068 23548
rect 29372 23492 29428 23502
rect 28140 23314 28196 23324
rect 29036 23380 29092 23390
rect 27692 23266 27860 23268
rect 27692 23214 27694 23266
rect 27746 23214 27860 23266
rect 27692 23212 27860 23214
rect 27692 23202 27748 23212
rect 26908 23062 26964 23100
rect 28140 23156 28196 23166
rect 28140 22484 28196 23100
rect 28588 22484 28644 22494
rect 26348 22194 26404 22204
rect 27692 22482 28644 22484
rect 27692 22430 28142 22482
rect 28194 22430 28590 22482
rect 28642 22430 28644 22482
rect 27692 22428 28644 22430
rect 25340 21534 25342 21586
rect 25394 21534 25396 21586
rect 23996 20850 24052 20860
rect 25116 20916 25172 20926
rect 25172 20860 25284 20916
rect 25116 20850 25172 20860
rect 23324 20130 23940 20132
rect 23324 20078 23326 20130
rect 23378 20078 23940 20130
rect 23324 20076 23940 20078
rect 23324 20066 23380 20076
rect 22988 20020 23044 20030
rect 22988 19926 23044 19964
rect 23884 20018 23940 20076
rect 23884 19966 23886 20018
rect 23938 19966 23940 20018
rect 23884 19954 23940 19966
rect 23996 20468 24052 20478
rect 22764 19796 22820 19806
rect 22764 19236 22820 19740
rect 23996 19348 24052 20412
rect 24668 20468 24724 20478
rect 24556 20244 24612 20254
rect 24556 20150 24612 20188
rect 24332 20130 24388 20142
rect 24332 20078 24334 20130
rect 24386 20078 24388 20130
rect 24332 20020 24388 20078
rect 24444 20132 24500 20142
rect 24444 20038 24500 20076
rect 24668 20130 24724 20412
rect 24668 20078 24670 20130
rect 24722 20078 24724 20130
rect 24668 20066 24724 20078
rect 25228 20130 25284 20860
rect 25340 20914 25396 21534
rect 25340 20862 25342 20914
rect 25394 20862 25396 20914
rect 25340 20850 25396 20862
rect 26012 21474 26068 21486
rect 26012 21422 26014 21474
rect 26066 21422 26068 21474
rect 26012 20244 26068 21422
rect 26908 21476 26964 21486
rect 26908 20188 26964 21420
rect 26012 20178 26068 20188
rect 25228 20078 25230 20130
rect 25282 20078 25284 20130
rect 25228 20066 25284 20078
rect 26236 20130 26292 20142
rect 26236 20078 26238 20130
rect 26290 20078 26292 20130
rect 24332 19954 24388 19964
rect 25564 20018 25620 20030
rect 25564 19966 25566 20018
rect 25618 19966 25620 20018
rect 25340 19908 25396 19918
rect 25340 19906 25508 19908
rect 25340 19854 25342 19906
rect 25394 19854 25508 19906
rect 25340 19852 25508 19854
rect 25340 19842 25396 19852
rect 22764 18564 22820 19180
rect 23660 19292 24052 19348
rect 23436 18676 23492 18686
rect 23436 18582 23492 18620
rect 22764 18498 22820 18508
rect 22988 17892 23044 17902
rect 22988 17798 23044 17836
rect 23660 17890 23716 19292
rect 23660 17838 23662 17890
rect 23714 17838 23716 17890
rect 23660 17826 23716 17838
rect 24332 19234 24388 19246
rect 24332 19182 24334 19234
rect 24386 19182 24388 19234
rect 22764 17780 22820 17790
rect 22428 17778 22820 17780
rect 22428 17726 22766 17778
rect 22818 17726 22820 17778
rect 22428 17724 22820 17726
rect 22428 17666 22484 17724
rect 22764 17714 22820 17724
rect 22428 17614 22430 17666
rect 22482 17614 22484 17666
rect 22428 17444 22484 17614
rect 23772 17668 23828 17678
rect 23772 17574 23828 17612
rect 23996 17668 24052 17678
rect 23996 17666 24164 17668
rect 23996 17614 23998 17666
rect 24050 17614 24164 17666
rect 23996 17612 24164 17614
rect 23996 17602 24052 17612
rect 22428 17378 22484 17388
rect 23324 17444 23380 17454
rect 23324 17350 23380 17388
rect 22316 16930 22372 16940
rect 21756 16270 21758 16322
rect 21810 16270 21812 16322
rect 21756 16258 21812 16270
rect 23548 16884 23604 16894
rect 21420 16210 21476 16222
rect 21420 16158 21422 16210
rect 21474 16158 21476 16210
rect 18508 16098 18564 16110
rect 18508 16046 18510 16098
rect 18562 16046 18564 16098
rect 18508 15314 18564 16046
rect 19628 16100 19684 16110
rect 19628 16006 19684 16044
rect 20524 16100 20580 16110
rect 20524 16006 20580 16044
rect 20748 16100 20804 16110
rect 21420 16100 21476 16158
rect 20748 16098 21476 16100
rect 20748 16046 20750 16098
rect 20802 16046 21476 16098
rect 20748 16044 21476 16046
rect 20748 16034 20804 16044
rect 20636 15876 20692 15886
rect 20524 15874 20692 15876
rect 20524 15822 20638 15874
rect 20690 15822 20692 15874
rect 20524 15820 20692 15822
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 18508 15262 18510 15314
rect 18562 15262 18564 15314
rect 18508 14756 18564 15262
rect 18732 15426 18788 15438
rect 18732 15374 18734 15426
rect 18786 15374 18788 15426
rect 18732 15148 18788 15374
rect 20188 15426 20244 15438
rect 20188 15374 20190 15426
rect 20242 15374 20244 15426
rect 18732 15092 19124 15148
rect 18956 14756 19012 14766
rect 18508 14754 19012 14756
rect 18508 14702 18958 14754
rect 19010 14702 19012 14754
rect 18508 14700 19012 14702
rect 18732 14642 18788 14700
rect 18956 14690 19012 14700
rect 18732 14590 18734 14642
rect 18786 14590 18788 14642
rect 18732 14578 18788 14590
rect 17724 8372 17892 8428
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 17500 5236 17556 5246
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 17500 800 17556 5180
rect 17724 5122 17780 8372
rect 18732 5236 18788 5246
rect 18732 5142 18788 5180
rect 17724 5070 17726 5122
rect 17778 5070 17780 5122
rect 17724 5058 17780 5070
rect 19068 4338 19124 15092
rect 19292 14756 19348 14766
rect 19292 14754 19684 14756
rect 19292 14702 19294 14754
rect 19346 14702 19684 14754
rect 19292 14700 19684 14702
rect 19292 14690 19348 14700
rect 19180 14308 19236 14318
rect 19180 13748 19236 14252
rect 19404 13748 19460 13758
rect 19180 13692 19404 13748
rect 19404 13654 19460 13692
rect 19068 4286 19070 4338
rect 19122 4286 19124 4338
rect 19068 4274 19124 4286
rect 18844 4116 18900 4126
rect 18172 3666 18228 3678
rect 18172 3614 18174 3666
rect 18226 3614 18228 3666
rect 18172 800 18228 3614
rect 18844 800 18900 4060
rect 19628 3556 19684 14700
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 20076 13860 20132 13870
rect 20188 13860 20244 15374
rect 20524 15426 20580 15820
rect 20636 15810 20692 15820
rect 21532 15874 21588 15886
rect 21532 15822 21534 15874
rect 21586 15822 21588 15874
rect 20524 15374 20526 15426
rect 20578 15374 20580 15426
rect 20524 15362 20580 15374
rect 20076 13858 20244 13860
rect 20076 13806 20078 13858
rect 20130 13806 20244 13858
rect 20076 13804 20244 13806
rect 20076 13794 20132 13804
rect 21420 13524 21476 13534
rect 21532 13524 21588 15822
rect 23548 14530 23604 16828
rect 23548 14478 23550 14530
rect 23602 14478 23604 14530
rect 23548 14466 23604 14478
rect 24108 16772 24164 17612
rect 24332 16884 24388 19182
rect 25116 19122 25172 19134
rect 25116 19070 25118 19122
rect 25170 19070 25172 19122
rect 25116 18340 25172 19070
rect 25340 18562 25396 18574
rect 25340 18510 25342 18562
rect 25394 18510 25396 18562
rect 25340 18452 25396 18510
rect 25452 18564 25508 19852
rect 25564 19348 25620 19966
rect 25564 19282 25620 19292
rect 25676 20018 25732 20030
rect 25676 19966 25678 20018
rect 25730 19966 25732 20018
rect 25676 18676 25732 19966
rect 25676 18610 25732 18620
rect 26124 20018 26180 20030
rect 26124 19966 26126 20018
rect 26178 19966 26180 20018
rect 25564 18564 25620 18574
rect 25452 18562 25620 18564
rect 25452 18510 25566 18562
rect 25618 18510 25620 18562
rect 25452 18508 25620 18510
rect 25564 18498 25620 18508
rect 25228 18340 25284 18350
rect 25116 18338 25284 18340
rect 25116 18286 25230 18338
rect 25282 18286 25284 18338
rect 25116 18284 25284 18286
rect 25228 18274 25284 18284
rect 24332 16818 24388 16828
rect 24444 18116 24500 18126
rect 24220 16772 24276 16782
rect 24108 16770 24276 16772
rect 24108 16718 24222 16770
rect 24274 16718 24276 16770
rect 24108 16716 24276 16718
rect 22652 13748 22708 13758
rect 22652 13654 22708 13692
rect 21476 13468 21588 13524
rect 22204 13634 22260 13646
rect 22204 13582 22206 13634
rect 22258 13582 22260 13634
rect 22204 13524 22260 13582
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 20076 4116 20132 4126
rect 20076 4022 20132 4060
rect 19740 3556 19796 3566
rect 19628 3554 19796 3556
rect 19628 3502 19742 3554
rect 19794 3502 19796 3554
rect 19628 3500 19796 3502
rect 19740 3490 19796 3500
rect 21420 3554 21476 13468
rect 22204 13458 22260 13468
rect 24108 8428 24164 16716
rect 24220 16706 24276 16716
rect 24444 15986 24500 18060
rect 24668 16884 24724 16894
rect 24668 16790 24724 16828
rect 24668 16212 24724 16222
rect 25116 16212 25172 16222
rect 24668 16210 25172 16212
rect 24668 16158 24670 16210
rect 24722 16158 25118 16210
rect 25170 16158 25172 16210
rect 24668 16156 25172 16158
rect 24668 16146 24724 16156
rect 25116 16146 25172 16156
rect 24444 15934 24446 15986
rect 24498 15934 24500 15986
rect 24444 15922 24500 15934
rect 25004 15988 25060 15998
rect 24556 15874 24612 15886
rect 24556 15822 24558 15874
rect 24610 15822 24612 15874
rect 24556 15148 24612 15822
rect 24332 15092 24612 15148
rect 25004 15204 25060 15932
rect 25340 15988 25396 18396
rect 26124 18116 26180 19966
rect 26236 19460 26292 20078
rect 26684 20132 26740 20142
rect 26684 20038 26740 20076
rect 26796 20132 26964 20188
rect 26796 20130 26852 20132
rect 26796 20078 26798 20130
rect 26850 20078 26852 20130
rect 26796 20066 26852 20078
rect 26460 20020 26516 20030
rect 26460 19926 26516 19964
rect 27692 20018 27748 22428
rect 28140 22418 28196 22428
rect 28588 21586 28644 22428
rect 29036 22370 29092 23324
rect 29036 22318 29038 22370
rect 29090 22318 29092 22370
rect 29036 22306 29092 22318
rect 29260 23044 29316 23054
rect 29260 22258 29316 22988
rect 29372 22372 29428 23436
rect 30268 23156 30324 23166
rect 30268 23062 30324 23100
rect 37660 23156 37716 23166
rect 37660 23062 37716 23100
rect 29820 23044 29876 23054
rect 29820 22950 29876 22988
rect 40012 22932 40068 22942
rect 40012 22838 40068 22876
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 40012 22482 40068 22494
rect 40012 22430 40014 22482
rect 40066 22430 40068 22482
rect 29372 22370 29764 22372
rect 29372 22318 29374 22370
rect 29426 22318 29764 22370
rect 29372 22316 29764 22318
rect 29372 22306 29428 22316
rect 29260 22206 29262 22258
rect 29314 22206 29316 22258
rect 29260 22194 29316 22206
rect 28588 21534 28590 21586
rect 28642 21534 28644 21586
rect 28588 21522 28644 21534
rect 28140 21476 28196 21486
rect 28140 21382 28196 21420
rect 29260 21476 29316 21486
rect 29260 21474 29652 21476
rect 29260 21422 29262 21474
rect 29314 21422 29652 21474
rect 29260 21420 29652 21422
rect 29260 21410 29316 21420
rect 29596 20914 29652 21420
rect 29596 20862 29598 20914
rect 29650 20862 29652 20914
rect 29596 20850 29652 20862
rect 29484 20804 29540 20814
rect 29484 20710 29540 20748
rect 29708 20804 29764 22316
rect 37884 22370 37940 22382
rect 37884 22318 37886 22370
rect 37938 22318 37940 22370
rect 37660 21588 37716 21598
rect 37548 21586 37716 21588
rect 37548 21534 37662 21586
rect 37714 21534 37716 21586
rect 37548 21532 37716 21534
rect 31388 21474 31444 21486
rect 31388 21422 31390 21474
rect 31442 21422 31444 21474
rect 30156 20916 30212 20926
rect 30044 20804 30100 20814
rect 29708 20802 30100 20804
rect 29708 20750 29710 20802
rect 29762 20750 30046 20802
rect 30098 20750 30100 20802
rect 29708 20748 30100 20750
rect 29148 20692 29204 20702
rect 29148 20598 29204 20636
rect 27692 19966 27694 20018
rect 27746 19966 27748 20018
rect 27356 19908 27412 19918
rect 27692 19908 27748 19966
rect 27356 19906 27748 19908
rect 27356 19854 27358 19906
rect 27410 19854 27748 19906
rect 27356 19852 27748 19854
rect 27356 19842 27412 19852
rect 26236 19012 26292 19404
rect 27244 19348 27300 19358
rect 27244 19254 27300 19292
rect 26236 18946 26292 18956
rect 27692 19010 27748 19852
rect 28252 20580 28308 20590
rect 28252 19236 28308 20524
rect 28476 19906 28532 19918
rect 28476 19854 28478 19906
rect 28530 19854 28532 19906
rect 28364 19460 28420 19470
rect 28476 19460 28532 19854
rect 28364 19458 28532 19460
rect 28364 19406 28366 19458
rect 28418 19406 28532 19458
rect 28364 19404 28532 19406
rect 28364 19394 28420 19404
rect 28476 19236 28532 19246
rect 28252 19234 28532 19236
rect 28252 19182 28478 19234
rect 28530 19182 28532 19234
rect 28252 19180 28532 19182
rect 28476 19170 28532 19180
rect 27692 18958 27694 19010
rect 27746 18958 27748 19010
rect 26124 18050 26180 18060
rect 27356 17554 27412 17566
rect 27356 17502 27358 17554
rect 27410 17502 27412 17554
rect 26572 17444 26628 17454
rect 27356 17444 27412 17502
rect 27580 17556 27636 17566
rect 27580 17462 27636 17500
rect 26628 17388 26740 17444
rect 26572 17378 26628 17388
rect 25676 16884 25732 16894
rect 25676 16098 25732 16828
rect 25676 16046 25678 16098
rect 25730 16046 25732 16098
rect 25676 16034 25732 16046
rect 25340 15922 25396 15932
rect 26460 15988 26516 15998
rect 26460 15986 26628 15988
rect 26460 15934 26462 15986
rect 26514 15934 26628 15986
rect 26460 15932 26628 15934
rect 26460 15922 26516 15932
rect 25004 15138 25060 15148
rect 25228 15874 25284 15886
rect 25228 15822 25230 15874
rect 25282 15822 25284 15874
rect 25228 15148 25284 15822
rect 26572 15202 26628 15932
rect 26684 15538 26740 17388
rect 27356 17378 27412 17388
rect 26908 16884 26964 16894
rect 27244 16884 27300 16894
rect 27692 16884 27748 18958
rect 28364 19012 28420 19022
rect 28364 18918 28420 18956
rect 28252 18788 28308 18798
rect 27916 17780 27972 17790
rect 27916 17778 28084 17780
rect 27916 17726 27918 17778
rect 27970 17726 28084 17778
rect 27916 17724 28084 17726
rect 27916 17714 27972 17724
rect 27804 17668 27860 17706
rect 27804 17602 27860 17612
rect 27916 17556 27972 17566
rect 27916 17462 27972 17500
rect 28028 16994 28084 17724
rect 28252 17556 28308 18732
rect 29708 18788 29764 20748
rect 30044 20738 30100 20748
rect 30156 20690 30212 20860
rect 30828 20916 30884 20926
rect 30604 20804 30660 20814
rect 30604 20710 30660 20748
rect 30156 20638 30158 20690
rect 30210 20638 30212 20690
rect 30156 20626 30212 20638
rect 30716 20692 30772 20702
rect 30716 20598 30772 20636
rect 30380 20580 30436 20590
rect 30380 20486 30436 20524
rect 30828 20188 30884 20860
rect 31388 20692 31444 21422
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 31388 20626 31444 20636
rect 37548 20692 37604 21532
rect 37660 21522 37716 21532
rect 37884 21476 37940 22318
rect 40012 21588 40068 22430
rect 40012 21522 40068 21532
rect 37884 21410 37940 21420
rect 39900 21474 39956 21486
rect 39900 21422 39902 21474
rect 39954 21422 39956 21474
rect 39900 20916 39956 21422
rect 39900 20850 39956 20860
rect 40012 20914 40068 20926
rect 40012 20862 40014 20914
rect 40066 20862 40068 20914
rect 37660 20804 37716 20814
rect 37660 20710 37716 20748
rect 37548 20626 37604 20636
rect 30604 20132 30884 20188
rect 40012 20244 40068 20862
rect 40012 20178 40068 20188
rect 30604 19906 30660 20132
rect 30604 19854 30606 19906
rect 30658 19854 30660 19906
rect 30604 19842 30660 19854
rect 37660 20018 37716 20030
rect 37660 19966 37662 20018
rect 37714 19966 37716 20018
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 37660 19348 37716 19966
rect 40012 19794 40068 19806
rect 40012 19742 40014 19794
rect 40066 19742 40068 19794
rect 40012 19572 40068 19742
rect 40012 19506 40068 19516
rect 37660 19282 37716 19292
rect 29708 18722 29764 18732
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 40012 17778 40068 17790
rect 40012 17726 40014 17778
rect 40066 17726 40068 17778
rect 29148 17668 29204 17678
rect 29148 17574 29204 17612
rect 37660 17668 37716 17678
rect 37660 17574 37716 17612
rect 28252 17490 28308 17500
rect 29260 17556 29316 17566
rect 29260 17462 29316 17500
rect 30156 17556 30212 17566
rect 28028 16942 28030 16994
rect 28082 16942 28084 16994
rect 28028 16930 28084 16942
rect 26908 16882 27748 16884
rect 26908 16830 26910 16882
rect 26962 16830 27246 16882
rect 27298 16830 27748 16882
rect 26908 16828 27748 16830
rect 26908 16772 26964 16828
rect 27244 16818 27300 16828
rect 26684 15486 26686 15538
rect 26738 15486 26740 15538
rect 26684 15474 26740 15486
rect 26796 16716 26908 16772
rect 26796 16212 26852 16716
rect 26908 16706 26964 16716
rect 28588 16772 28644 16782
rect 26572 15150 26574 15202
rect 26626 15150 26628 15202
rect 25228 15092 25396 15148
rect 26572 15138 26628 15150
rect 24220 14644 24276 14654
rect 24332 14644 24388 15092
rect 24220 14642 24388 14644
rect 24220 14590 24222 14642
rect 24274 14590 24388 14642
rect 24220 14588 24388 14590
rect 25340 14644 25396 15092
rect 26796 15092 26852 16156
rect 28588 16210 28644 16716
rect 30156 16770 30212 17500
rect 40012 17556 40068 17726
rect 40012 17490 40068 17500
rect 30156 16718 30158 16770
rect 30210 16718 30212 16770
rect 30156 16706 30212 16718
rect 37660 16882 37716 16894
rect 37660 16830 37662 16882
rect 37714 16830 37716 16882
rect 37660 16772 37716 16830
rect 37660 16706 37716 16716
rect 40012 16658 40068 16670
rect 40012 16606 40014 16658
rect 40066 16606 40068 16658
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 28588 16158 28590 16210
rect 28642 16158 28644 16210
rect 27580 15540 27636 15550
rect 26908 15316 26964 15326
rect 27356 15316 27412 15326
rect 26908 15314 27412 15316
rect 26908 15262 26910 15314
rect 26962 15262 27358 15314
rect 27410 15262 27412 15314
rect 26908 15260 27412 15262
rect 26908 15250 26964 15260
rect 27356 15250 27412 15260
rect 27580 15314 27636 15484
rect 28588 15540 28644 16158
rect 29260 16212 29316 16222
rect 29260 16118 29316 16156
rect 40012 16212 40068 16606
rect 40012 16146 40068 16156
rect 28588 15474 28644 15484
rect 27580 15262 27582 15314
rect 27634 15262 27636 15314
rect 27580 15250 27636 15262
rect 27244 15092 27300 15102
rect 26796 15036 26964 15092
rect 26348 14644 26404 14654
rect 25340 14642 26404 14644
rect 25340 14590 26350 14642
rect 26402 14590 26404 14642
rect 25340 14588 26404 14590
rect 24220 14578 24276 14588
rect 26348 8428 26404 14588
rect 26908 14642 26964 15036
rect 27244 14998 27300 15036
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 26908 14590 26910 14642
rect 26962 14590 26964 14642
rect 26908 14578 26964 14590
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 24108 8372 24612 8428
rect 24444 4452 24500 4462
rect 24220 4450 24500 4452
rect 24220 4398 24446 4450
rect 24498 4398 24500 4450
rect 24220 4396 24500 4398
rect 21420 3502 21422 3554
rect 21474 3502 21476 3554
rect 21420 3490 21476 3502
rect 23548 3668 23604 3678
rect 22428 3332 22484 3342
rect 22204 3330 22484 3332
rect 22204 3278 22430 3330
rect 22482 3278 22484 3330
rect 22204 3276 22484 3278
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 22204 800 22260 3276
rect 22428 3266 22484 3276
rect 23548 800 23604 3612
rect 24220 800 24276 4396
rect 24444 4386 24500 4396
rect 24556 3554 24612 8372
rect 25788 8372 26404 8428
rect 25788 4338 25844 8372
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 25788 4286 25790 4338
rect 25842 4286 25844 4338
rect 25788 4274 25844 4286
rect 26796 4114 26852 4126
rect 26796 4062 26798 4114
rect 26850 4062 26852 4114
rect 25564 3668 25620 3678
rect 25564 3574 25620 3612
rect 24556 3502 24558 3554
rect 24610 3502 24612 3554
rect 24556 3490 24612 3502
rect 25564 3444 25620 3454
rect 25564 800 25620 3388
rect 26796 3444 26852 4062
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 26796 3378 26852 3388
rect 17472 0 17584 800
rect 18144 0 18256 800
rect 18816 0 18928 800
rect 22176 0 22288 800
rect 23520 0 23632 800
rect 24192 0 24304 800
rect 25536 0 25648 800
<< via2 >>
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 4172 27580 4228 27636
rect 1932 26236 1988 26292
rect 2044 26908 2100 26964
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 4284 27074 4340 27076
rect 4284 27022 4286 27074
rect 4286 27022 4338 27074
rect 4338 27022 4340 27074
rect 4284 27020 4340 27022
rect 11452 26908 11508 26964
rect 13468 26684 13524 26740
rect 4284 26290 4340 26292
rect 4284 26238 4286 26290
rect 4286 26238 4338 26290
rect 4338 26238 4340 26290
rect 4284 26236 4340 26238
rect 11788 26236 11844 26292
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 14364 26908 14420 26964
rect 17724 26962 17780 26964
rect 17724 26910 17726 26962
rect 17726 26910 17778 26962
rect 17778 26910 17780 26962
rect 17724 26908 17780 26910
rect 17052 26796 17108 26852
rect 18732 27804 18788 27860
rect 17836 26796 17892 26852
rect 14924 26460 14980 26516
rect 15372 26684 15428 26740
rect 15596 26460 15652 26516
rect 14588 25676 14644 25732
rect 15260 26290 15316 26292
rect 15260 26238 15262 26290
rect 15262 26238 15314 26290
rect 15314 26238 15316 26290
rect 15260 26236 15316 26238
rect 15036 25676 15092 25732
rect 14028 25340 14084 25396
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 13468 24162 13524 24164
rect 13468 24110 13470 24162
rect 13470 24110 13522 24162
rect 13522 24110 13524 24162
rect 13468 24108 13524 24110
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 4172 21644 4228 21700
rect 4284 21586 4340 21588
rect 4284 21534 4286 21586
rect 4286 21534 4338 21586
rect 4338 21534 4340 21586
rect 4284 21532 4340 21534
rect 9996 21532 10052 21588
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 1932 20860 1988 20916
rect 11564 21586 11620 21588
rect 11564 21534 11566 21586
rect 11566 21534 11618 21586
rect 11618 21534 11620 21586
rect 11564 21532 11620 21534
rect 15372 25340 15428 25396
rect 15484 25564 15540 25620
rect 14252 24050 14308 24052
rect 14252 23998 14254 24050
rect 14254 23998 14306 24050
rect 14306 23998 14308 24050
rect 14252 23996 14308 23998
rect 18620 27020 18676 27076
rect 18732 26908 18788 26964
rect 19292 27858 19348 27860
rect 19292 27806 19294 27858
rect 19294 27806 19346 27858
rect 19346 27806 19348 27858
rect 19292 27804 19348 27806
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 22876 38220 22932 38276
rect 25564 38274 25620 38276
rect 25564 38222 25566 38274
rect 25566 38222 25618 38274
rect 25618 38222 25620 38274
rect 25564 38220 25620 38222
rect 20860 37436 20916 37492
rect 22092 37490 22148 37492
rect 22092 37438 22094 37490
rect 22094 37438 22146 37490
rect 22146 37438 22148 37490
rect 22092 37436 22148 37438
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 18956 26908 19012 26964
rect 17836 25564 17892 25620
rect 18284 25676 18340 25732
rect 16156 24892 16212 24948
rect 16492 25340 16548 25396
rect 15708 23996 15764 24052
rect 17948 25228 18004 25284
rect 17500 24946 17556 24948
rect 17500 24894 17502 24946
rect 17502 24894 17554 24946
rect 17554 24894 17556 24946
rect 17500 24892 17556 24894
rect 16492 24668 16548 24724
rect 14140 23884 14196 23940
rect 15596 23884 15652 23940
rect 14812 22876 14868 22932
rect 14476 22316 14532 22372
rect 12348 22092 12404 22148
rect 13580 22146 13636 22148
rect 13580 22094 13582 22146
rect 13582 22094 13634 22146
rect 13634 22094 13636 22146
rect 13580 22092 13636 22094
rect 14028 22092 14084 22148
rect 12236 21532 12292 21588
rect 12796 21532 12852 21588
rect 14252 21308 14308 21364
rect 12796 20860 12852 20916
rect 12124 20802 12180 20804
rect 12124 20750 12126 20802
rect 12126 20750 12178 20802
rect 12178 20750 12180 20802
rect 12124 20748 12180 20750
rect 13580 20914 13636 20916
rect 13580 20862 13582 20914
rect 13582 20862 13634 20914
rect 13634 20862 13636 20914
rect 13580 20860 13636 20862
rect 9996 20636 10052 20692
rect 13468 20188 13524 20244
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 4284 19234 4340 19236
rect 4284 19182 4286 19234
rect 4286 19182 4338 19234
rect 4338 19182 4340 19234
rect 4284 19180 4340 19182
rect 14252 20748 14308 20804
rect 15148 22764 15204 22820
rect 15148 22092 15204 22148
rect 14924 20860 14980 20916
rect 14140 20188 14196 20244
rect 14588 20578 14644 20580
rect 14588 20526 14590 20578
rect 14590 20526 14642 20578
rect 14642 20526 14644 20578
rect 14588 20524 14644 20526
rect 15372 20690 15428 20692
rect 15372 20638 15374 20690
rect 15374 20638 15426 20690
rect 15426 20638 15428 20690
rect 15372 20636 15428 20638
rect 13804 19234 13860 19236
rect 13804 19182 13806 19234
rect 13806 19182 13858 19234
rect 13858 19182 13860 19234
rect 13804 19180 13860 19182
rect 14028 19122 14084 19124
rect 14028 19070 14030 19122
rect 14030 19070 14082 19122
rect 14082 19070 14084 19122
rect 14028 19068 14084 19070
rect 1932 18844 1988 18900
rect 11004 18844 11060 18900
rect 4284 18284 4340 18340
rect 14812 19234 14868 19236
rect 14812 19182 14814 19234
rect 14814 19182 14866 19234
rect 14866 19182 14868 19234
rect 14812 19180 14868 19182
rect 15036 19292 15092 19348
rect 14700 19122 14756 19124
rect 14700 19070 14702 19122
rect 14702 19070 14754 19122
rect 14754 19070 14756 19122
rect 14700 19068 14756 19070
rect 14364 18844 14420 18900
rect 15036 18508 15092 18564
rect 13468 18284 13524 18340
rect 1932 18226 1988 18228
rect 1932 18174 1934 18226
rect 1934 18174 1986 18226
rect 1986 18174 1988 18226
rect 1932 18172 1988 18174
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 14588 18450 14644 18452
rect 14588 18398 14590 18450
rect 14590 18398 14642 18450
rect 14642 18398 14644 18450
rect 14588 18396 14644 18398
rect 14812 18450 14868 18452
rect 14812 18398 14814 18450
rect 14814 18398 14866 18450
rect 14866 18398 14868 18450
rect 14812 18396 14868 18398
rect 14140 18284 14196 18340
rect 15260 20578 15316 20580
rect 15260 20526 15262 20578
rect 15262 20526 15314 20578
rect 15314 20526 15316 20578
rect 15260 20524 15316 20526
rect 16268 23436 16324 23492
rect 15596 22370 15652 22372
rect 15596 22318 15598 22370
rect 15598 22318 15650 22370
rect 15650 22318 15652 22370
rect 15596 22316 15652 22318
rect 16156 22316 16212 22372
rect 17388 24780 17444 24836
rect 20636 27858 20692 27860
rect 20636 27806 20638 27858
rect 20638 27806 20690 27858
rect 20690 27806 20692 27858
rect 20636 27804 20692 27806
rect 19404 26908 19460 26964
rect 19068 25676 19124 25732
rect 18284 24834 18340 24836
rect 18284 24782 18286 24834
rect 18286 24782 18338 24834
rect 18338 24782 18340 24834
rect 18284 24780 18340 24782
rect 17612 24722 17668 24724
rect 17612 24670 17614 24722
rect 17614 24670 17666 24722
rect 17666 24670 17668 24722
rect 17612 24668 17668 24670
rect 18620 24780 18676 24836
rect 17500 23996 17556 24052
rect 17388 23212 17444 23268
rect 16380 21868 16436 21924
rect 16492 21980 16548 22036
rect 15708 21362 15764 21364
rect 15708 21310 15710 21362
rect 15710 21310 15762 21362
rect 15762 21310 15764 21362
rect 15708 21308 15764 21310
rect 15820 20860 15876 20916
rect 15484 19740 15540 19796
rect 15484 19180 15540 19236
rect 16716 20972 16772 21028
rect 16828 21868 16884 21924
rect 16604 19180 16660 19236
rect 15260 18450 15316 18452
rect 15260 18398 15262 18450
rect 15262 18398 15314 18450
rect 15314 18398 15316 18450
rect 15260 18396 15316 18398
rect 15148 17836 15204 17892
rect 14700 17388 14756 17444
rect 18060 23660 18116 23716
rect 17612 22764 17668 22820
rect 17612 22428 17668 22484
rect 17724 22146 17780 22148
rect 17724 22094 17726 22146
rect 17726 22094 17778 22146
rect 17778 22094 17780 22146
rect 17724 22092 17780 22094
rect 17612 21868 17668 21924
rect 17724 21810 17780 21812
rect 17724 21758 17726 21810
rect 17726 21758 17778 21810
rect 17778 21758 17780 21810
rect 17724 21756 17780 21758
rect 18956 25282 19012 25284
rect 18956 25230 18958 25282
rect 18958 25230 19010 25282
rect 19010 25230 19012 25282
rect 18956 25228 19012 25230
rect 19180 25282 19236 25284
rect 19180 25230 19182 25282
rect 19182 25230 19234 25282
rect 19234 25230 19236 25282
rect 19180 25228 19236 25230
rect 18284 22258 18340 22260
rect 18284 22206 18286 22258
rect 18286 22206 18338 22258
rect 18338 22206 18340 22258
rect 18284 22204 18340 22206
rect 18956 24780 19012 24836
rect 18508 24108 18564 24164
rect 18620 23938 18676 23940
rect 18620 23886 18622 23938
rect 18622 23886 18674 23938
rect 18674 23886 18676 23938
rect 18620 23884 18676 23886
rect 18620 23436 18676 23492
rect 18844 23660 18900 23716
rect 18732 23378 18788 23380
rect 18732 23326 18734 23378
rect 18734 23326 18786 23378
rect 18786 23326 18788 23378
rect 18732 23324 18788 23326
rect 18508 23266 18564 23268
rect 18508 23214 18510 23266
rect 18510 23214 18562 23266
rect 18562 23214 18564 23266
rect 18508 23212 18564 23214
rect 18396 23154 18452 23156
rect 18396 23102 18398 23154
rect 18398 23102 18450 23154
rect 18450 23102 18452 23154
rect 18396 23100 18452 23102
rect 18060 21756 18116 21812
rect 18508 22764 18564 22820
rect 19068 23660 19124 23716
rect 18956 22930 19012 22932
rect 18956 22878 18958 22930
rect 18958 22878 19010 22930
rect 19010 22878 19012 22930
rect 18956 22876 19012 22878
rect 18844 22540 18900 22596
rect 18620 22316 18676 22372
rect 18732 21756 18788 21812
rect 18844 22204 18900 22260
rect 18732 21474 18788 21476
rect 18732 21422 18734 21474
rect 18734 21422 18786 21474
rect 18786 21422 18788 21474
rect 18732 21420 18788 21422
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 20300 27132 20356 27188
rect 20748 27074 20804 27076
rect 20748 27022 20750 27074
rect 20750 27022 20802 27074
rect 20802 27022 20804 27074
rect 20748 27020 20804 27022
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 22204 27074 22260 27076
rect 22204 27022 22206 27074
rect 22206 27022 22258 27074
rect 22258 27022 22260 27074
rect 22204 27020 22260 27022
rect 21308 26962 21364 26964
rect 21308 26910 21310 26962
rect 21310 26910 21362 26962
rect 21362 26910 21364 26962
rect 21308 26908 21364 26910
rect 22316 26962 22372 26964
rect 22316 26910 22318 26962
rect 22318 26910 22370 26962
rect 22370 26910 22372 26962
rect 22316 26908 22372 26910
rect 23436 26908 23492 26964
rect 24668 27858 24724 27860
rect 24668 27806 24670 27858
rect 24670 27806 24722 27858
rect 24722 27806 24724 27858
rect 24668 27804 24724 27806
rect 20300 25788 20356 25844
rect 20636 26290 20692 26292
rect 20636 26238 20638 26290
rect 20638 26238 20690 26290
rect 20690 26238 20692 26290
rect 20636 26236 20692 26238
rect 19740 25618 19796 25620
rect 19740 25566 19742 25618
rect 19742 25566 19794 25618
rect 19794 25566 19796 25618
rect 19740 25564 19796 25566
rect 19292 23324 19348 23380
rect 19516 23772 19572 23828
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 19740 23714 19796 23716
rect 19740 23662 19742 23714
rect 19742 23662 19794 23714
rect 19794 23662 19796 23714
rect 19740 23660 19796 23662
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 19852 23154 19908 23156
rect 19852 23102 19854 23154
rect 19854 23102 19906 23154
rect 19906 23102 19908 23154
rect 19852 23100 19908 23102
rect 19180 22370 19236 22372
rect 19180 22318 19182 22370
rect 19182 22318 19234 22370
rect 19234 22318 19236 22370
rect 19180 22316 19236 22318
rect 19292 21980 19348 22036
rect 19404 21644 19460 21700
rect 20412 22988 20468 23044
rect 20076 22428 20132 22484
rect 21532 26236 21588 26292
rect 21084 25564 21140 25620
rect 21644 25788 21700 25844
rect 21420 25228 21476 25284
rect 23548 24668 23604 24724
rect 21420 24050 21476 24052
rect 21420 23998 21422 24050
rect 21422 23998 21474 24050
rect 21474 23998 21476 24050
rect 21420 23996 21476 23998
rect 21308 23660 21364 23716
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 19628 21756 19684 21812
rect 17164 20188 17220 20244
rect 16044 18508 16100 18564
rect 16940 18508 16996 18564
rect 16604 18450 16660 18452
rect 16604 18398 16606 18450
rect 16606 18398 16658 18450
rect 16658 18398 16660 18450
rect 16604 18396 16660 18398
rect 15932 17836 15988 17892
rect 16268 18284 16324 18340
rect 15820 17276 15876 17332
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 16604 15372 16660 15428
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 16044 14252 16100 14308
rect 17500 18844 17556 18900
rect 17052 18284 17108 18340
rect 17500 18396 17556 18452
rect 16828 17500 16884 17556
rect 17052 17442 17108 17444
rect 17052 17390 17054 17442
rect 17054 17390 17106 17442
rect 17106 17390 17108 17442
rect 17052 17388 17108 17390
rect 17276 17442 17332 17444
rect 17276 17390 17278 17442
rect 17278 17390 17330 17442
rect 17330 17390 17332 17442
rect 17276 17388 17332 17390
rect 17724 18172 17780 18228
rect 18060 20188 18116 20244
rect 18284 19964 18340 20020
rect 18508 20578 18564 20580
rect 18508 20526 18510 20578
rect 18510 20526 18562 20578
rect 18562 20526 18564 20578
rect 18508 20524 18564 20526
rect 18396 19180 18452 19236
rect 18508 20300 18564 20356
rect 19292 20972 19348 21028
rect 19292 20412 19348 20468
rect 19068 20188 19124 20244
rect 20524 21644 20580 21700
rect 20412 21420 20468 21476
rect 19852 20802 19908 20804
rect 19852 20750 19854 20802
rect 19854 20750 19906 20802
rect 19906 20750 19908 20802
rect 19852 20748 19908 20750
rect 18956 19964 19012 20020
rect 18732 19292 18788 19348
rect 18284 18956 18340 19012
rect 18844 19234 18900 19236
rect 18844 19182 18846 19234
rect 18846 19182 18898 19234
rect 18898 19182 18900 19234
rect 18844 19180 18900 19182
rect 19180 18844 19236 18900
rect 19628 20636 19684 20692
rect 19516 20300 19572 20356
rect 19404 19740 19460 19796
rect 19404 18732 19460 18788
rect 19292 18620 19348 18676
rect 18620 18562 18676 18564
rect 18620 18510 18622 18562
rect 18622 18510 18674 18562
rect 18674 18510 18676 18562
rect 18620 18508 18676 18510
rect 19068 18508 19124 18564
rect 17612 17554 17668 17556
rect 17612 17502 17614 17554
rect 17614 17502 17666 17554
rect 17666 17502 17668 17554
rect 17612 17500 17668 17502
rect 17724 16492 17780 16548
rect 17388 15426 17444 15428
rect 17388 15374 17390 15426
rect 17390 15374 17442 15426
rect 17442 15374 17444 15426
rect 17388 15372 17444 15374
rect 16716 14252 16772 14308
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 18284 18284 18340 18340
rect 19180 18284 19236 18340
rect 18172 17388 18228 17444
rect 18844 18172 18900 18228
rect 19292 17948 19348 18004
rect 19404 18172 19460 18228
rect 18844 17612 18900 17668
rect 18732 16828 18788 16884
rect 19180 17388 19236 17444
rect 19068 17276 19124 17332
rect 19068 17052 19124 17108
rect 19292 16658 19348 16660
rect 19292 16606 19294 16658
rect 19294 16606 19346 16658
rect 19346 16606 19348 16658
rect 19292 16604 19348 16606
rect 19628 20412 19684 20468
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 20300 20188 20356 20244
rect 19628 19068 19684 19124
rect 19964 19292 20020 19348
rect 20300 19234 20356 19236
rect 20300 19182 20302 19234
rect 20302 19182 20354 19234
rect 20354 19182 20356 19234
rect 20300 19180 20356 19182
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 19740 18508 19796 18564
rect 19852 18450 19908 18452
rect 19852 18398 19854 18450
rect 19854 18398 19906 18450
rect 19906 18398 19908 18450
rect 19852 18396 19908 18398
rect 21308 22370 21364 22372
rect 21308 22318 21310 22370
rect 21310 22318 21362 22370
rect 21362 22318 21364 22370
rect 21308 22316 21364 22318
rect 22652 24556 22708 24612
rect 22540 24108 22596 24164
rect 23436 24108 23492 24164
rect 23212 23772 23268 23828
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 40236 26236 40292 26292
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 24668 24722 24724 24724
rect 24668 24670 24670 24722
rect 24670 24670 24722 24722
rect 24722 24670 24724 24722
rect 24668 24668 24724 24670
rect 25340 24722 25396 24724
rect 25340 24670 25342 24722
rect 25342 24670 25394 24722
rect 25394 24670 25396 24722
rect 25340 24668 25396 24670
rect 23884 24610 23940 24612
rect 23884 24558 23886 24610
rect 23886 24558 23938 24610
rect 23938 24558 23940 24610
rect 23884 24556 23940 24558
rect 22204 23154 22260 23156
rect 22204 23102 22206 23154
rect 22206 23102 22258 23154
rect 22258 23102 22260 23154
rect 22204 23100 22260 23102
rect 21644 22988 21700 23044
rect 21532 22092 21588 22148
rect 20636 20748 20692 20804
rect 21532 20802 21588 20804
rect 21532 20750 21534 20802
rect 21534 20750 21586 20802
rect 21586 20750 21588 20802
rect 21532 20748 21588 20750
rect 21308 20690 21364 20692
rect 21308 20638 21310 20690
rect 21310 20638 21362 20690
rect 21362 20638 21364 20690
rect 21308 20636 21364 20638
rect 21532 20300 21588 20356
rect 21196 19068 21252 19124
rect 21868 20802 21924 20804
rect 21868 20750 21870 20802
rect 21870 20750 21922 20802
rect 21922 20750 21924 20802
rect 21868 20748 21924 20750
rect 21756 20578 21812 20580
rect 21756 20526 21758 20578
rect 21758 20526 21810 20578
rect 21810 20526 21812 20578
rect 21756 20524 21812 20526
rect 21868 19964 21924 20020
rect 21756 19404 21812 19460
rect 20748 18620 20804 18676
rect 20188 17666 20244 17668
rect 20188 17614 20190 17666
rect 20190 17614 20242 17666
rect 20242 17614 20244 17666
rect 20188 17612 20244 17614
rect 19964 17554 20020 17556
rect 19964 17502 19966 17554
rect 19966 17502 20018 17554
rect 20018 17502 20020 17554
rect 19964 17500 20020 17502
rect 19740 17388 19796 17444
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 21644 18508 21700 18564
rect 22092 20076 22148 20132
rect 22092 19740 22148 19796
rect 22540 20748 22596 20804
rect 22540 19740 22596 19796
rect 22540 18956 22596 19012
rect 21980 18620 22036 18676
rect 22092 18508 22148 18564
rect 22428 18396 22484 18452
rect 21868 17666 21924 17668
rect 21868 17614 21870 17666
rect 21870 17614 21922 17666
rect 21922 17614 21924 17666
rect 21868 17612 21924 17614
rect 22092 17554 22148 17556
rect 22092 17502 22094 17554
rect 22094 17502 22146 17554
rect 22146 17502 22148 17554
rect 22092 17500 22148 17502
rect 21420 17052 21476 17108
rect 21756 17388 21812 17444
rect 19740 16658 19796 16660
rect 19740 16606 19742 16658
rect 19742 16606 19794 16658
rect 19794 16606 19796 16658
rect 19740 16604 19796 16606
rect 19852 16492 19908 16548
rect 19404 16380 19460 16436
rect 20300 16604 20356 16660
rect 20188 16492 20244 16548
rect 21420 16882 21476 16884
rect 21420 16830 21422 16882
rect 21422 16830 21474 16882
rect 21474 16830 21476 16882
rect 21420 16828 21476 16830
rect 20412 16380 20468 16436
rect 22876 23154 22932 23156
rect 22876 23102 22878 23154
rect 22878 23102 22930 23154
rect 22930 23102 22932 23154
rect 22876 23100 22932 23102
rect 22988 22988 23044 23044
rect 22764 20860 22820 20916
rect 23324 20802 23380 20804
rect 23324 20750 23326 20802
rect 23326 20750 23378 20802
rect 23378 20750 23380 20802
rect 23324 20748 23380 20750
rect 23660 20300 23716 20356
rect 23100 20130 23156 20132
rect 23100 20078 23102 20130
rect 23102 20078 23154 20130
rect 23154 20078 23156 20130
rect 23100 20076 23156 20078
rect 24220 22258 24276 22260
rect 24220 22206 24222 22258
rect 24222 22206 24274 22258
rect 24274 22206 24276 22258
rect 24220 22204 24276 22206
rect 26572 24668 26628 24724
rect 26348 23548 26404 23604
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 27356 23996 27412 24052
rect 27020 23714 27076 23716
rect 27020 23662 27022 23714
rect 27022 23662 27074 23714
rect 27074 23662 27076 23714
rect 27020 23660 27076 23662
rect 26684 23548 26740 23604
rect 27692 23436 27748 23492
rect 37660 23938 37716 23940
rect 37660 23886 37662 23938
rect 37662 23886 37714 23938
rect 37714 23886 37716 23938
rect 37660 23884 37716 23886
rect 28028 23826 28084 23828
rect 28028 23774 28030 23826
rect 28030 23774 28082 23826
rect 28082 23774 28084 23826
rect 28028 23772 28084 23774
rect 40012 24220 40068 24276
rect 37884 23548 37940 23604
rect 40012 23548 40068 23604
rect 29372 23436 29428 23492
rect 28140 23324 28196 23380
rect 29036 23324 29092 23380
rect 26908 23154 26964 23156
rect 26908 23102 26910 23154
rect 26910 23102 26962 23154
rect 26962 23102 26964 23154
rect 26908 23100 26964 23102
rect 28140 23100 28196 23156
rect 26348 22204 26404 22260
rect 23996 20860 24052 20916
rect 25116 20860 25172 20916
rect 22988 20018 23044 20020
rect 22988 19966 22990 20018
rect 22990 19966 23042 20018
rect 23042 19966 23044 20018
rect 22988 19964 23044 19966
rect 23996 20412 24052 20468
rect 22764 19740 22820 19796
rect 24668 20412 24724 20468
rect 24556 20242 24612 20244
rect 24556 20190 24558 20242
rect 24558 20190 24610 20242
rect 24610 20190 24612 20242
rect 24556 20188 24612 20190
rect 24444 20130 24500 20132
rect 24444 20078 24446 20130
rect 24446 20078 24498 20130
rect 24498 20078 24500 20130
rect 24444 20076 24500 20078
rect 26012 20188 26068 20244
rect 26908 21420 26964 21476
rect 24332 19964 24388 20020
rect 22764 19180 22820 19236
rect 23436 18674 23492 18676
rect 23436 18622 23438 18674
rect 23438 18622 23490 18674
rect 23490 18622 23492 18674
rect 23436 18620 23492 18622
rect 22764 18508 22820 18564
rect 22988 17890 23044 17892
rect 22988 17838 22990 17890
rect 22990 17838 23042 17890
rect 23042 17838 23044 17890
rect 22988 17836 23044 17838
rect 23772 17666 23828 17668
rect 23772 17614 23774 17666
rect 23774 17614 23826 17666
rect 23826 17614 23828 17666
rect 23772 17612 23828 17614
rect 22428 17388 22484 17444
rect 23324 17442 23380 17444
rect 23324 17390 23326 17442
rect 23326 17390 23378 17442
rect 23378 17390 23380 17442
rect 23324 17388 23380 17390
rect 22316 16940 22372 16996
rect 23548 16828 23604 16884
rect 19628 16098 19684 16100
rect 19628 16046 19630 16098
rect 19630 16046 19682 16098
rect 19682 16046 19684 16098
rect 19628 16044 19684 16046
rect 20524 16098 20580 16100
rect 20524 16046 20526 16098
rect 20526 16046 20578 16098
rect 20578 16046 20580 16098
rect 20524 16044 20580 16046
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 17500 5180 17556 5236
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 18732 5234 18788 5236
rect 18732 5182 18734 5234
rect 18734 5182 18786 5234
rect 18786 5182 18788 5234
rect 18732 5180 18788 5182
rect 19180 14306 19236 14308
rect 19180 14254 19182 14306
rect 19182 14254 19234 14306
rect 19234 14254 19236 14306
rect 19180 14252 19236 14254
rect 19404 13746 19460 13748
rect 19404 13694 19406 13746
rect 19406 13694 19458 13746
rect 19458 13694 19460 13746
rect 19404 13692 19460 13694
rect 18844 4060 18900 4116
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 25564 19292 25620 19348
rect 25676 18620 25732 18676
rect 25340 18396 25396 18452
rect 24332 16828 24388 16884
rect 24444 18060 24500 18116
rect 22652 13746 22708 13748
rect 22652 13694 22654 13746
rect 22654 13694 22706 13746
rect 22706 13694 22708 13746
rect 22652 13692 22708 13694
rect 21420 13468 21476 13524
rect 22204 13468 22260 13524
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 20076 4114 20132 4116
rect 20076 4062 20078 4114
rect 20078 4062 20130 4114
rect 20130 4062 20132 4114
rect 20076 4060 20132 4062
rect 24668 16882 24724 16884
rect 24668 16830 24670 16882
rect 24670 16830 24722 16882
rect 24722 16830 24724 16882
rect 24668 16828 24724 16830
rect 25004 15986 25060 15988
rect 25004 15934 25006 15986
rect 25006 15934 25058 15986
rect 25058 15934 25060 15986
rect 25004 15932 25060 15934
rect 26684 20130 26740 20132
rect 26684 20078 26686 20130
rect 26686 20078 26738 20130
rect 26738 20078 26740 20130
rect 26684 20076 26740 20078
rect 26460 20018 26516 20020
rect 26460 19966 26462 20018
rect 26462 19966 26514 20018
rect 26514 19966 26516 20018
rect 26460 19964 26516 19966
rect 29260 22988 29316 23044
rect 30268 23154 30324 23156
rect 30268 23102 30270 23154
rect 30270 23102 30322 23154
rect 30322 23102 30324 23154
rect 30268 23100 30324 23102
rect 37660 23154 37716 23156
rect 37660 23102 37662 23154
rect 37662 23102 37714 23154
rect 37714 23102 37716 23154
rect 37660 23100 37716 23102
rect 29820 23042 29876 23044
rect 29820 22990 29822 23042
rect 29822 22990 29874 23042
rect 29874 22990 29876 23042
rect 29820 22988 29876 22990
rect 40012 22930 40068 22932
rect 40012 22878 40014 22930
rect 40014 22878 40066 22930
rect 40066 22878 40068 22930
rect 40012 22876 40068 22878
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 28140 21474 28196 21476
rect 28140 21422 28142 21474
rect 28142 21422 28194 21474
rect 28194 21422 28196 21474
rect 28140 21420 28196 21422
rect 29484 20802 29540 20804
rect 29484 20750 29486 20802
rect 29486 20750 29538 20802
rect 29538 20750 29540 20802
rect 29484 20748 29540 20750
rect 30156 20860 30212 20916
rect 29148 20690 29204 20692
rect 29148 20638 29150 20690
rect 29150 20638 29202 20690
rect 29202 20638 29204 20690
rect 29148 20636 29204 20638
rect 26236 19404 26292 19460
rect 27244 19346 27300 19348
rect 27244 19294 27246 19346
rect 27246 19294 27298 19346
rect 27298 19294 27300 19346
rect 27244 19292 27300 19294
rect 26236 18956 26292 19012
rect 28252 20524 28308 20580
rect 26124 18060 26180 18116
rect 27580 17554 27636 17556
rect 27580 17502 27582 17554
rect 27582 17502 27634 17554
rect 27634 17502 27636 17554
rect 27580 17500 27636 17502
rect 26572 17388 26628 17444
rect 25676 16828 25732 16884
rect 25340 15932 25396 15988
rect 25004 15148 25060 15204
rect 27356 17388 27412 17444
rect 28364 19010 28420 19012
rect 28364 18958 28366 19010
rect 28366 18958 28418 19010
rect 28418 18958 28420 19010
rect 28364 18956 28420 18958
rect 28252 18732 28308 18788
rect 27804 17666 27860 17668
rect 27804 17614 27806 17666
rect 27806 17614 27858 17666
rect 27858 17614 27860 17666
rect 27804 17612 27860 17614
rect 27916 17554 27972 17556
rect 27916 17502 27918 17554
rect 27918 17502 27970 17554
rect 27970 17502 27972 17554
rect 27916 17500 27972 17502
rect 30828 20860 30884 20916
rect 30604 20802 30660 20804
rect 30604 20750 30606 20802
rect 30606 20750 30658 20802
rect 30658 20750 30660 20802
rect 30604 20748 30660 20750
rect 30716 20690 30772 20692
rect 30716 20638 30718 20690
rect 30718 20638 30770 20690
rect 30770 20638 30772 20690
rect 30716 20636 30772 20638
rect 30380 20578 30436 20580
rect 30380 20526 30382 20578
rect 30382 20526 30434 20578
rect 30434 20526 30436 20578
rect 30380 20524 30436 20526
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 31388 20636 31444 20692
rect 40012 21532 40068 21588
rect 37884 21420 37940 21476
rect 39900 20860 39956 20916
rect 37660 20802 37716 20804
rect 37660 20750 37662 20802
rect 37662 20750 37714 20802
rect 37714 20750 37716 20802
rect 37660 20748 37716 20750
rect 37548 20636 37604 20692
rect 40012 20188 40068 20244
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 40012 19516 40068 19572
rect 37660 19292 37716 19348
rect 29708 18732 29764 18788
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 29148 17666 29204 17668
rect 29148 17614 29150 17666
rect 29150 17614 29202 17666
rect 29202 17614 29204 17666
rect 29148 17612 29204 17614
rect 37660 17666 37716 17668
rect 37660 17614 37662 17666
rect 37662 17614 37714 17666
rect 37714 17614 37716 17666
rect 37660 17612 37716 17614
rect 28252 17500 28308 17556
rect 29260 17554 29316 17556
rect 29260 17502 29262 17554
rect 29262 17502 29314 17554
rect 29314 17502 29316 17554
rect 29260 17500 29316 17502
rect 30156 17500 30212 17556
rect 26908 16716 26964 16772
rect 28588 16716 28644 16772
rect 26796 16156 26852 16212
rect 40012 17500 40068 17556
rect 37660 16716 37716 16772
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 27580 15484 27636 15540
rect 29260 16210 29316 16212
rect 29260 16158 29262 16210
rect 29262 16158 29314 16210
rect 29314 16158 29316 16210
rect 29260 16156 29316 16158
rect 40012 16156 40068 16212
rect 28588 15484 28644 15540
rect 27244 15090 27300 15092
rect 27244 15038 27246 15090
rect 27246 15038 27298 15090
rect 27298 15038 27300 15090
rect 27244 15036 27300 15038
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 23548 3612 23604 3668
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 25564 3666 25620 3668
rect 25564 3614 25566 3666
rect 25566 3614 25618 3666
rect 25618 3614 25620 3666
rect 25564 3612 25620 3614
rect 25564 3388 25620 3444
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 26796 3388 26852 3444
<< metal3 >>
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 22866 38220 22876 38276
rect 22932 38220 25564 38276
rect 25620 38220 25630 38276
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 20850 37436 20860 37492
rect 20916 37436 22092 37492
rect 22148 37436 22158 37492
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 18722 27804 18732 27860
rect 18788 27804 19292 27860
rect 19348 27804 19358 27860
rect 20626 27804 20636 27860
rect 20692 27804 24668 27860
rect 24724 27804 24734 27860
rect 0 27636 800 27664
rect 0 27580 4172 27636
rect 4228 27580 4238 27636
rect 0 27552 800 27580
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 20290 27132 20300 27188
rect 20356 27132 22260 27188
rect 22204 27076 22260 27132
rect 4274 27020 4284 27076
rect 4340 27020 8428 27076
rect 18610 27020 18620 27076
rect 18676 27020 20748 27076
rect 20804 27020 20814 27076
rect 22194 27020 22204 27076
rect 22260 27020 22270 27076
rect 0 26964 800 26992
rect 8372 26964 8428 27020
rect 0 26908 2044 26964
rect 2100 26908 2110 26964
rect 8372 26908 11452 26964
rect 11508 26908 14364 26964
rect 14420 26908 14430 26964
rect 17714 26908 17724 26964
rect 17780 26908 18620 26964
rect 18676 26908 18732 26964
rect 18788 26908 18798 26964
rect 18946 26908 18956 26964
rect 19012 26908 19404 26964
rect 19460 26908 21308 26964
rect 21364 26908 21374 26964
rect 22306 26908 22316 26964
rect 22372 26908 23436 26964
rect 23492 26908 23502 26964
rect 0 26880 800 26908
rect 17042 26796 17052 26852
rect 17108 26796 17836 26852
rect 17892 26796 17902 26852
rect 13458 26684 13468 26740
rect 13524 26684 15372 26740
rect 15428 26684 15438 26740
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 14914 26460 14924 26516
rect 14980 26460 15596 26516
rect 15652 26460 15662 26516
rect 0 26292 800 26320
rect 41200 26292 42000 26320
rect 0 26236 1932 26292
rect 1988 26236 1998 26292
rect 4274 26236 4284 26292
rect 4340 26236 11788 26292
rect 11844 26236 15260 26292
rect 15316 26236 15326 26292
rect 20626 26236 20636 26292
rect 20692 26236 21532 26292
rect 21588 26236 21598 26292
rect 40226 26236 40236 26292
rect 40292 26236 42000 26292
rect 0 26208 800 26236
rect 41200 26208 42000 26236
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 15092 25788 20300 25844
rect 20356 25788 21644 25844
rect 21700 25788 21710 25844
rect 14578 25676 14588 25732
rect 14644 25676 15036 25732
rect 15092 25676 15148 25788
rect 18274 25676 18284 25732
rect 18340 25676 19068 25732
rect 19124 25676 19134 25732
rect 15474 25564 15484 25620
rect 15540 25564 17836 25620
rect 17892 25564 19740 25620
rect 19796 25564 21084 25620
rect 21140 25564 21150 25620
rect 14018 25340 14028 25396
rect 14084 25340 15372 25396
rect 15428 25340 16492 25396
rect 16548 25340 16558 25396
rect 17938 25228 17948 25284
rect 18004 25228 18956 25284
rect 19012 25228 19022 25284
rect 19170 25228 19180 25284
rect 19236 25228 21420 25284
rect 21476 25228 21486 25284
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 16146 24892 16156 24948
rect 16212 24892 17500 24948
rect 17556 24892 17566 24948
rect 17378 24780 17388 24836
rect 17444 24780 18284 24836
rect 18340 24780 18350 24836
rect 18610 24780 18620 24836
rect 18676 24780 18956 24836
rect 19012 24780 19022 24836
rect 16482 24668 16492 24724
rect 16548 24668 17612 24724
rect 17668 24668 17678 24724
rect 23538 24668 23548 24724
rect 23604 24668 24668 24724
rect 24724 24668 25340 24724
rect 25396 24668 26572 24724
rect 26628 24668 26638 24724
rect 22642 24556 22652 24612
rect 22708 24556 23884 24612
rect 23940 24556 23950 24612
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 41200 24276 42000 24304
rect 40002 24220 40012 24276
rect 40068 24220 42000 24276
rect 41200 24192 42000 24220
rect 13458 24108 13468 24164
rect 13524 24108 18508 24164
rect 18564 24108 22540 24164
rect 22596 24108 23436 24164
rect 23492 24108 23502 24164
rect 14242 23996 14252 24052
rect 14308 23996 15708 24052
rect 15764 23996 17500 24052
rect 17556 23996 17566 24052
rect 21410 23996 21420 24052
rect 21476 23996 27356 24052
rect 27412 23996 27422 24052
rect 14130 23884 14140 23940
rect 14196 23884 15596 23940
rect 15652 23884 15662 23940
rect 18582 23884 18620 23940
rect 18676 23884 18686 23940
rect 31892 23884 37660 23940
rect 37716 23884 37726 23940
rect 19506 23772 19516 23828
rect 19572 23772 23212 23828
rect 23268 23772 28028 23828
rect 28084 23772 28094 23828
rect 31892 23716 31948 23884
rect 18050 23660 18060 23716
rect 18116 23660 18844 23716
rect 18900 23660 18910 23716
rect 19058 23660 19068 23716
rect 19124 23660 19740 23716
rect 19796 23660 21308 23716
rect 21364 23660 21374 23716
rect 27010 23660 27020 23716
rect 27076 23660 31948 23716
rect 41200 23604 42000 23632
rect 26338 23548 26348 23604
rect 26404 23548 26684 23604
rect 26740 23548 37884 23604
rect 37940 23548 37950 23604
rect 40002 23548 40012 23604
rect 40068 23548 42000 23604
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 41200 23520 42000 23548
rect 16258 23436 16268 23492
rect 16324 23436 18620 23492
rect 18676 23436 18686 23492
rect 27682 23436 27692 23492
rect 27748 23436 29372 23492
rect 29428 23436 29438 23492
rect 18722 23324 18732 23380
rect 18788 23324 19292 23380
rect 19348 23324 19358 23380
rect 28130 23324 28140 23380
rect 28196 23324 29036 23380
rect 29092 23324 29102 23380
rect 17378 23212 17388 23268
rect 17444 23212 18508 23268
rect 18564 23212 18574 23268
rect 18386 23100 18396 23156
rect 18452 23100 19852 23156
rect 19908 23100 19918 23156
rect 22194 23100 22204 23156
rect 22260 23100 22876 23156
rect 22932 23100 22942 23156
rect 26898 23100 26908 23156
rect 26964 23100 28140 23156
rect 28196 23100 30268 23156
rect 30324 23100 30334 23156
rect 31892 23100 37660 23156
rect 37716 23100 37726 23156
rect 31892 23044 31948 23100
rect 20402 22988 20412 23044
rect 20468 22988 21644 23044
rect 21700 22988 22988 23044
rect 23044 22988 23054 23044
rect 29250 22988 29260 23044
rect 29316 22988 29820 23044
rect 29876 22988 31948 23044
rect 41200 22932 42000 22960
rect 14802 22876 14812 22932
rect 14868 22876 18956 22932
rect 19012 22876 19022 22932
rect 40002 22876 40012 22932
rect 40068 22876 42000 22932
rect 41200 22848 42000 22876
rect 15138 22764 15148 22820
rect 15204 22764 17612 22820
rect 17668 22764 18508 22820
rect 18564 22764 18574 22820
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 18834 22540 18844 22596
rect 18900 22540 19628 22596
rect 19684 22540 19694 22596
rect 17602 22428 17612 22484
rect 17668 22428 20076 22484
rect 20132 22428 20142 22484
rect 14466 22316 14476 22372
rect 14532 22316 15596 22372
rect 15652 22316 15662 22372
rect 16146 22316 16156 22372
rect 16212 22316 18620 22372
rect 18676 22316 19180 22372
rect 19236 22316 21308 22372
rect 21364 22316 21374 22372
rect 18274 22204 18284 22260
rect 18340 22204 18844 22260
rect 18900 22204 18910 22260
rect 24210 22204 24220 22260
rect 24276 22204 26348 22260
rect 26404 22204 26414 22260
rect 12338 22092 12348 22148
rect 12404 22092 13580 22148
rect 13636 22092 13646 22148
rect 14018 22092 14028 22148
rect 14084 22092 15148 22148
rect 15204 22092 17724 22148
rect 17780 22092 17790 22148
rect 19292 22092 21532 22148
rect 21588 22092 21598 22148
rect 19292 22036 19348 22092
rect 16482 21980 16492 22036
rect 16548 21980 19292 22036
rect 19348 21980 19358 22036
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 16370 21868 16380 21924
rect 16436 21868 16828 21924
rect 16884 21868 17612 21924
rect 17668 21868 17678 21924
rect 17714 21756 17724 21812
rect 17780 21756 18060 21812
rect 18116 21756 18732 21812
rect 18788 21756 19628 21812
rect 19684 21756 19694 21812
rect 4162 21644 4172 21700
rect 4228 21644 19404 21700
rect 19460 21644 20524 21700
rect 20580 21644 20590 21700
rect 41200 21588 42000 21616
rect 4274 21532 4284 21588
rect 4340 21532 9996 21588
rect 10052 21532 10062 21588
rect 11554 21532 11564 21588
rect 11620 21532 12236 21588
rect 12292 21532 12796 21588
rect 12852 21532 12862 21588
rect 40002 21532 40012 21588
rect 40068 21532 42000 21588
rect 41200 21504 42000 21532
rect 18722 21420 18732 21476
rect 18788 21420 20412 21476
rect 20468 21420 20478 21476
rect 26898 21420 26908 21476
rect 26964 21420 28140 21476
rect 28196 21420 37884 21476
rect 37940 21420 37950 21476
rect 14242 21308 14252 21364
rect 14308 21308 15708 21364
rect 15764 21308 15774 21364
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 16706 20972 16716 21028
rect 16772 20972 19292 21028
rect 19348 20972 19358 21028
rect 0 20916 800 20944
rect 41200 20916 42000 20944
rect 0 20860 1932 20916
rect 1988 20860 1998 20916
rect 12786 20860 12796 20916
rect 12852 20860 13580 20916
rect 13636 20860 14924 20916
rect 14980 20860 14990 20916
rect 15810 20860 15820 20916
rect 15876 20860 22764 20916
rect 22820 20860 23996 20916
rect 24052 20860 25116 20916
rect 25172 20860 25182 20916
rect 30146 20860 30156 20916
rect 30212 20860 30828 20916
rect 30884 20860 31948 20916
rect 39890 20860 39900 20916
rect 39956 20860 42000 20916
rect 0 20832 800 20860
rect 21868 20804 21924 20860
rect 31892 20804 31948 20860
rect 41200 20832 42000 20860
rect 12114 20748 12124 20804
rect 12180 20748 14252 20804
rect 14308 20748 14318 20804
rect 19842 20748 19852 20804
rect 19908 20748 20636 20804
rect 20692 20748 21532 20804
rect 21588 20748 21598 20804
rect 21858 20748 21868 20804
rect 21924 20748 21934 20804
rect 22530 20748 22540 20804
rect 22596 20748 23324 20804
rect 23380 20748 23390 20804
rect 29474 20748 29484 20804
rect 29540 20748 30604 20804
rect 30660 20748 30670 20804
rect 31892 20748 37660 20804
rect 37716 20748 37726 20804
rect 9986 20636 9996 20692
rect 10052 20636 15372 20692
rect 15428 20636 15438 20692
rect 19618 20636 19628 20692
rect 19684 20636 21308 20692
rect 21364 20636 21374 20692
rect 26852 20636 29148 20692
rect 29204 20636 29214 20692
rect 30706 20636 30716 20692
rect 30772 20636 31388 20692
rect 31444 20636 37548 20692
rect 37604 20636 37614 20692
rect 26852 20580 26908 20636
rect 14578 20524 14588 20580
rect 14644 20524 15260 20580
rect 15316 20524 15326 20580
rect 18498 20524 18508 20580
rect 18564 20524 21588 20580
rect 21746 20524 21756 20580
rect 21812 20524 26908 20580
rect 28242 20524 28252 20580
rect 28308 20524 30380 20580
rect 30436 20524 30446 20580
rect 21532 20468 21588 20524
rect 19282 20412 19292 20468
rect 19348 20412 19628 20468
rect 19684 20412 19694 20468
rect 21532 20412 23996 20468
rect 24052 20412 24668 20468
rect 24724 20412 24734 20468
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 18498 20300 18508 20356
rect 18564 20300 19516 20356
rect 19572 20300 19582 20356
rect 20524 20300 21532 20356
rect 21588 20300 23660 20356
rect 23716 20300 23726 20356
rect 13458 20188 13468 20244
rect 13524 20188 14140 20244
rect 14196 20188 14206 20244
rect 17154 20188 17164 20244
rect 17220 20188 18060 20244
rect 18116 20188 18900 20244
rect 19058 20188 19068 20244
rect 19124 20188 20300 20244
rect 20356 20188 20366 20244
rect 18844 20132 18900 20188
rect 20524 20132 20580 20300
rect 41200 20244 42000 20272
rect 24546 20188 24556 20244
rect 24612 20188 26012 20244
rect 26068 20188 26078 20244
rect 40002 20188 40012 20244
rect 40068 20188 42000 20244
rect 41200 20160 42000 20188
rect 18844 20076 20580 20132
rect 22082 20076 22092 20132
rect 22148 20076 23100 20132
rect 23156 20076 23166 20132
rect 24434 20076 24444 20132
rect 24500 20076 26684 20132
rect 26740 20076 26750 20132
rect 18274 19964 18284 20020
rect 18340 19964 18956 20020
rect 19012 19964 19022 20020
rect 21858 19964 21868 20020
rect 21924 19964 22988 20020
rect 23044 19964 23054 20020
rect 24322 19964 24332 20020
rect 24388 19964 26460 20020
rect 26516 19964 26526 20020
rect 15092 19740 15484 19796
rect 15540 19740 19404 19796
rect 19460 19740 22092 19796
rect 22148 19740 22158 19796
rect 22530 19740 22540 19796
rect 22596 19740 22764 19796
rect 22820 19740 22830 19796
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 15026 19292 15036 19348
rect 15092 19292 15148 19740
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 41200 19572 42000 19600
rect 40002 19516 40012 19572
rect 40068 19516 42000 19572
rect 41200 19488 42000 19516
rect 21746 19404 21756 19460
rect 21812 19404 26236 19460
rect 26292 19404 26302 19460
rect 18722 19292 18732 19348
rect 18788 19292 19964 19348
rect 20020 19292 20030 19348
rect 25554 19292 25564 19348
rect 25620 19292 27244 19348
rect 27300 19292 37660 19348
rect 37716 19292 37726 19348
rect 4274 19180 4284 19236
rect 4340 19180 8428 19236
rect 13794 19180 13804 19236
rect 13860 19180 14812 19236
rect 14868 19180 15484 19236
rect 15540 19180 16604 19236
rect 16660 19180 16670 19236
rect 18386 19180 18396 19236
rect 18452 19180 18844 19236
rect 18900 19180 18910 19236
rect 20290 19180 20300 19236
rect 20356 19180 22764 19236
rect 22820 19180 22830 19236
rect 0 18900 800 18928
rect 8372 18900 8428 19180
rect 14018 19068 14028 19124
rect 14084 19068 14700 19124
rect 14756 19068 14766 19124
rect 19618 19068 19628 19124
rect 19684 19068 21196 19124
rect 21252 19068 21262 19124
rect 18274 18956 18284 19012
rect 18340 18956 22540 19012
rect 22596 18956 22606 19012
rect 26226 18956 26236 19012
rect 26292 18956 28364 19012
rect 28420 18956 28430 19012
rect 0 18844 1932 18900
rect 1988 18844 1998 18900
rect 8372 18844 11004 18900
rect 11060 18844 14364 18900
rect 14420 18844 14430 18900
rect 17490 18844 17500 18900
rect 17556 18844 19180 18900
rect 19236 18844 19684 18900
rect 0 18816 800 18844
rect 19394 18732 19404 18788
rect 19460 18732 19572 18788
rect 19282 18620 19292 18676
rect 19348 18620 19358 18676
rect 15026 18508 15036 18564
rect 15092 18508 16044 18564
rect 16100 18508 16940 18564
rect 16996 18508 17006 18564
rect 18610 18508 18620 18564
rect 18676 18508 19068 18564
rect 19124 18508 19134 18564
rect 19292 18452 19348 18620
rect 19516 18564 19572 18732
rect 13468 18396 14588 18452
rect 14644 18396 14654 18452
rect 14802 18396 14812 18452
rect 14868 18396 15260 18452
rect 15316 18396 15326 18452
rect 16594 18396 16604 18452
rect 16660 18396 17500 18452
rect 17556 18396 19348 18452
rect 19404 18508 19572 18564
rect 19628 18564 19684 18844
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 28242 18732 28252 18788
rect 28308 18732 29708 18788
rect 29764 18732 29774 18788
rect 20738 18620 20748 18676
rect 20804 18620 21980 18676
rect 22036 18620 23436 18676
rect 23492 18620 25676 18676
rect 25732 18620 25742 18676
rect 19628 18508 19740 18564
rect 19796 18508 21644 18564
rect 21700 18508 21710 18564
rect 22082 18508 22092 18564
rect 22148 18508 22764 18564
rect 22820 18508 22830 18564
rect 13468 18340 13524 18396
rect 16604 18340 16660 18396
rect 4274 18284 4284 18340
rect 4340 18284 13468 18340
rect 13524 18284 13534 18340
rect 14130 18284 14140 18340
rect 14196 18284 16268 18340
rect 16324 18284 16660 18340
rect 17042 18284 17052 18340
rect 17108 18284 18284 18340
rect 18340 18284 19180 18340
rect 19236 18284 19246 18340
rect 0 18228 800 18256
rect 19404 18228 19460 18508
rect 19618 18396 19628 18452
rect 19684 18396 19852 18452
rect 19908 18396 19918 18452
rect 22418 18396 22428 18452
rect 22484 18396 25340 18452
rect 25396 18396 25406 18452
rect 0 18172 1932 18228
rect 1988 18172 1998 18228
rect 17714 18172 17724 18228
rect 17780 18172 18844 18228
rect 18900 18172 18910 18228
rect 19394 18172 19404 18228
rect 19460 18172 19470 18228
rect 0 18144 800 18172
rect 24434 18060 24444 18116
rect 24500 18060 26124 18116
rect 26180 18060 26190 18116
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 24444 18004 24500 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 19282 17948 19292 18004
rect 19348 17948 24500 18004
rect 15138 17836 15148 17892
rect 15204 17836 15932 17892
rect 15988 17836 22988 17892
rect 23044 17836 23054 17892
rect 18834 17612 18844 17668
rect 18900 17612 20188 17668
rect 20244 17612 20254 17668
rect 21858 17612 21868 17668
rect 21924 17612 23772 17668
rect 23828 17612 23838 17668
rect 27794 17612 27804 17668
rect 27860 17612 29148 17668
rect 29204 17612 29214 17668
rect 31892 17612 37660 17668
rect 37716 17612 37726 17668
rect 31892 17556 31948 17612
rect 41200 17556 42000 17584
rect 16818 17500 16828 17556
rect 16884 17500 17612 17556
rect 17668 17500 17678 17556
rect 19954 17500 19964 17556
rect 20020 17500 22092 17556
rect 22148 17500 27580 17556
rect 27636 17500 27646 17556
rect 27906 17500 27916 17556
rect 27972 17500 28252 17556
rect 28308 17500 28318 17556
rect 29250 17500 29260 17556
rect 29316 17500 30156 17556
rect 30212 17500 31948 17556
rect 40002 17500 40012 17556
rect 40068 17500 42000 17556
rect 41200 17472 42000 17500
rect 14690 17388 14700 17444
rect 14756 17388 17052 17444
rect 17108 17388 17118 17444
rect 17266 17388 17276 17444
rect 17332 17388 18172 17444
rect 18228 17388 18238 17444
rect 19170 17388 19180 17444
rect 19236 17388 19740 17444
rect 19796 17388 19806 17444
rect 21746 17388 21756 17444
rect 21812 17388 22428 17444
rect 22484 17388 22494 17444
rect 23314 17388 23324 17444
rect 23380 17388 26572 17444
rect 26628 17388 27356 17444
rect 27412 17388 27422 17444
rect 15810 17276 15820 17332
rect 15876 17276 19068 17332
rect 19124 17276 19134 17332
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 19058 17052 19068 17108
rect 19124 17052 21420 17108
rect 21476 17052 21486 17108
rect 21084 16940 22316 16996
rect 22372 16940 22382 16996
rect 21084 16884 21140 16940
rect 17724 16828 18732 16884
rect 18788 16828 18798 16884
rect 20524 16828 21140 16884
rect 21410 16828 21420 16884
rect 21476 16828 23548 16884
rect 23604 16828 24332 16884
rect 24388 16828 24668 16884
rect 24724 16828 25676 16884
rect 25732 16828 26908 16884
rect 17724 16548 17780 16828
rect 19282 16604 19292 16660
rect 19348 16604 19740 16660
rect 19796 16604 20300 16660
rect 20356 16604 20366 16660
rect 20524 16548 20580 16828
rect 26852 16716 26908 16828
rect 26964 16716 26974 16772
rect 28578 16716 28588 16772
rect 28644 16716 37660 16772
rect 37716 16716 37726 16772
rect 17714 16492 17724 16548
rect 17780 16492 17790 16548
rect 19618 16492 19628 16548
rect 19684 16492 19852 16548
rect 19908 16492 19918 16548
rect 20178 16492 20188 16548
rect 20244 16492 20580 16548
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 19394 16380 19404 16436
rect 19460 16380 20412 16436
rect 20468 16380 20478 16436
rect 41200 16212 42000 16240
rect 26786 16156 26796 16212
rect 26852 16156 29260 16212
rect 29316 16156 29326 16212
rect 40002 16156 40012 16212
rect 40068 16156 42000 16212
rect 41200 16128 42000 16156
rect 19618 16044 19628 16100
rect 19684 16044 20524 16100
rect 20580 16044 20590 16100
rect 24994 15932 25004 15988
rect 25060 15932 25340 15988
rect 25396 15932 25406 15988
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 27570 15484 27580 15540
rect 27636 15484 28588 15540
rect 28644 15484 28654 15540
rect 16594 15372 16604 15428
rect 16660 15372 17388 15428
rect 17444 15372 17454 15428
rect 24994 15148 25004 15204
rect 25060 15148 27300 15204
rect 27244 15092 27300 15148
rect 27234 15036 27244 15092
rect 27300 15036 27310 15092
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 16034 14252 16044 14308
rect 16100 14252 16716 14308
rect 16772 14252 19180 14308
rect 19236 14252 19246 14308
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 19394 13692 19404 13748
rect 19460 13692 22652 13748
rect 22708 13692 22718 13748
rect 21410 13468 21420 13524
rect 21476 13468 22204 13524
rect 22260 13468 22270 13524
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 17490 5180 17500 5236
rect 17556 5180 18732 5236
rect 18788 5180 18798 5236
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 18834 4060 18844 4116
rect 18900 4060 20076 4116
rect 20132 4060 20142 4116
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 23538 3612 23548 3668
rect 23604 3612 25564 3668
rect 25620 3612 25630 3668
rect 25554 3388 25564 3444
rect 25620 3388 26796 3444
rect 26852 3388 26862 3444
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
<< via3 >>
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 18620 26908 18676 26964
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 18620 23884 18676 23940
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 19628 22540 19684 22596
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 19628 18396 19684 18452
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 19628 16492 19684 16548
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
<< metal4 >>
rect 4448 38444 4768 38476
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 19808 37660 20128 38476
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19808 34524 20128 36036
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 18620 26964 18676 26974
rect 18620 23940 18676 26908
rect 18620 23874 18676 23884
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 19808 23548 20128 25060
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 19628 22596 19684 22606
rect 19628 18452 19684 22540
rect 19628 16548 19684 18396
rect 19628 16482 19684 16492
rect 19808 21980 20128 23492
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 38444 35488 38476
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _099_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 23184 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _100_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 15680 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _101_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 20048 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _102_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21168 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _103_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 27216 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _104_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 29568 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _105_
timestamp 1698175906
transform 1 0 19936 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _106_
timestamp 1698175906
transform 1 0 17360 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _107_
timestamp 1698175906
transform -1 0 22064 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _108_
timestamp 1698175906
transform 1 0 15344 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _109_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 20720 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _110_
timestamp 1698175906
transform 1 0 27888 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _111_
timestamp 1698175906
transform -1 0 22624 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _112_
timestamp 1698175906
transform 1 0 17584 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _113_
timestamp 1698175906
transform -1 0 23184 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _114_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 20496 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _115_
timestamp 1698175906
transform 1 0 18032 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _116_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 20496 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _117_
timestamp 1698175906
transform 1 0 20048 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _118_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 18928 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _119_
timestamp 1698175906
transform 1 0 18704 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _120_
timestamp 1698175906
transform 1 0 18928 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _121_
timestamp 1698175906
transform 1 0 22064 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _122_
timestamp 1698175906
transform -1 0 21952 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _123_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 20944 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _124_
timestamp 1698175906
transform -1 0 20720 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _125_
timestamp 1698175906
transform 1 0 16688 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _126_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 20272 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _127_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21168 0 1 18816
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _128_
timestamp 1698175906
transform 1 0 29904 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _129_
timestamp 1698175906
transform -1 0 28672 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _130_
timestamp 1698175906
transform 1 0 21168 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _131_
timestamp 1698175906
transform 1 0 21168 0 1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _132_
timestamp 1698175906
transform 1 0 15232 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _133_
timestamp 1698175906
transform -1 0 17024 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _134_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 13776 0 1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _135_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 14224 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _136_
timestamp 1698175906
transform 1 0 18480 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _137_
timestamp 1698175906
transform 1 0 18256 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _138_
timestamp 1698175906
transform 1 0 13328 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _139_
timestamp 1698175906
transform -1 0 20832 0 -1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _140_
timestamp 1698175906
transform -1 0 18816 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _141_
timestamp 1698175906
transform -1 0 14448 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _142_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17472 0 1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _143_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 13328 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _144_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 22400 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _145_
timestamp 1698175906
transform -1 0 17920 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _146_
timestamp 1698175906
transform 1 0 18256 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _147_
timestamp 1698175906
transform -1 0 20384 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _148_
timestamp 1698175906
transform 1 0 18928 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _149_
timestamp 1698175906
transform 1 0 18480 0 1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _150_
timestamp 1698175906
transform 1 0 17248 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _151_
timestamp 1698175906
transform -1 0 15904 0 -1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _152_
timestamp 1698175906
transform 1 0 13328 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _153_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 23856 0 -1 18816
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _154_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 18256 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _155_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19040 0 1 17248
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _156_
timestamp 1698175906
transform 1 0 18256 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _157_
timestamp 1698175906
transform 1 0 23520 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _158_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 22512 0 1 17248
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _159_
timestamp 1698175906
transform -1 0 26992 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _160_
timestamp 1698175906
transform -1 0 19712 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _161_
timestamp 1698175906
transform 1 0 25984 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _162_
timestamp 1698175906
transform 1 0 22848 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _163_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 24864 0 -1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _164_
timestamp 1698175906
transform -1 0 30912 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _165_
timestamp 1698175906
transform 1 0 22288 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _166_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21168 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _167_
timestamp 1698175906
transform -1 0 29904 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _168_
timestamp 1698175906
transform 1 0 24864 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _169_
timestamp 1698175906
transform -1 0 24864 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _170_
timestamp 1698175906
transform 1 0 17920 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _171_
timestamp 1698175906
transform 1 0 18032 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _172_
timestamp 1698175906
transform 1 0 18480 0 -1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _173_
timestamp 1698175906
transform -1 0 17920 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _174_
timestamp 1698175906
transform 1 0 22064 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _175_
timestamp 1698175906
transform 1 0 21168 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _176_
timestamp 1698175906
transform 1 0 25088 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _177_
timestamp 1698175906
transform -1 0 25760 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _178_
timestamp 1698175906
transform -1 0 17136 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _179_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 15456 0 -1 21952
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _180_
timestamp 1698175906
transform 1 0 15792 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _181_
timestamp 1698175906
transform 1 0 14224 0 1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _182_
timestamp 1698175906
transform 1 0 13328 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _183_
timestamp 1698175906
transform 1 0 22624 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _184_
timestamp 1698175906
transform 1 0 27104 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _185_
timestamp 1698175906
transform -1 0 27104 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _186_
timestamp 1698175906
transform 1 0 23632 0 1 21952
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _187_
timestamp 1698175906
transform 1 0 23408 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _188_
timestamp 1698175906
transform -1 0 29456 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _189_
timestamp 1698175906
transform 1 0 27216 0 1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _190_
timestamp 1698175906
transform -1 0 17808 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _191_
timestamp 1698175906
transform -1 0 18144 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _192_
timestamp 1698175906
transform 1 0 16576 0 1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _193_
timestamp 1698175906
transform 1 0 15008 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _194_
timestamp 1698175906
transform -1 0 19712 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _195_
timestamp 1698175906
transform -1 0 15008 0 1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _196_
timestamp 1698175906
transform -1 0 15120 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _197_
timestamp 1698175906
transform -1 0 16016 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _198_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 26768 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _199_
timestamp 1698175906
transform 1 0 19152 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _200_
timestamp 1698175906
transform 1 0 27552 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _201_
timestamp 1698175906
transform -1 0 14560 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _202_
timestamp 1698175906
transform 1 0 16800 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _203_
timestamp 1698175906
transform 1 0 12096 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _204_
timestamp 1698175906
transform 1 0 11424 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _205_
timestamp 1698175906
transform -1 0 24864 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _206_
timestamp 1698175906
transform 1 0 17696 0 1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _207_
timestamp 1698175906
transform 1 0 15232 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _208_
timestamp 1698175906
transform -1 0 14896 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _209_
timestamp 1698175906
transform 1 0 21168 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _210_
timestamp 1698175906
transform 1 0 25088 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _211_
timestamp 1698175906
transform 1 0 28336 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _212_
timestamp 1698175906
transform 1 0 23296 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _213_
timestamp 1698175906
transform 1 0 15680 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _214_
timestamp 1698175906
transform 1 0 20384 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _215_
timestamp 1698175906
transform 1 0 24192 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _216_
timestamp 1698175906
transform -1 0 14112 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _217_
timestamp 1698175906
transform 1 0 25536 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _218_
timestamp 1698175906
transform 1 0 23296 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _219_
timestamp 1698175906
transform 1 0 27104 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _220_
timestamp 1698175906
transform 1 0 13776 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _221_
timestamp 1698175906
transform -1 0 13104 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _222_
timestamp 1698175906
transform -1 0 16576 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _225_
timestamp 1698175906
transform 1 0 26544 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _226_
timestamp 1698175906
transform 1 0 18256 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _227_
timestamp 1698175906
transform 1 0 23632 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__198__CLK dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 30240 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__199__CLK
timestamp 1698175906
transform 1 0 22624 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__200__CLK
timestamp 1698175906
transform 1 0 27328 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__201__CLK
timestamp 1698175906
transform 1 0 14784 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__202__CLK
timestamp 1698175906
transform 1 0 21056 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__203__CLK
timestamp 1698175906
transform 1 0 15344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__204__CLK
timestamp 1698175906
transform 1 0 14896 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__205__CLK
timestamp 1698175906
transform 1 0 25312 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__206__CLK
timestamp 1698175906
transform 1 0 21392 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__207__CLK
timestamp 1698175906
transform 1 0 19712 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__208__CLK
timestamp 1698175906
transform 1 0 14896 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__209__CLK
timestamp 1698175906
transform 1 0 24640 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__210__CLK
timestamp 1698175906
transform 1 0 28560 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__211__CLK
timestamp 1698175906
transform 1 0 28112 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__212__CLK
timestamp 1698175906
transform -1 0 26992 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__213__CLK
timestamp 1698175906
transform 1 0 19152 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__214__CLK
timestamp 1698175906
transform -1 0 24752 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__215__CLK
timestamp 1698175906
transform 1 0 27664 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__216__CLK
timestamp 1698175906
transform 1 0 14112 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__217__CLK
timestamp 1698175906
transform 1 0 29232 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__218__CLK
timestamp 1698175906
transform 1 0 26544 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__219__CLK
timestamp 1698175906
transform 1 0 26880 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__220__CLK
timestamp 1698175906
transform 1 0 17472 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__221__CLK
timestamp 1698175906
transform 1 0 13552 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__222__CLK
timestamp 1698175906
transform 1 0 16576 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1698175906
transform 1 0 20496 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19264 0 -1 21952
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1698175906
transform -1 0 22848 0 -1 20384
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1698175906
transform 1 0 23184 0 1 20384
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1568 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698175906
transform 1 0 5376 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698175906
transform 1 0 9184 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698175906
transform 1 0 12992 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_138 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 16800 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_142 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17248 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_172
timestamp 1698175906
transform 1 0 20608 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_176
timestamp 1698175906
transform 1 0 21056 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_232
timestamp 1698175906
transform 1 0 27328 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_236
timestamp 1698175906
transform 1 0 27776 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_240
timestamp 1698175906
transform 1 0 28224 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_274
timestamp 1698175906
transform 1 0 32032 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_308
timestamp 1698175906
transform 1 0 35840 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_342
timestamp 1698175906
transform 1 0 39648 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_346
timestamp 1698175906
transform 1 0 40096 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_348 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 40320 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1568 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698175906
transform 1 0 8736 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698175906
transform 1 0 9408 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698175906
transform 1 0 16576 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_142 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17248 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_150
timestamp 1698175906
transform 1 0 18144 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_154
timestamp 1698175906
transform 1 0 18592 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_156
timestamp 1698175906
transform 1 0 18816 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_183 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21840 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_199
timestamp 1698175906
transform 1 0 23632 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_203
timestamp 1698175906
transform 1 0 24080 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_209
timestamp 1698175906
transform 1 0 24752 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_212
timestamp 1698175906
transform 1 0 25088 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_216
timestamp 1698175906
transform 1 0 25536 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_243
timestamp 1698175906
transform 1 0 28560 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_275
timestamp 1698175906
transform 1 0 32144 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_279
timestamp 1698175906
transform 1 0 32592 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_282
timestamp 1698175906
transform 1 0 32928 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_346
timestamp 1698175906
transform 1 0 40096 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_348
timestamp 1698175906
transform 1 0 40320 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698175906
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698175906
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698175906
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698175906
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_107
timestamp 1698175906
transform 1 0 13328 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_139
timestamp 1698175906
transform 1 0 16912 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_143
timestamp 1698175906
transform 1 0 17360 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_171
timestamp 1698175906
transform 1 0 20496 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_177
timestamp 1698175906
transform 1 0 21168 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_241
timestamp 1698175906
transform 1 0 28336 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698175906
transform 1 0 29008 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698175906
transform 1 0 36176 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_317
timestamp 1698175906
transform 1 0 36848 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698175906
transform 1 0 1568 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698175906
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698175906
transform 1 0 9408 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698175906
transform 1 0 16576 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_142
timestamp 1698175906
transform 1 0 17248 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_206
timestamp 1698175906
transform 1 0 24416 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_212
timestamp 1698175906
transform 1 0 25088 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_276
timestamp 1698175906
transform 1 0 32256 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_282
timestamp 1698175906
transform 1 0 32928 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_346
timestamp 1698175906
transform 1 0 40096 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_348
timestamp 1698175906
transform 1 0 40320 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698175906
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698175906
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698175906
transform 1 0 5488 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698175906
transform 1 0 12656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_107
timestamp 1698175906
transform 1 0 13328 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698175906
transform 1 0 20496 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_177
timestamp 1698175906
transform 1 0 21168 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_241
timestamp 1698175906
transform 1 0 28336 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698175906
transform 1 0 29008 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698175906
transform 1 0 36176 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_317
timestamp 1698175906
transform 1 0 36848 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698175906
transform 1 0 1568 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698175906
transform 1 0 8736 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698175906
transform 1 0 9408 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698175906
transform 1 0 16576 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_142
timestamp 1698175906
transform 1 0 17248 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_206
timestamp 1698175906
transform 1 0 24416 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_212
timestamp 1698175906
transform 1 0 25088 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698175906
transform 1 0 32256 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_282
timestamp 1698175906
transform 1 0 32928 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_346
timestamp 1698175906
transform 1 0 40096 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_348
timestamp 1698175906
transform 1 0 40320 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698175906
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698175906
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698175906
transform 1 0 5488 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698175906
transform 1 0 12656 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_107
timestamp 1698175906
transform 1 0 13328 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_171
timestamp 1698175906
transform 1 0 20496 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_177
timestamp 1698175906
transform 1 0 21168 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_241
timestamp 1698175906
transform 1 0 28336 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_247
timestamp 1698175906
transform 1 0 29008 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_311
timestamp 1698175906
transform 1 0 36176 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_317
timestamp 1698175906
transform 1 0 36848 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698175906
transform 1 0 1568 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698175906
transform 1 0 8736 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_72
timestamp 1698175906
transform 1 0 9408 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698175906
transform 1 0 16576 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_142
timestamp 1698175906
transform 1 0 17248 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_206
timestamp 1698175906
transform 1 0 24416 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_212
timestamp 1698175906
transform 1 0 25088 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_276
timestamp 1698175906
transform 1 0 32256 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_282
timestamp 1698175906
transform 1 0 32928 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_346
timestamp 1698175906
transform 1 0 40096 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_348
timestamp 1698175906
transform 1 0 40320 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698175906
transform 1 0 1568 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698175906
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_37
timestamp 1698175906
transform 1 0 5488 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_101
timestamp 1698175906
transform 1 0 12656 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_107
timestamp 1698175906
transform 1 0 13328 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_171
timestamp 1698175906
transform 1 0 20496 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_177
timestamp 1698175906
transform 1 0 21168 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_241
timestamp 1698175906
transform 1 0 28336 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_247
timestamp 1698175906
transform 1 0 29008 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_311
timestamp 1698175906
transform 1 0 36176 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_317
timestamp 1698175906
transform 1 0 36848 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698175906
transform 1 0 1568 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698175906
transform 1 0 8736 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_72
timestamp 1698175906
transform 1 0 9408 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_136
timestamp 1698175906
transform 1 0 16576 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_142
timestamp 1698175906
transform 1 0 17248 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_206
timestamp 1698175906
transform 1 0 24416 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_212
timestamp 1698175906
transform 1 0 25088 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_276
timestamp 1698175906
transform 1 0 32256 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_282
timestamp 1698175906
transform 1 0 32928 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_346
timestamp 1698175906
transform 1 0 40096 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_348
timestamp 1698175906
transform 1 0 40320 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698175906
transform 1 0 1568 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698175906
transform 1 0 5152 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_37
timestamp 1698175906
transform 1 0 5488 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698175906
transform 1 0 12656 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_107
timestamp 1698175906
transform 1 0 13328 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_171
timestamp 1698175906
transform 1 0 20496 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_177
timestamp 1698175906
transform 1 0 21168 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_241
timestamp 1698175906
transform 1 0 28336 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_247
timestamp 1698175906
transform 1 0 29008 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_311
timestamp 1698175906
transform 1 0 36176 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_317
timestamp 1698175906
transform 1 0 36848 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2
timestamp 1698175906
transform 1 0 1568 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698175906
transform 1 0 8736 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_72
timestamp 1698175906
transform 1 0 9408 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698175906
transform 1 0 16576 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_142
timestamp 1698175906
transform 1 0 17248 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_206
timestamp 1698175906
transform 1 0 24416 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_212
timestamp 1698175906
transform 1 0 25088 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_276
timestamp 1698175906
transform 1 0 32256 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_282
timestamp 1698175906
transform 1 0 32928 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_346
timestamp 1698175906
transform 1 0 40096 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_348
timestamp 1698175906
transform 1 0 40320 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698175906
transform 1 0 1568 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698175906
transform 1 0 5152 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_37
timestamp 1698175906
transform 1 0 5488 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698175906
transform 1 0 12656 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_107
timestamp 1698175906
transform 1 0 13328 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_171
timestamp 1698175906
transform 1 0 20496 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_177
timestamp 1698175906
transform 1 0 21168 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_241
timestamp 1698175906
transform 1 0 28336 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_247
timestamp 1698175906
transform 1 0 29008 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_311
timestamp 1698175906
transform 1 0 36176 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_317
timestamp 1698175906
transform 1 0 36848 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_2
timestamp 1698175906
transform 1 0 1568 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_66
timestamp 1698175906
transform 1 0 8736 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_72
timestamp 1698175906
transform 1 0 9408 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_136
timestamp 1698175906
transform 1 0 16576 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_142
timestamp 1698175906
transform 1 0 17248 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_158
timestamp 1698175906
transform 1 0 19040 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_188
timestamp 1698175906
transform 1 0 22400 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_192
timestamp 1698175906
transform 1 0 22848 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_208
timestamp 1698175906
transform 1 0 24640 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_212
timestamp 1698175906
transform 1 0 25088 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_276
timestamp 1698175906
transform 1 0 32256 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_282
timestamp 1698175906
transform 1 0 32928 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_346
timestamp 1698175906
transform 1 0 40096 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_348
timestamp 1698175906
transform 1 0 40320 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698175906
transform 1 0 1568 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698175906
transform 1 0 5152 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_37
timestamp 1698175906
transform 1 0 5488 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_101
timestamp 1698175906
transform 1 0 12656 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_107
timestamp 1698175906
transform 1 0 13328 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_123
timestamp 1698175906
transform 1 0 15120 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_127
timestamp 1698175906
transform 1 0 15568 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_157
timestamp 1698175906
transform 1 0 18928 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_161
timestamp 1698175906
transform 1 0 19376 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_169
timestamp 1698175906
transform 1 0 20272 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_173
timestamp 1698175906
transform 1 0 20720 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_177
timestamp 1698175906
transform 1 0 21168 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_193
timestamp 1698175906
transform 1 0 22960 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_195
timestamp 1698175906
transform 1 0 23184 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_225
timestamp 1698175906
transform 1 0 26544 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_229
timestamp 1698175906
transform 1 0 26992 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_247
timestamp 1698175906
transform 1 0 29008 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_311
timestamp 1698175906
transform 1 0 36176 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_317
timestamp 1698175906
transform 1 0 36848 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_2
timestamp 1698175906
transform 1 0 1568 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_66
timestamp 1698175906
transform 1 0 8736 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_72
timestamp 1698175906
transform 1 0 9408 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_136
timestamp 1698175906
transform 1 0 16576 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_148
timestamp 1698175906
transform 1 0 17920 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_150
timestamp 1698175906
transform 1 0 18144 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_157
timestamp 1698175906
transform 1 0 18928 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_165
timestamp 1698175906
transform 1 0 19824 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_173
timestamp 1698175906
transform 1 0 20720 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_205
timestamp 1698175906
transform 1 0 24304 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_209
timestamp 1698175906
transform 1 0 24752 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_212
timestamp 1698175906
transform 1 0 25088 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_220
timestamp 1698175906
transform 1 0 25984 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_236
timestamp 1698175906
transform 1 0 27776 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_268
timestamp 1698175906
transform 1 0 31360 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_276
timestamp 1698175906
transform 1 0 32256 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_282
timestamp 1698175906
transform 1 0 32928 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_346
timestamp 1698175906
transform 1 0 40096 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_348
timestamp 1698175906
transform 1 0 40320 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_2
timestamp 1698175906
transform 1 0 1568 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698175906
transform 1 0 5152 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_37
timestamp 1698175906
transform 1 0 5488 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_101
timestamp 1698175906
transform 1 0 12656 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_107
timestamp 1698175906
transform 1 0 13328 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_139
timestamp 1698175906
transform 1 0 16912 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_147
timestamp 1698175906
transform 1 0 17808 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_155
timestamp 1698175906
transform 1 0 18704 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_177
timestamp 1698175906
transform 1 0 21168 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_184
timestamp 1698175906
transform 1 0 21952 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_200
timestamp 1698175906
transform 1 0 23744 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_247
timestamp 1698175906
transform 1 0 29008 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_251
timestamp 1698175906
transform 1 0 29456 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_317
timestamp 1698175906
transform 1 0 36848 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_2
timestamp 1698175906
transform 1 0 1568 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_66
timestamp 1698175906
transform 1 0 8736 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_72
timestamp 1698175906
transform 1 0 9408 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_104
timestamp 1698175906
transform 1 0 12992 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_108
timestamp 1698175906
transform 1 0 13440 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_110
timestamp 1698175906
transform 1 0 13664 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_142
timestamp 1698175906
transform 1 0 17248 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_146
timestamp 1698175906
transform 1 0 17696 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_150
timestamp 1698175906
transform 1 0 18144 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_152
timestamp 1698175906
transform 1 0 18368 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_171
timestamp 1698175906
transform 1 0 20496 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_175
timestamp 1698175906
transform 1 0 20944 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_206
timestamp 1698175906
transform 1 0 24416 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_212
timestamp 1698175906
transform 1 0 25088 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_259
timestamp 1698175906
transform 1 0 30352 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_275
timestamp 1698175906
transform 1 0 32144 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_279
timestamp 1698175906
transform 1 0 32592 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_282
timestamp 1698175906
transform 1 0 32928 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_314
timestamp 1698175906
transform 1 0 36512 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_322
timestamp 1698175906
transform 1 0 37408 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_2
timestamp 1698175906
transform 1 0 1568 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698175906
transform 1 0 5152 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_37
timestamp 1698175906
transform 1 0 5488 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_101
timestamp 1698175906
transform 1 0 12656 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_150
timestamp 1698175906
transform 1 0 18144 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_177
timestamp 1698175906
transform 1 0 21168 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_189
timestamp 1698175906
transform 1 0 22512 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_204
timestamp 1698175906
transform 1 0 24192 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_220
timestamp 1698175906
transform 1 0 25984 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_228
timestamp 1698175906
transform 1 0 26880 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_230
timestamp 1698175906
transform 1 0 27104 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_240
timestamp 1698175906
transform 1 0 28224 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_244
timestamp 1698175906
transform 1 0 28672 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_251
timestamp 1698175906
transform 1 0 29456 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_317
timestamp 1698175906
transform 1 0 36848 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_321
timestamp 1698175906
transform 1 0 37296 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_28
timestamp 1698175906
transform 1 0 4480 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_60
timestamp 1698175906
transform 1 0 8064 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_68
timestamp 1698175906
transform 1 0 8960 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_72
timestamp 1698175906
transform 1 0 9408 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_80
timestamp 1698175906
transform 1 0 10304 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_84
timestamp 1698175906
transform 1 0 10752 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_114
timestamp 1698175906
transform 1 0 14112 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_131
timestamp 1698175906
transform 1 0 16016 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_135
timestamp 1698175906
transform 1 0 16464 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_138
timestamp 1698175906
transform 1 0 16800 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_147
timestamp 1698175906
transform 1 0 17808 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_201
timestamp 1698175906
transform 1 0 23856 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_209
timestamp 1698175906
transform 1 0 24752 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_218
timestamp 1698175906
transform 1 0 25760 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_250
timestamp 1698175906
transform 1 0 29344 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_266
timestamp 1698175906
transform 1 0 31136 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_274
timestamp 1698175906
transform 1 0 32032 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_278
timestamp 1698175906
transform 1 0 32480 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_282
timestamp 1698175906
transform 1 0 32928 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_346
timestamp 1698175906
transform 1 0 40096 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_348
timestamp 1698175906
transform 1 0 40320 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_28
timestamp 1698175906
transform 1 0 4480 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_32
timestamp 1698175906
transform 1 0 4928 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698175906
transform 1 0 5152 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_37
timestamp 1698175906
transform 1 0 5488 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_101
timestamp 1698175906
transform 1 0 12656 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_124
timestamp 1698175906
transform 1 0 15232 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_128
timestamp 1698175906
transform 1 0 15680 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_141
timestamp 1698175906
transform 1 0 17136 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_161
timestamp 1698175906
transform 1 0 19376 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_171
timestamp 1698175906
transform 1 0 20496 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_190
timestamp 1698175906
transform 1 0 22624 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_198
timestamp 1698175906
transform 1 0 23520 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_202
timestamp 1698175906
transform 1 0 23968 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_233
timestamp 1698175906
transform 1 0 27440 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_237
timestamp 1698175906
transform 1 0 27888 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_244
timestamp 1698175906
transform 1 0 28672 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_247
timestamp 1698175906
transform 1 0 29008 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_311
timestamp 1698175906
transform 1 0 36176 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_317
timestamp 1698175906
transform 1 0 36848 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_2
timestamp 1698175906
transform 1 0 1568 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_66
timestamp 1698175906
transform 1 0 8736 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_72
timestamp 1698175906
transform 1 0 9408 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_104
timestamp 1698175906
transform 1 0 12992 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_112
timestamp 1698175906
transform 1 0 13888 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_116
timestamp 1698175906
transform 1 0 14336 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_130
timestamp 1698175906
transform 1 0 15904 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_138
timestamp 1698175906
transform 1 0 16800 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_197
timestamp 1698175906
transform 1 0 23408 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_199
timestamp 1698175906
transform 1 0 23632 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_229
timestamp 1698175906
transform 1 0 26992 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_231
timestamp 1698175906
transform 1 0 27216 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_263
timestamp 1698175906
transform 1 0 30800 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_279
timestamp 1698175906
transform 1 0 32592 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_282
timestamp 1698175906
transform 1 0 32928 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_314
timestamp 1698175906
transform 1 0 36512 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_322
timestamp 1698175906
transform 1 0 37408 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_2
timestamp 1698175906
transform 1 0 1568 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698175906
transform 1 0 5152 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_37
timestamp 1698175906
transform 1 0 5488 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_69
timestamp 1698175906
transform 1 0 9072 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_73
timestamp 1698175906
transform 1 0 9520 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_75
timestamp 1698175906
transform 1 0 9744 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_107
timestamp 1698175906
transform 1 0 13328 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_111
timestamp 1698175906
transform 1 0 13776 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_130
timestamp 1698175906
transform 1 0 15904 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_134
timestamp 1698175906
transform 1 0 16352 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_136
timestamp 1698175906
transform 1 0 16576 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_169
timestamp 1698175906
transform 1 0 20272 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_173
timestamp 1698175906
transform 1 0 20720 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_193
timestamp 1698175906
transform 1 0 22960 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_264
timestamp 1698175906
transform 1 0 30912 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_296
timestamp 1698175906
transform 1 0 34496 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_312
timestamp 1698175906
transform 1 0 36288 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_314
timestamp 1698175906
transform 1 0 36512 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_317
timestamp 1698175906
transform 1 0 36848 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_321
timestamp 1698175906
transform 1 0 37296 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_28
timestamp 1698175906
transform 1 0 4480 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_60
timestamp 1698175906
transform 1 0 8064 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_68
timestamp 1698175906
transform 1 0 8960 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_72
timestamp 1698175906
transform 1 0 9408 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_88
timestamp 1698175906
transform 1 0 11200 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_119
timestamp 1698175906
transform 1 0 14672 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_123
timestamp 1698175906
transform 1 0 15120 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_125
timestamp 1698175906
transform 1 0 15344 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_148
timestamp 1698175906
transform 1 0 17920 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_157
timestamp 1698175906
transform 1 0 18928 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_159
timestamp 1698175906
transform 1 0 19152 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_270
timestamp 1698175906
transform 1 0 31584 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_278
timestamp 1698175906
transform 1 0 32480 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_282
timestamp 1698175906
transform 1 0 32928 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_314
timestamp 1698175906
transform 1 0 36512 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_322
timestamp 1698175906
transform 1 0 37408 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_2
timestamp 1698175906
transform 1 0 1568 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698175906
transform 1 0 5152 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_37
timestamp 1698175906
transform 1 0 5488 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_101
timestamp 1698175906
transform 1 0 12656 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_115
timestamp 1698175906
transform 1 0 14224 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_123
timestamp 1698175906
transform 1 0 15120 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_133
timestamp 1698175906
transform 1 0 16240 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_140
timestamp 1698175906
transform 1 0 17024 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_173
timestamp 1698175906
transform 1 0 20720 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_195
timestamp 1698175906
transform 1 0 23184 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_206
timestamp 1698175906
transform 1 0 24416 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_238
timestamp 1698175906
transform 1 0 28000 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_241
timestamp 1698175906
transform 1 0 28336 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_252
timestamp 1698175906
transform 1 0 29568 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_284
timestamp 1698175906
transform 1 0 33152 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_300
timestamp 1698175906
transform 1 0 34944 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_308
timestamp 1698175906
transform 1 0 35840 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_312
timestamp 1698175906
transform 1 0 36288 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_314
timestamp 1698175906
transform 1 0 36512 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_317
timestamp 1698175906
transform 1 0 36848 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_321
timestamp 1698175906
transform 1 0 37296 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_2
timestamp 1698175906
transform 1 0 1568 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_66
timestamp 1698175906
transform 1 0 8736 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_72
timestamp 1698175906
transform 1 0 9408 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_88
timestamp 1698175906
transform 1 0 11200 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_125
timestamp 1698175906
transform 1 0 15344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_127
timestamp 1698175906
transform 1 0 15568 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_136
timestamp 1698175906
transform 1 0 16576 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_142
timestamp 1698175906
transform 1 0 17248 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_174
timestamp 1698175906
transform 1 0 20832 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_176
timestamp 1698175906
transform 1 0 21056 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_195
timestamp 1698175906
transform 1 0 23184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_205
timestamp 1698175906
transform 1 0 24304 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_209
timestamp 1698175906
transform 1 0 24752 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_212
timestamp 1698175906
transform 1 0 25088 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_220
timestamp 1698175906
transform 1 0 25984 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_224
timestamp 1698175906
transform 1 0 26432 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_256
timestamp 1698175906
transform 1 0 30016 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_260
timestamp 1698175906
transform 1 0 30464 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_276
timestamp 1698175906
transform 1 0 32256 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_282
timestamp 1698175906
transform 1 0 32928 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_314
timestamp 1698175906
transform 1 0 36512 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_322
timestamp 1698175906
transform 1 0 37408 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_2
timestamp 1698175906
transform 1 0 1568 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698175906
transform 1 0 5152 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_37
timestamp 1698175906
transform 1 0 5488 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_101
timestamp 1698175906
transform 1 0 12656 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_117
timestamp 1698175906
transform 1 0 14448 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_127
timestamp 1698175906
transform 1 0 15568 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_143
timestamp 1698175906
transform 1 0 17360 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_167
timestamp 1698175906
transform 1 0 20048 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_183
timestamp 1698175906
transform 1 0 21840 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_187
timestamp 1698175906
transform 1 0 22288 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_242
timestamp 1698175906
transform 1 0 28448 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_244
timestamp 1698175906
transform 1 0 28672 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_247
timestamp 1698175906
transform 1 0 29008 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_311
timestamp 1698175906
transform 1 0 36176 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_317
timestamp 1698175906
transform 1 0 36848 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_321
timestamp 1698175906
transform 1 0 37296 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_2
timestamp 1698175906
transform 1 0 1568 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_66
timestamp 1698175906
transform 1 0 8736 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_72
timestamp 1698175906
transform 1 0 9408 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_136
timestamp 1698175906
transform 1 0 16576 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_156
timestamp 1698175906
transform 1 0 18816 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_172
timestamp 1698175906
transform 1 0 20608 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_180
timestamp 1698175906
transform 1 0 21504 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_212
timestamp 1698175906
transform 1 0 25088 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_216
timestamp 1698175906
transform 1 0 25536 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_282
timestamp 1698175906
transform 1 0 32928 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_314
timestamp 1698175906
transform 1 0 36512 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_322
timestamp 1698175906
transform 1 0 37408 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_2
timestamp 1698175906
transform 1 0 1568 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698175906
transform 1 0 5152 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_37
timestamp 1698175906
transform 1 0 5488 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_101
timestamp 1698175906
transform 1 0 12656 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_107
timestamp 1698175906
transform 1 0 13328 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_120
timestamp 1698175906
transform 1 0 14784 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_162
timestamp 1698175906
transform 1 0 19488 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_166
timestamp 1698175906
transform 1 0 19936 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_174
timestamp 1698175906
transform 1 0 20832 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_183
timestamp 1698175906
transform 1 0 21840 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_215
timestamp 1698175906
transform 1 0 25424 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_231
timestamp 1698175906
transform 1 0 27216 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_239
timestamp 1698175906
transform 1 0 28112 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_243
timestamp 1698175906
transform 1 0 28560 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_247
timestamp 1698175906
transform 1 0 29008 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_311
timestamp 1698175906
transform 1 0 36176 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_317
timestamp 1698175906
transform 1 0 36848 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_28
timestamp 1698175906
transform 1 0 4480 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_60
timestamp 1698175906
transform 1 0 8064 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_68
timestamp 1698175906
transform 1 0 8960 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_72
timestamp 1698175906
transform 1 0 9408 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_88
timestamp 1698175906
transform 1 0 11200 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_130
timestamp 1698175906
transform 1 0 15904 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_138
timestamp 1698175906
transform 1 0 16800 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_142
timestamp 1698175906
transform 1 0 17248 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_150
timestamp 1698175906
transform 1 0 18144 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_152
timestamp 1698175906
transform 1 0 18368 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_157
timestamp 1698175906
transform 1 0 18928 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_165
timestamp 1698175906
transform 1 0 19824 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_174
timestamp 1698175906
transform 1 0 20832 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_178
timestamp 1698175906
transform 1 0 21280 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_212
timestamp 1698175906
transform 1 0 25088 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_276
timestamp 1698175906
transform 1 0 32256 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_282
timestamp 1698175906
transform 1 0 32928 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_346
timestamp 1698175906
transform 1 0 40096 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_348
timestamp 1698175906
transform 1 0 40320 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_28
timestamp 1698175906
transform 1 0 4480 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_32
timestamp 1698175906
transform 1 0 4928 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698175906
transform 1 0 5152 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_37
timestamp 1698175906
transform 1 0 5488 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_101
timestamp 1698175906
transform 1 0 12656 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_115
timestamp 1698175906
transform 1 0 14224 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_119
timestamp 1698175906
transform 1 0 14672 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_123
timestamp 1698175906
transform 1 0 15120 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_131
timestamp 1698175906
transform 1 0 16016 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_135
timestamp 1698175906
transform 1 0 16464 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_137
timestamp 1698175906
transform 1 0 16688 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_190
timestamp 1698175906
transform 1 0 22624 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_222
timestamp 1698175906
transform 1 0 26208 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_238
timestamp 1698175906
transform 1 0 28000 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_242
timestamp 1698175906
transform 1 0 28448 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_244
timestamp 1698175906
transform 1 0 28672 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_247
timestamp 1698175906
transform 1 0 29008 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_311
timestamp 1698175906
transform 1 0 36176 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_317
timestamp 1698175906
transform 1 0 36848 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_333
timestamp 1698175906
transform 1 0 38640 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_341
timestamp 1698175906
transform 1 0 39536 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_2
timestamp 1698175906
transform 1 0 1568 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_66
timestamp 1698175906
transform 1 0 8736 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_72
timestamp 1698175906
transform 1 0 9408 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_88
timestamp 1698175906
transform 1 0 11200 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_118
timestamp 1698175906
transform 1 0 14560 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_122
timestamp 1698175906
transform 1 0 15008 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_138
timestamp 1698175906
transform 1 0 16800 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_142
timestamp 1698175906
transform 1 0 17248 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_150
timestamp 1698175906
transform 1 0 18144 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_154
timestamp 1698175906
transform 1 0 18592 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_156
timestamp 1698175906
transform 1 0 18816 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_205
timestamp 1698175906
transform 1 0 24304 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_209
timestamp 1698175906
transform 1 0 24752 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_212
timestamp 1698175906
transform 1 0 25088 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_276
timestamp 1698175906
transform 1 0 32256 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_282
timestamp 1698175906
transform 1 0 32928 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_346
timestamp 1698175906
transform 1 0 40096 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_348
timestamp 1698175906
transform 1 0 40320 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_2
timestamp 1698175906
transform 1 0 1568 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698175906
transform 1 0 5152 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_37
timestamp 1698175906
transform 1 0 5488 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_101
timestamp 1698175906
transform 1 0 12656 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_107
timestamp 1698175906
transform 1 0 13328 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_139
timestamp 1698175906
transform 1 0 16912 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_143
timestamp 1698175906
transform 1 0 17360 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_145
timestamp 1698175906
transform 1 0 17584 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_177
timestamp 1698175906
transform 1 0 21168 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_181
timestamp 1698175906
transform 1 0 21616 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_247
timestamp 1698175906
transform 1 0 29008 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_311
timestamp 1698175906
transform 1 0 36176 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_317
timestamp 1698175906
transform 1 0 36848 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_2
timestamp 1698175906
transform 1 0 1568 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_66
timestamp 1698175906
transform 1 0 8736 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_72
timestamp 1698175906
transform 1 0 9408 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_136
timestamp 1698175906
transform 1 0 16576 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_142
timestamp 1698175906
transform 1 0 17248 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_206
timestamp 1698175906
transform 1 0 24416 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_212
timestamp 1698175906
transform 1 0 25088 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_276
timestamp 1698175906
transform 1 0 32256 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_282
timestamp 1698175906
transform 1 0 32928 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_346
timestamp 1698175906
transform 1 0 40096 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_348
timestamp 1698175906
transform 1 0 40320 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698175906
transform 1 0 1568 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698175906
transform 1 0 5152 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_37
timestamp 1698175906
transform 1 0 5488 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_101
timestamp 1698175906
transform 1 0 12656 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_107
timestamp 1698175906
transform 1 0 13328 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_171
timestamp 1698175906
transform 1 0 20496 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_177
timestamp 1698175906
transform 1 0 21168 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_241
timestamp 1698175906
transform 1 0 28336 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_247
timestamp 1698175906
transform 1 0 29008 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_311
timestamp 1698175906
transform 1 0 36176 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_317
timestamp 1698175906
transform 1 0 36848 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2
timestamp 1698175906
transform 1 0 1568 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_66
timestamp 1698175906
transform 1 0 8736 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_72
timestamp 1698175906
transform 1 0 9408 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_136
timestamp 1698175906
transform 1 0 16576 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_142
timestamp 1698175906
transform 1 0 17248 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_206
timestamp 1698175906
transform 1 0 24416 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_212
timestamp 1698175906
transform 1 0 25088 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_276
timestamp 1698175906
transform 1 0 32256 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_282
timestamp 1698175906
transform 1 0 32928 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_346
timestamp 1698175906
transform 1 0 40096 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_348
timestamp 1698175906
transform 1 0 40320 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_2
timestamp 1698175906
transform 1 0 1568 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698175906
transform 1 0 5152 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_37
timestamp 1698175906
transform 1 0 5488 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_101
timestamp 1698175906
transform 1 0 12656 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_107
timestamp 1698175906
transform 1 0 13328 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_171
timestamp 1698175906
transform 1 0 20496 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_177
timestamp 1698175906
transform 1 0 21168 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_241
timestamp 1698175906
transform 1 0 28336 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_247
timestamp 1698175906
transform 1 0 29008 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_311
timestamp 1698175906
transform 1 0 36176 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_317
timestamp 1698175906
transform 1 0 36848 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2
timestamp 1698175906
transform 1 0 1568 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_66
timestamp 1698175906
transform 1 0 8736 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_72
timestamp 1698175906
transform 1 0 9408 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_136
timestamp 1698175906
transform 1 0 16576 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_142
timestamp 1698175906
transform 1 0 17248 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_206
timestamp 1698175906
transform 1 0 24416 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_212
timestamp 1698175906
transform 1 0 25088 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_276
timestamp 1698175906
transform 1 0 32256 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_282
timestamp 1698175906
transform 1 0 32928 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_346
timestamp 1698175906
transform 1 0 40096 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_348
timestamp 1698175906
transform 1 0 40320 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698175906
transform 1 0 1568 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698175906
transform 1 0 5152 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_37
timestamp 1698175906
transform 1 0 5488 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_101
timestamp 1698175906
transform 1 0 12656 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_107
timestamp 1698175906
transform 1 0 13328 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_171
timestamp 1698175906
transform 1 0 20496 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_177
timestamp 1698175906
transform 1 0 21168 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_241
timestamp 1698175906
transform 1 0 28336 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_247
timestamp 1698175906
transform 1 0 29008 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_311
timestamp 1698175906
transform 1 0 36176 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_317
timestamp 1698175906
transform 1 0 36848 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_2
timestamp 1698175906
transform 1 0 1568 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_66
timestamp 1698175906
transform 1 0 8736 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_72
timestamp 1698175906
transform 1 0 9408 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_136
timestamp 1698175906
transform 1 0 16576 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_142
timestamp 1698175906
transform 1 0 17248 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_206
timestamp 1698175906
transform 1 0 24416 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_212
timestamp 1698175906
transform 1 0 25088 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_276
timestamp 1698175906
transform 1 0 32256 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_282
timestamp 1698175906
transform 1 0 32928 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_346
timestamp 1698175906
transform 1 0 40096 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_348
timestamp 1698175906
transform 1 0 40320 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698175906
transform 1 0 1568 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698175906
transform 1 0 5152 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_37
timestamp 1698175906
transform 1 0 5488 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_101
timestamp 1698175906
transform 1 0 12656 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_107
timestamp 1698175906
transform 1 0 13328 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_171
timestamp 1698175906
transform 1 0 20496 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_177
timestamp 1698175906
transform 1 0 21168 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_241
timestamp 1698175906
transform 1 0 28336 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_247
timestamp 1698175906
transform 1 0 29008 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_311
timestamp 1698175906
transform 1 0 36176 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_317
timestamp 1698175906
transform 1 0 36848 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2
timestamp 1698175906
transform 1 0 1568 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1698175906
transform 1 0 8736 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_72
timestamp 1698175906
transform 1 0 9408 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_136
timestamp 1698175906
transform 1 0 16576 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_142
timestamp 1698175906
transform 1 0 17248 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_206
timestamp 1698175906
transform 1 0 24416 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_212
timestamp 1698175906
transform 1 0 25088 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_276
timestamp 1698175906
transform 1 0 32256 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_282
timestamp 1698175906
transform 1 0 32928 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_346
timestamp 1698175906
transform 1 0 40096 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_348
timestamp 1698175906
transform 1 0 40320 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_2
timestamp 1698175906
transform 1 0 1568 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698175906
transform 1 0 5152 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_37
timestamp 1698175906
transform 1 0 5488 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_101
timestamp 1698175906
transform 1 0 12656 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_107
timestamp 1698175906
transform 1 0 13328 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_171
timestamp 1698175906
transform 1 0 20496 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_177
timestamp 1698175906
transform 1 0 21168 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_241
timestamp 1698175906
transform 1 0 28336 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_247
timestamp 1698175906
transform 1 0 29008 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_311
timestamp 1698175906
transform 1 0 36176 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_317
timestamp 1698175906
transform 1 0 36848 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_2
timestamp 1698175906
transform 1 0 1568 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_66
timestamp 1698175906
transform 1 0 8736 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_72
timestamp 1698175906
transform 1 0 9408 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_136
timestamp 1698175906
transform 1 0 16576 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_142
timestamp 1698175906
transform 1 0 17248 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_174
timestamp 1698175906
transform 1 0 20832 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_201
timestamp 1698175906
transform 1 0 23856 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_209
timestamp 1698175906
transform 1 0 24752 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_212
timestamp 1698175906
transform 1 0 25088 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_276
timestamp 1698175906
transform 1 0 32256 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_282
timestamp 1698175906
transform 1 0 32928 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_346
timestamp 1698175906
transform 1 0 40096 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_348
timestamp 1698175906
transform 1 0 40320 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_2
timestamp 1698175906
transform 1 0 1568 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_36
timestamp 1698175906
transform 1 0 5376 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_70
timestamp 1698175906
transform 1 0 9184 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_104
timestamp 1698175906
transform 1 0 12992 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_138
timestamp 1698175906
transform 1 0 16800 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_142
timestamp 1698175906
transform 1 0 17248 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_172
timestamp 1698175906
transform 1 0 20608 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_176
timestamp 1698175906
transform 1 0 21056 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_232
timestamp 1698175906
transform 1 0 27328 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_236
timestamp 1698175906
transform 1 0 27776 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_240
timestamp 1698175906
transform 1 0 28224 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_274
timestamp 1698175906
transform 1 0 32032 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_308
timestamp 1698175906
transform 1 0 35840 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_342
timestamp 1698175906
transform 1 0 39648 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_346
timestamp 1698175906
transform 1 0 40096 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_348
timestamp 1698175906
transform 1 0 40320 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita9_25 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 24752 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  ita9_26 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 39984 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 37520 0 1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output2
timestamp 1698175906
transform 1 0 37520 0 1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output3
timestamp 1698175906
transform 1 0 37520 0 -1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output4
timestamp 1698175906
transform 1 0 25648 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output5
timestamp 1698175906
transform 1 0 18928 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output6
timestamp 1698175906
transform -1 0 24192 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output7
timestamp 1698175906
transform 1 0 37520 0 -1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output8
timestamp 1698175906
transform -1 0 20384 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output9
timestamp 1698175906
transform 1 0 37520 0 1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output10
timestamp 1698175906
transform 1 0 24416 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output11
timestamp 1698175906
transform 1 0 17584 0 1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output12
timestamp 1698175906
transform -1 0 4480 0 -1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output13
timestamp 1698175906
transform -1 0 4480 0 -1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output14
timestamp 1698175906
transform -1 0 4480 0 1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output15
timestamp 1698175906
transform 1 0 37520 0 -1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output16
timestamp 1698175906
transform -1 0 20384 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output17
timestamp 1698175906
transform 1 0 24416 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output18
timestamp 1698175906
transform 1 0 20944 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output19
timestamp 1698175906
transform 1 0 37520 0 1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output20
timestamp 1698175906
transform 1 0 21280 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output21
timestamp 1698175906
transform 1 0 37520 0 -1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output22
timestamp 1698175906
transform 1 0 37520 0 -1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output23
timestamp 1698175906
transform -1 0 4480 0 1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output24
timestamp 1698175906
transform -1 0 4480 0 -1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_45 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698175906
transform -1 0 40656 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_46
timestamp 1698175906
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698175906
transform -1 0 40656 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_47
timestamp 1698175906
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698175906
transform -1 0 40656 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_48
timestamp 1698175906
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698175906
transform -1 0 40656 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_49
timestamp 1698175906
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698175906
transform -1 0 40656 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_50
timestamp 1698175906
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698175906
transform -1 0 40656 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_51
timestamp 1698175906
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698175906
transform -1 0 40656 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_52
timestamp 1698175906
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698175906
transform -1 0 40656 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_53
timestamp 1698175906
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698175906
transform -1 0 40656 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_54
timestamp 1698175906
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698175906
transform -1 0 40656 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_55
timestamp 1698175906
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698175906
transform -1 0 40656 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_56
timestamp 1698175906
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698175906
transform -1 0 40656 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_57
timestamp 1698175906
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698175906
transform -1 0 40656 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_58
timestamp 1698175906
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698175906
transform -1 0 40656 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_59
timestamp 1698175906
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698175906
transform -1 0 40656 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_60
timestamp 1698175906
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698175906
transform -1 0 40656 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_61
timestamp 1698175906
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698175906
transform -1 0 40656 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_62
timestamp 1698175906
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698175906
transform -1 0 40656 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_63
timestamp 1698175906
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698175906
transform -1 0 40656 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_64
timestamp 1698175906
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698175906
transform -1 0 40656 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_65
timestamp 1698175906
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698175906
transform -1 0 40656 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_66
timestamp 1698175906
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698175906
transform -1 0 40656 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_67
timestamp 1698175906
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698175906
transform -1 0 40656 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_68
timestamp 1698175906
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698175906
transform -1 0 40656 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_69
timestamp 1698175906
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698175906
transform -1 0 40656 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_70
timestamp 1698175906
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698175906
transform -1 0 40656 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_71
timestamp 1698175906
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698175906
transform -1 0 40656 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_72
timestamp 1698175906
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698175906
transform -1 0 40656 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_73
timestamp 1698175906
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698175906
transform -1 0 40656 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_74
timestamp 1698175906
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698175906
transform -1 0 40656 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_75
timestamp 1698175906
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698175906
transform -1 0 40656 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_76
timestamp 1698175906
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698175906
transform -1 0 40656 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_77
timestamp 1698175906
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698175906
transform -1 0 40656 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_78
timestamp 1698175906
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698175906
transform -1 0 40656 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_79
timestamp 1698175906
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698175906
transform -1 0 40656 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_80
timestamp 1698175906
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698175906
transform -1 0 40656 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_81
timestamp 1698175906
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698175906
transform -1 0 40656 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_82
timestamp 1698175906
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698175906
transform -1 0 40656 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_83
timestamp 1698175906
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698175906
transform -1 0 40656 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_84
timestamp 1698175906
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698175906
transform -1 0 40656 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_85
timestamp 1698175906
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698175906
transform -1 0 40656 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_86
timestamp 1698175906
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698175906
transform -1 0 40656 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_87
timestamp 1698175906
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698175906
transform -1 0 40656 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_88
timestamp 1698175906
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698175906
transform -1 0 40656 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_89
timestamp 1698175906
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698175906
transform -1 0 40656 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_90 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_91
timestamp 1698175906
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_92
timestamp 1698175906
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_93
timestamp 1698175906
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_94
timestamp 1698175906
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_95
timestamp 1698175906
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_96
timestamp 1698175906
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_97
timestamp 1698175906
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_98
timestamp 1698175906
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_99
timestamp 1698175906
transform 1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_100
timestamp 1698175906
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_101
timestamp 1698175906
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_102
timestamp 1698175906
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_103
timestamp 1698175906
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_104
timestamp 1698175906
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_105
timestamp 1698175906
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_106
timestamp 1698175906
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_107
timestamp 1698175906
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_108
timestamp 1698175906
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_109
timestamp 1698175906
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_110
timestamp 1698175906
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_111
timestamp 1698175906
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_112
timestamp 1698175906
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_113
timestamp 1698175906
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_114
timestamp 1698175906
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_115
timestamp 1698175906
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_116
timestamp 1698175906
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_117
timestamp 1698175906
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_118
timestamp 1698175906
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_119
timestamp 1698175906
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_120
timestamp 1698175906
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_121
timestamp 1698175906
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_122
timestamp 1698175906
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_123
timestamp 1698175906
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_124
timestamp 1698175906
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_125
timestamp 1698175906
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_126
timestamp 1698175906
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_127
timestamp 1698175906
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_128
timestamp 1698175906
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_129
timestamp 1698175906
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_130
timestamp 1698175906
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_131
timestamp 1698175906
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_132
timestamp 1698175906
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_133
timestamp 1698175906
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_134
timestamp 1698175906
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_135
timestamp 1698175906
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_136
timestamp 1698175906
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_137
timestamp 1698175906
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_138
timestamp 1698175906
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_139
timestamp 1698175906
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_140
timestamp 1698175906
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_141
timestamp 1698175906
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_142
timestamp 1698175906
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_143
timestamp 1698175906
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_144
timestamp 1698175906
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_145
timestamp 1698175906
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_146
timestamp 1698175906
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_147
timestamp 1698175906
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_148
timestamp 1698175906
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_149
timestamp 1698175906
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_150
timestamp 1698175906
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_151
timestamp 1698175906
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_152
timestamp 1698175906
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_153
timestamp 1698175906
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_154
timestamp 1698175906
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_155
timestamp 1698175906
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_156
timestamp 1698175906
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_157
timestamp 1698175906
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_158
timestamp 1698175906
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_159
timestamp 1698175906
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_160
timestamp 1698175906
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_161
timestamp 1698175906
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_162
timestamp 1698175906
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_163
timestamp 1698175906
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_164
timestamp 1698175906
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_165
timestamp 1698175906
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_166
timestamp 1698175906
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_167
timestamp 1698175906
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_168
timestamp 1698175906
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_169
timestamp 1698175906
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_170
timestamp 1698175906
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_171
timestamp 1698175906
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_172
timestamp 1698175906
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_173
timestamp 1698175906
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_174
timestamp 1698175906
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_175
timestamp 1698175906
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_176
timestamp 1698175906
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_177
timestamp 1698175906
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_178
timestamp 1698175906
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_179
timestamp 1698175906
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_180
timestamp 1698175906
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_181
timestamp 1698175906
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_182
timestamp 1698175906
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_183
timestamp 1698175906
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_184
timestamp 1698175906
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_185
timestamp 1698175906
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_186
timestamp 1698175906
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_187
timestamp 1698175906
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_188
timestamp 1698175906
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_189
timestamp 1698175906
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_190
timestamp 1698175906
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_191
timestamp 1698175906
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_192
timestamp 1698175906
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_193
timestamp 1698175906
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_194
timestamp 1698175906
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_195
timestamp 1698175906
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_196
timestamp 1698175906
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_197
timestamp 1698175906
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_198
timestamp 1698175906
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_199
timestamp 1698175906
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_200
timestamp 1698175906
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_201
timestamp 1698175906
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_202
timestamp 1698175906
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_203
timestamp 1698175906
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_204
timestamp 1698175906
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_205
timestamp 1698175906
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_206
timestamp 1698175906
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_207
timestamp 1698175906
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_208
timestamp 1698175906
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_209
timestamp 1698175906
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_210
timestamp 1698175906
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_211
timestamp 1698175906
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_212
timestamp 1698175906
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_213
timestamp 1698175906
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_214
timestamp 1698175906
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_215
timestamp 1698175906
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_216
timestamp 1698175906
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_217
timestamp 1698175906
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_218
timestamp 1698175906
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_219
timestamp 1698175906
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_220
timestamp 1698175906
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_221
timestamp 1698175906
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_222
timestamp 1698175906
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_223
timestamp 1698175906
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_224
timestamp 1698175906
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_225
timestamp 1698175906
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_226
timestamp 1698175906
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_227
timestamp 1698175906
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_228
timestamp 1698175906
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_229
timestamp 1698175906
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_230
timestamp 1698175906
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_231
timestamp 1698175906
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_232
timestamp 1698175906
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_233
timestamp 1698175906
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_234
timestamp 1698175906
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_235
timestamp 1698175906
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_236
timestamp 1698175906
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_237
timestamp 1698175906
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_238
timestamp 1698175906
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_239
timestamp 1698175906
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_240
timestamp 1698175906
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_241
timestamp 1698175906
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_242
timestamp 1698175906
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_243
timestamp 1698175906
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_244
timestamp 1698175906
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_245
timestamp 1698175906
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_246
timestamp 1698175906
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_247
timestamp 1698175906
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_248
timestamp 1698175906
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_249
timestamp 1698175906
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_250
timestamp 1698175906
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_251
timestamp 1698175906
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_252
timestamp 1698175906
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_253
timestamp 1698175906
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_254
timestamp 1698175906
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_255
timestamp 1698175906
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_256
timestamp 1698175906
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_257
timestamp 1698175906
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_258
timestamp 1698175906
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_259
timestamp 1698175906
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_260
timestamp 1698175906
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_261
timestamp 1698175906
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_262
timestamp 1698175906
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_263
timestamp 1698175906
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_264
timestamp 1698175906
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_265
timestamp 1698175906
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_266
timestamp 1698175906
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_267
timestamp 1698175906
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_268
timestamp 1698175906
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_269
timestamp 1698175906
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_270
timestamp 1698175906
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_271
timestamp 1698175906
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_272
timestamp 1698175906
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_273
timestamp 1698175906
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_274
timestamp 1698175906
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_275
timestamp 1698175906
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_276
timestamp 1698175906
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_277
timestamp 1698175906
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_278
timestamp 1698175906
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_279
timestamp 1698175906
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_280
timestamp 1698175906
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_281
timestamp 1698175906
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_282
timestamp 1698175906
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_283
timestamp 1698175906
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_284
timestamp 1698175906
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_285
timestamp 1698175906
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_286
timestamp 1698175906
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_287
timestamp 1698175906
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_288
timestamp 1698175906
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_289
timestamp 1698175906
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_290
timestamp 1698175906
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_291
timestamp 1698175906
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_292
timestamp 1698175906
transform 1 0 32704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_293
timestamp 1698175906
transform 1 0 5152 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_294
timestamp 1698175906
transform 1 0 8960 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_295
timestamp 1698175906
transform 1 0 12768 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_296
timestamp 1698175906
transform 1 0 16576 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_297
timestamp 1698175906
transform 1 0 20384 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_298
timestamp 1698175906
transform 1 0 24192 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_299
timestamp 1698175906
transform 1 0 28000 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_300
timestamp 1698175906
transform 1 0 31808 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_301
timestamp 1698175906
transform 1 0 35616 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_302
timestamp 1698175906
transform 1 0 39424 0 1 37632
box -86 -86 310 870
<< labels >>
flabel metal3 s 0 27552 800 27664 0 FreeSans 448 0 0 0 clk
port 0 nsew signal input
flabel metal3 s 41200 23520 42000 23632 0 FreeSans 448 0 0 0 segm[0]
port 1 nsew signal tristate
flabel metal3 s 41200 21504 42000 21616 0 FreeSans 448 0 0 0 segm[10]
port 2 nsew signal tristate
flabel metal3 s 41200 20832 42000 20944 0 FreeSans 448 0 0 0 segm[11]
port 3 nsew signal tristate
flabel metal2 s 25536 0 25648 800 0 FreeSans 448 90 0 0 segm[12]
port 4 nsew signal tristate
flabel metal3 s 41200 26208 42000 26320 0 FreeSans 448 0 0 0 segm[13]
port 5 nsew signal tristate
flabel metal2 s 18816 0 18928 800 0 FreeSans 448 90 0 0 segm[1]
port 6 nsew signal tristate
flabel metal2 s 22176 41200 22288 42000 0 FreeSans 448 90 0 0 segm[2]
port 7 nsew signal tristate
flabel metal3 s 41200 24192 42000 24304 0 FreeSans 448 0 0 0 segm[3]
port 8 nsew signal tristate
flabel metal2 s 18144 0 18256 800 0 FreeSans 448 90 0 0 segm[4]
port 9 nsew signal tristate
flabel metal2 s 24192 0 24304 800 0 FreeSans 448 90 0 0 segm[5]
port 10 nsew signal tristate
flabel metal3 s 41200 17472 42000 17584 0 FreeSans 448 0 0 0 segm[6]
port 11 nsew signal tristate
flabel metal2 s 23520 0 23632 800 0 FreeSans 448 90 0 0 segm[7]
port 12 nsew signal tristate
flabel metal2 s 17472 0 17584 800 0 FreeSans 448 90 0 0 segm[8]
port 13 nsew signal tristate
flabel metal3 s 0 20832 800 20944 0 FreeSans 448 0 0 0 segm[9]
port 14 nsew signal tristate
flabel metal3 s 0 26880 800 26992 0 FreeSans 448 0 0 0 sel[0]
port 15 nsew signal tristate
flabel metal3 s 0 18816 800 18928 0 FreeSans 448 0 0 0 sel[10]
port 16 nsew signal tristate
flabel metal3 s 41200 16128 42000 16240 0 FreeSans 448 0 0 0 sel[11]
port 17 nsew signal tristate
flabel metal2 s 18144 41200 18256 42000 0 FreeSans 448 90 0 0 sel[1]
port 18 nsew signal tristate
flabel metal2 s 22848 41200 22960 42000 0 FreeSans 448 90 0 0 sel[2]
port 19 nsew signal tristate
flabel metal2 s 20832 41200 20944 42000 0 FreeSans 448 90 0 0 sel[3]
port 20 nsew signal tristate
flabel metal3 s 41200 20160 42000 20272 0 FreeSans 448 0 0 0 sel[4]
port 21 nsew signal tristate
flabel metal2 s 22176 0 22288 800 0 FreeSans 448 90 0 0 sel[5]
port 22 nsew signal tristate
flabel metal3 s 41200 19488 42000 19600 0 FreeSans 448 0 0 0 sel[6]
port 23 nsew signal tristate
flabel metal3 s 41200 22848 42000 22960 0 FreeSans 448 0 0 0 sel[7]
port 24 nsew signal tristate
flabel metal3 s 0 26208 800 26320 0 FreeSans 448 0 0 0 sel[8]
port 25 nsew signal tristate
flabel metal3 s 0 18144 800 18256 0 FreeSans 448 0 0 0 sel[9]
port 26 nsew signal tristate
flabel metal4 s 4448 3076 4768 38476 0 FreeSans 1280 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 35168 3076 35488 38476 0 FreeSans 1280 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 19808 3076 20128 38476 0 FreeSans 1280 90 0 0 vss
port 28 nsew ground bidirectional
rlabel metal1 21000 38416 21000 38416 0 vdd
rlabel metal1 21000 37632 21000 37632 0 vss
rlabel metal2 22064 16968 22064 16968 0 _000_
rlabel metal2 26040 20832 26040 20832 0 _001_
rlabel metal2 29624 21168 29624 21168 0 _002_
rlabel metal2 24304 14616 24304 14616 0 _003_
rlabel metal3 17024 15400 17024 15400 0 _004_
rlabel metal2 21392 27160 21392 27160 0 _005_
rlabel metal2 25200 18312 25200 18312 0 _006_
rlabel metal2 13160 18704 13160 18704 0 _007_
rlabel metal2 26600 15568 26600 15568 0 _008_
rlabel metal2 23688 23576 23688 23576 0 _009_
rlabel metal2 28056 17360 28056 17360 0 _010_
rlabel metal2 14728 17192 14728 17192 0 _011_
rlabel metal2 14280 20832 14280 20832 0 _012_
rlabel metal2 15624 18032 15624 18032 0 _013_
rlabel metal2 27776 23240 27776 23240 0 _014_
rlabel metal2 20160 13832 20160 13832 0 _015_
rlabel metal2 28448 19432 28448 19432 0 _016_
rlabel metal2 13944 27496 13944 27496 0 _017_
rlabel metal3 17472 23464 17472 23464 0 _018_
rlabel metal2 13048 23408 13048 23408 0 _019_
rlabel metal2 12376 21896 12376 21896 0 _020_
rlabel metal2 22680 24304 22680 24304 0 _021_
rlabel metal2 19208 28280 19208 28280 0 _022_
rlabel metal3 16856 24920 16856 24920 0 _023_
rlabel metal2 13888 26376 13888 26376 0 _024_
rlabel metal2 17976 25032 17976 25032 0 _025_
rlabel metal2 13496 26824 13496 26824 0 _026_
rlabel metal3 24584 18648 24584 18648 0 _027_
rlabel metal2 18872 17472 18872 17472 0 _028_
rlabel metal3 21056 17528 21056 17528 0 _029_
rlabel metal2 24696 20272 24696 20272 0 _030_
rlabel metal3 22848 17640 22848 17640 0 _031_
rlabel metal3 25592 20104 25592 20104 0 _032_
rlabel metal2 24472 17024 24472 17024 0 _033_
rlabel metal2 24360 20048 24360 20048 0 _034_
rlabel metal2 23912 21560 23912 21560 0 _035_
rlabel metal3 30072 20776 30072 20776 0 _036_
rlabel metal3 21896 20832 21896 20832 0 _037_
rlabel metal3 28028 20664 28028 20664 0 _038_
rlabel metal2 24920 16184 24920 16184 0 _039_
rlabel metal2 18200 17304 18200 17304 0 _040_
rlabel metal2 18536 16464 18536 16464 0 _041_
rlabel metal2 17752 15960 17752 15960 0 _042_
rlabel metal2 22008 27160 22008 27160 0 _043_
rlabel metal2 25536 18536 25536 18536 0 _044_
rlabel metal2 14392 20356 14392 20356 0 _045_
rlabel metal2 14168 21056 14168 21056 0 _046_
rlabel metal2 15064 18480 15064 18480 0 _047_
rlabel metal3 14392 19096 14392 19096 0 _048_
rlabel metal2 27384 17472 27384 17472 0 _049_
rlabel metal2 27160 15288 27160 15288 0 _050_
rlabel metal2 24248 22792 24248 22792 0 _051_
rlabel metal3 28504 17640 28504 17640 0 _052_
rlabel metal2 17248 17640 17248 17640 0 _053_
rlabel metal2 16856 17584 16856 17584 0 _054_
rlabel metal3 14952 20552 14952 20552 0 _055_
rlabel metal2 14840 21840 14840 21840 0 _056_
rlabel metal3 15064 18424 15064 18424 0 _057_
rlabel metal2 21784 23520 21784 23520 0 _058_
rlabel metal2 17640 22120 17640 22120 0 _059_
rlabel metal2 22512 19096 22512 19096 0 _060_
rlabel metal2 27384 23968 27384 23968 0 _061_
rlabel metal2 29400 22904 29400 22904 0 _062_
rlabel metal2 29064 22848 29064 22848 0 _063_
rlabel metal3 21112 26264 21112 26264 0 _064_
rlabel metal2 19656 22064 19656 22064 0 _065_
rlabel metal2 16408 20384 16408 20384 0 _066_
rlabel metal3 20272 22344 20272 22344 0 _067_
rlabel metal2 23240 23856 23240 23856 0 _068_
rlabel metal3 27272 15120 27272 15120 0 _069_
rlabel metal2 18088 23744 18088 23744 0 _070_
rlabel metal2 22456 20160 22456 20160 0 _071_
rlabel metal2 18648 18928 18648 18928 0 _072_
rlabel metal2 19544 19600 19544 19600 0 _073_
rlabel metal3 19544 16632 19544 16632 0 _074_
rlabel metal3 19712 27048 19712 27048 0 _075_
rlabel metal2 18424 19880 18424 19880 0 _076_
rlabel metal2 21672 18088 21672 18088 0 _077_
rlabel metal3 20104 16072 20104 16072 0 _078_
rlabel metal2 22624 23352 22624 23352 0 _079_
rlabel metal2 21448 16128 21448 16128 0 _080_
rlabel metal2 20552 15624 20552 15624 0 _081_
rlabel metal2 21560 19768 21560 19768 0 _082_
rlabel metal2 19320 20944 19320 20944 0 _083_
rlabel metal2 26264 19768 26264 19768 0 _084_
rlabel metal3 29344 20552 29344 20552 0 _085_
rlabel metal3 22232 27104 22232 27104 0 _086_
rlabel metal2 15064 19264 15064 19264 0 _087_
rlabel metal2 14168 24584 14168 24584 0 _088_
rlabel metal2 14056 25424 14056 25424 0 _089_
rlabel metal2 14280 26264 14280 26264 0 _090_
rlabel metal2 13496 22624 13496 22624 0 _091_
rlabel metal2 18424 22344 18424 22344 0 _092_
rlabel metal2 17472 24696 17472 24696 0 _093_
rlabel metal2 13832 23016 13832 23016 0 _094_
rlabel metal2 14056 22176 14056 22176 0 _095_
rlabel metal2 17416 22512 17416 22512 0 _096_
rlabel metal2 19040 27832 19040 27832 0 _097_
rlabel metal2 19880 27888 19880 27888 0 _098_
rlabel metal3 2478 27608 2478 27608 0 clk
rlabel metal2 23352 21112 23352 21112 0 clknet_0_clk
rlabel metal2 21280 28392 21280 28392 0 clknet_1_0__leaf_clk
rlabel metal3 22680 27832 22680 27832 0 clknet_1_1__leaf_clk
rlabel metal2 20216 27104 20216 27104 0 dut9.count\[0\]
rlabel metal2 17640 22960 17640 22960 0 dut9.count\[1\]
rlabel metal2 14504 21896 14504 21896 0 dut9.count\[2\]
rlabel metal2 23016 22736 23016 22736 0 dut9.count\[3\]
rlabel metal3 29484 23688 29484 23688 0 net1
rlabel metal2 24584 5964 24584 5964 0 net10
rlabel metal2 17752 6748 17752 6748 0 net11
rlabel metal2 10024 20776 10024 20776 0 net12
rlabel metal2 11816 26208 11816 26208 0 net13
rlabel metal3 6356 19208 6356 19208 0 net14
rlabel metal2 28616 16464 28616 16464 0 net15
rlabel metal2 19264 27608 19264 27608 0 net16
rlabel metal2 24136 29988 24136 29988 0 net17
rlabel metal2 20216 28392 20216 28392 0 net18
rlabel metal2 30184 20776 30184 20776 0 net19
rlabel metal3 27552 21448 27552 21448 0 net2
rlabel metal2 22232 13552 22232 13552 0 net20
rlabel metal2 37688 19656 37688 19656 0 net21
rlabel metal2 29288 22624 29288 22624 0 net22
rlabel metal3 6356 27048 6356 27048 0 net23
rlabel metal2 4312 18368 4312 18368 0 net24
rlabel metal2 24248 2590 24248 2590 0 net25
rlabel metal2 40264 26712 40264 26712 0 net26
rlabel metal2 31416 21056 31416 21056 0 net3
rlabel metal2 25816 6356 25816 6356 0 net4
rlabel metal2 19096 9716 19096 9716 0 net5
rlabel metal2 23464 27888 23464 27888 0 net6
rlabel metal2 37912 24136 37912 24136 0 net7
rlabel metal2 19712 3528 19712 3528 0 net8
rlabel metal2 30184 17136 30184 17136 0 net9
rlabel metal2 40040 23800 40040 23800 0 segm[0]
rlabel metal2 40040 22008 40040 22008 0 segm[10]
rlabel metal2 39928 21168 39928 21168 0 segm[11]
rlabel metal2 25592 2086 25592 2086 0 segm[12]
rlabel metal2 18872 2422 18872 2422 0 segm[1]
rlabel metal2 22232 39690 22232 39690 0 segm[2]
rlabel metal2 40040 24360 40040 24360 0 segm[3]
rlabel metal2 18200 2198 18200 2198 0 segm[4]
rlabel metal2 40040 17640 40040 17640 0 segm[6]
rlabel metal2 23576 2198 23576 2198 0 segm[7]
rlabel metal2 17528 2982 17528 2982 0 segm[8]
rlabel metal3 1358 20888 1358 20888 0 segm[9]
rlabel metal3 1414 26936 1414 26936 0 sel[0]
rlabel metal3 1358 18872 1358 18872 0 sel[10]
rlabel metal2 40040 16408 40040 16408 0 sel[11]
rlabel metal2 18200 39690 18200 39690 0 sel[1]
rlabel metal2 22904 39746 22904 39746 0 sel[2]
rlabel metal2 20888 39354 20888 39354 0 sel[3]
rlabel metal2 40040 20552 40040 20552 0 sel[4]
rlabel metal2 22232 2030 22232 2030 0 sel[5]
rlabel metal2 40040 19656 40040 19656 0 sel[6]
rlabel metal3 40642 22904 40642 22904 0 sel[7]
rlabel metal3 1358 26264 1358 26264 0 sel[8]
rlabel metal3 1358 18200 1358 18200 0 sel[9]
<< properties >>
string FIXED_BBOX 0 0 42000 42000
<< end >>
