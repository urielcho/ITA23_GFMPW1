magic
tech gf180mcuD
magscale 1 10
timestamp 1699641146
<< metal1 >>
rect 1344 38442 40656 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 40656 38442
rect 1344 38356 40656 38390
rect 18622 38274 18674 38286
rect 18622 38210 18674 38222
rect 22094 38274 22146 38286
rect 22094 38210 22146 38222
rect 25566 38274 25618 38286
rect 25566 38210 25618 38222
rect 18050 37998 18062 38050
rect 18114 37998 18126 38050
rect 21298 37998 21310 38050
rect 21362 37998 21374 38050
rect 24546 37998 24558 38050
rect 24610 37998 24622 38050
rect 1344 37658 40656 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 40656 37658
rect 1344 37572 40656 37606
rect 18398 37490 18450 37502
rect 18398 37426 18450 37438
rect 28142 37490 28194 37502
rect 28142 37426 28194 37438
rect 17378 37214 17390 37266
rect 17442 37214 17454 37266
rect 27570 37214 27582 37266
rect 27634 37214 27646 37266
rect 1344 36874 40656 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 40656 36874
rect 1344 36788 40656 36822
rect 17390 36706 17442 36718
rect 17390 36642 17442 36654
rect 16370 36430 16382 36482
rect 16434 36430 16446 36482
rect 40238 36370 40290 36382
rect 40238 36306 40290 36318
rect 1344 36090 40656 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 40656 36090
rect 1344 36004 40656 36038
rect 1344 35306 40656 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 40656 35306
rect 1344 35220 40656 35254
rect 1344 34522 40656 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 40656 34522
rect 1344 34436 40656 34470
rect 1344 33738 40656 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 40656 33738
rect 1344 33652 40656 33686
rect 1344 32954 40656 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 40656 32954
rect 1344 32868 40656 32902
rect 1344 32170 40656 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 40656 32170
rect 1344 32084 40656 32118
rect 1344 31386 40656 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 40656 31386
rect 1344 31300 40656 31334
rect 1344 30602 40656 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 40656 30602
rect 1344 30516 40656 30550
rect 1344 29818 40656 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 40656 29818
rect 1344 29732 40656 29766
rect 17614 29314 17666 29326
rect 17614 29250 17666 29262
rect 1344 29034 40656 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 40656 29034
rect 1344 28948 40656 28982
rect 18062 28754 18114 28766
rect 18062 28690 18114 28702
rect 16158 28530 16210 28542
rect 16158 28466 16210 28478
rect 16270 28530 16322 28542
rect 16270 28466 16322 28478
rect 16942 28530 16994 28542
rect 17266 28478 17278 28530
rect 17330 28478 17342 28530
rect 16942 28466 16994 28478
rect 16494 28418 16546 28430
rect 16494 28354 16546 28366
rect 1344 28250 40656 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 40656 28250
rect 1344 28164 40656 28198
rect 17390 27970 17442 27982
rect 17390 27906 17442 27918
rect 17726 27858 17778 27870
rect 13906 27806 13918 27858
rect 13970 27806 13982 27858
rect 17726 27794 17778 27806
rect 17950 27858 18002 27870
rect 18498 27806 18510 27858
rect 18562 27806 18574 27858
rect 25218 27806 25230 27858
rect 25282 27806 25294 27858
rect 17950 27794 18002 27806
rect 17502 27746 17554 27758
rect 28702 27746 28754 27758
rect 14690 27694 14702 27746
rect 14754 27694 14766 27746
rect 16818 27694 16830 27746
rect 16882 27694 16894 27746
rect 19170 27694 19182 27746
rect 19234 27694 19246 27746
rect 21298 27694 21310 27746
rect 21362 27694 21374 27746
rect 26002 27694 26014 27746
rect 26066 27694 26078 27746
rect 28130 27694 28142 27746
rect 28194 27694 28206 27746
rect 17502 27682 17554 27694
rect 28702 27682 28754 27694
rect 1344 27466 40656 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 40656 27466
rect 1344 27380 40656 27414
rect 19630 27298 19682 27310
rect 19630 27234 19682 27246
rect 19070 27186 19122 27198
rect 40014 27186 40066 27198
rect 17154 27134 17166 27186
rect 17218 27134 17230 27186
rect 24210 27134 24222 27186
rect 24274 27134 24286 27186
rect 27682 27134 27694 27186
rect 27746 27134 27758 27186
rect 19070 27122 19122 27134
rect 40014 27122 40066 27134
rect 17390 27074 17442 27086
rect 14354 27022 14366 27074
rect 14418 27022 14430 27074
rect 17390 27010 17442 27022
rect 17950 27074 18002 27086
rect 17950 27010 18002 27022
rect 18286 27074 18338 27086
rect 18286 27010 18338 27022
rect 18622 27074 18674 27086
rect 28142 27074 28194 27086
rect 19618 27022 19630 27074
rect 19682 27022 19694 27074
rect 21410 27022 21422 27074
rect 21474 27022 21486 27074
rect 24770 27022 24782 27074
rect 24834 27022 24846 27074
rect 37650 27022 37662 27074
rect 37714 27022 37726 27074
rect 18622 27010 18674 27022
rect 28142 27010 28194 27022
rect 17614 26962 17666 26974
rect 15026 26910 15038 26962
rect 15090 26910 15102 26962
rect 17614 26898 17666 26910
rect 17838 26962 17890 26974
rect 17838 26898 17890 26910
rect 18510 26962 18562 26974
rect 18510 26898 18562 26910
rect 19966 26962 20018 26974
rect 22082 26910 22094 26962
rect 22146 26910 22158 26962
rect 25554 26910 25566 26962
rect 25618 26910 25630 26962
rect 19966 26898 20018 26910
rect 1344 26682 40656 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 40656 26682
rect 1344 26596 40656 26630
rect 20414 26514 20466 26526
rect 17490 26462 17502 26514
rect 17554 26462 17566 26514
rect 20414 26450 20466 26462
rect 20526 26514 20578 26526
rect 20526 26450 20578 26462
rect 23326 26514 23378 26526
rect 23326 26450 23378 26462
rect 24446 26514 24498 26526
rect 26574 26514 26626 26526
rect 25554 26462 25566 26514
rect 25618 26462 25630 26514
rect 24446 26450 24498 26462
rect 26574 26450 26626 26462
rect 18510 26402 18562 26414
rect 18510 26338 18562 26350
rect 20638 26402 20690 26414
rect 20638 26338 20690 26350
rect 22654 26402 22706 26414
rect 27134 26402 27186 26414
rect 25442 26350 25454 26402
rect 25506 26350 25518 26402
rect 22654 26338 22706 26350
rect 27134 26338 27186 26350
rect 18062 26290 18114 26302
rect 20302 26290 20354 26302
rect 22766 26290 22818 26302
rect 25678 26290 25730 26302
rect 18722 26238 18734 26290
rect 18786 26238 18798 26290
rect 21074 26238 21086 26290
rect 21138 26238 21150 26290
rect 23538 26238 23550 26290
rect 23602 26238 23614 26290
rect 25218 26238 25230 26290
rect 25282 26238 25294 26290
rect 18062 26226 18114 26238
rect 20302 26226 20354 26238
rect 22766 26226 22818 26238
rect 25678 26226 25730 26238
rect 26126 26290 26178 26302
rect 26126 26226 26178 26238
rect 26350 26290 26402 26302
rect 26350 26226 26402 26238
rect 26686 26290 26738 26302
rect 26686 26226 26738 26238
rect 27022 26290 27074 26302
rect 27022 26226 27074 26238
rect 25902 26178 25954 26190
rect 25902 26114 25954 26126
rect 17838 26066 17890 26078
rect 17838 26002 17890 26014
rect 22654 26066 22706 26078
rect 22654 26002 22706 26014
rect 23214 26066 23266 26078
rect 23214 26002 23266 26014
rect 1344 25898 40656 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 40656 25898
rect 1344 25812 40656 25846
rect 23202 25678 23214 25730
rect 23266 25678 23278 25730
rect 25566 25618 25618 25630
rect 25566 25554 25618 25566
rect 40014 25618 40066 25630
rect 40014 25554 40066 25566
rect 22318 25506 22370 25518
rect 25118 25506 25170 25518
rect 21746 25454 21758 25506
rect 21810 25454 21822 25506
rect 22418 25454 22430 25506
rect 22482 25454 22494 25506
rect 23314 25454 23326 25506
rect 23378 25454 23390 25506
rect 23762 25454 23774 25506
rect 23826 25454 23838 25506
rect 22318 25442 22370 25454
rect 25118 25442 25170 25454
rect 25454 25506 25506 25518
rect 25454 25442 25506 25454
rect 25790 25506 25842 25518
rect 37650 25454 37662 25506
rect 37714 25454 37726 25506
rect 25790 25442 25842 25454
rect 21310 25394 21362 25406
rect 21310 25330 21362 25342
rect 29262 25394 29314 25406
rect 29262 25330 29314 25342
rect 29374 25394 29426 25406
rect 29374 25330 29426 25342
rect 29038 25282 29090 25294
rect 29038 25218 29090 25230
rect 1344 25114 40656 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 40656 25114
rect 1344 25028 40656 25062
rect 16382 24946 16434 24958
rect 16382 24882 16434 24894
rect 17278 24946 17330 24958
rect 17278 24882 17330 24894
rect 17502 24946 17554 24958
rect 17502 24882 17554 24894
rect 19854 24946 19906 24958
rect 27358 24946 27410 24958
rect 23202 24894 23214 24946
rect 23266 24894 23278 24946
rect 19854 24882 19906 24894
rect 27358 24882 27410 24894
rect 17614 24722 17666 24734
rect 4274 24670 4286 24722
rect 4338 24670 4350 24722
rect 15922 24670 15934 24722
rect 15986 24670 15998 24722
rect 17614 24658 17666 24670
rect 19742 24722 19794 24734
rect 20974 24722 21026 24734
rect 22878 24722 22930 24734
rect 20738 24670 20750 24722
rect 20802 24670 20814 24722
rect 21634 24670 21646 24722
rect 21698 24670 21710 24722
rect 27682 24670 27694 24722
rect 27746 24670 27758 24722
rect 19742 24658 19794 24670
rect 20974 24658 21026 24670
rect 22878 24658 22930 24670
rect 22654 24610 22706 24622
rect 13010 24558 13022 24610
rect 13074 24558 13086 24610
rect 15138 24558 15150 24610
rect 15202 24558 15214 24610
rect 20850 24558 20862 24610
rect 20914 24558 20926 24610
rect 21298 24558 21310 24610
rect 21362 24558 21374 24610
rect 28466 24558 28478 24610
rect 28530 24558 28542 24610
rect 30594 24558 30606 24610
rect 30658 24558 30670 24610
rect 22654 24546 22706 24558
rect 1934 24498 1986 24510
rect 1934 24434 1986 24446
rect 19854 24498 19906 24510
rect 19854 24434 19906 24446
rect 1344 24330 40656 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 40656 24330
rect 1344 24244 40656 24278
rect 14814 24162 14866 24174
rect 14814 24098 14866 24110
rect 16158 24162 16210 24174
rect 16158 24098 16210 24110
rect 23214 24162 23266 24174
rect 23214 24098 23266 24110
rect 1934 24050 1986 24062
rect 15262 24050 15314 24062
rect 9986 23998 9998 24050
rect 10050 23998 10062 24050
rect 1934 23986 1986 23998
rect 15262 23986 15314 23998
rect 15822 24050 15874 24062
rect 29262 24050 29314 24062
rect 16930 23998 16942 24050
rect 16994 23998 17006 24050
rect 15822 23986 15874 23998
rect 29262 23986 29314 23998
rect 13806 23938 13858 23950
rect 4274 23886 4286 23938
rect 4338 23886 4350 23938
rect 12898 23886 12910 23938
rect 12962 23886 12974 23938
rect 13806 23874 13858 23886
rect 13918 23938 13970 23950
rect 13918 23874 13970 23886
rect 14926 23938 14978 23950
rect 14926 23874 14978 23886
rect 15150 23938 15202 23950
rect 17614 23938 17666 23950
rect 21870 23938 21922 23950
rect 22878 23938 22930 23950
rect 16482 23886 16494 23938
rect 16546 23886 16558 23938
rect 17938 23886 17950 23938
rect 18002 23886 18014 23938
rect 18162 23886 18174 23938
rect 18226 23886 18238 23938
rect 22418 23886 22430 23938
rect 22482 23886 22494 23938
rect 15150 23874 15202 23886
rect 17614 23874 17666 23886
rect 21870 23874 21922 23886
rect 22878 23874 22930 23886
rect 29038 23938 29090 23950
rect 29038 23874 29090 23886
rect 29486 23938 29538 23950
rect 29486 23874 29538 23886
rect 29598 23938 29650 23950
rect 29598 23874 29650 23886
rect 13470 23826 13522 23838
rect 12114 23774 12126 23826
rect 12178 23774 12190 23826
rect 13470 23762 13522 23774
rect 13582 23826 13634 23838
rect 13582 23762 13634 23774
rect 15710 23826 15762 23838
rect 19406 23826 19458 23838
rect 23102 23826 23154 23838
rect 15922 23774 15934 23826
rect 15986 23774 15998 23826
rect 20290 23774 20302 23826
rect 20354 23774 20366 23826
rect 21970 23774 21982 23826
rect 22034 23774 22046 23826
rect 22306 23774 22318 23826
rect 22370 23774 22382 23826
rect 15710 23762 15762 23774
rect 19406 23762 19458 23774
rect 23102 23762 23154 23774
rect 23214 23826 23266 23838
rect 23214 23762 23266 23774
rect 17390 23714 17442 23726
rect 17390 23650 17442 23662
rect 17726 23714 17778 23726
rect 17726 23650 17778 23662
rect 19294 23714 19346 23726
rect 19294 23650 19346 23662
rect 20638 23714 20690 23726
rect 20638 23650 20690 23662
rect 1344 23546 40656 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 40656 23546
rect 1344 23460 40656 23494
rect 12798 23378 12850 23390
rect 12798 23314 12850 23326
rect 13022 23378 13074 23390
rect 13022 23314 13074 23326
rect 13358 23378 13410 23390
rect 13358 23314 13410 23326
rect 15934 23378 15986 23390
rect 22542 23378 22594 23390
rect 18722 23326 18734 23378
rect 18786 23326 18798 23378
rect 15934 23314 15986 23326
rect 22542 23314 22594 23326
rect 24222 23378 24274 23390
rect 24222 23314 24274 23326
rect 25230 23378 25282 23390
rect 25230 23314 25282 23326
rect 26126 23378 26178 23390
rect 26126 23314 26178 23326
rect 28478 23378 28530 23390
rect 28478 23314 28530 23326
rect 15822 23266 15874 23278
rect 15822 23202 15874 23214
rect 16046 23266 16098 23278
rect 19406 23266 19458 23278
rect 18274 23214 18286 23266
rect 18338 23214 18350 23266
rect 18498 23214 18510 23266
rect 18562 23214 18574 23266
rect 16046 23202 16098 23214
rect 19406 23202 19458 23214
rect 19854 23266 19906 23278
rect 23102 23266 23154 23278
rect 20738 23214 20750 23266
rect 20802 23214 20814 23266
rect 21634 23214 21646 23266
rect 21698 23214 21710 23266
rect 21970 23214 21982 23266
rect 22034 23214 22046 23266
rect 19854 23202 19906 23214
rect 23102 23202 23154 23214
rect 23214 23266 23266 23278
rect 23998 23266 24050 23278
rect 23314 23214 23326 23266
rect 23378 23214 23390 23266
rect 23214 23202 23266 23214
rect 23998 23202 24050 23214
rect 26910 23266 26962 23278
rect 26910 23202 26962 23214
rect 12686 23154 12738 23166
rect 20414 23154 20466 23166
rect 22878 23154 22930 23166
rect 18050 23102 18062 23154
rect 18114 23102 18126 23154
rect 19618 23102 19630 23154
rect 19682 23102 19694 23154
rect 22194 23102 22206 23154
rect 22258 23102 22270 23154
rect 12686 23090 12738 23102
rect 20414 23090 20466 23102
rect 22878 23090 22930 23102
rect 22990 23154 23042 23166
rect 26574 23154 26626 23166
rect 25442 23102 25454 23154
rect 25506 23102 25518 23154
rect 22990 23090 23042 23102
rect 26574 23090 26626 23102
rect 28142 23154 28194 23166
rect 28142 23090 28194 23102
rect 28590 23154 28642 23166
rect 28590 23090 28642 23102
rect 28702 23154 28754 23166
rect 37650 23102 37662 23154
rect 37714 23102 37726 23154
rect 28702 23090 28754 23102
rect 19294 23042 19346 23054
rect 19294 22978 19346 22990
rect 21534 23042 21586 23054
rect 26014 23042 26066 23054
rect 24322 22990 24334 23042
rect 24386 22990 24398 23042
rect 21534 22978 21586 22990
rect 26014 22978 26066 22990
rect 25902 22930 25954 22942
rect 25902 22866 25954 22878
rect 40014 22930 40066 22942
rect 40014 22866 40066 22878
rect 1344 22762 40656 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 40656 22762
rect 1344 22676 40656 22710
rect 16718 22594 16770 22606
rect 29934 22594 29986 22606
rect 28354 22542 28366 22594
rect 28418 22591 28430 22594
rect 28690 22591 28702 22594
rect 28418 22545 28702 22591
rect 28418 22542 28430 22545
rect 28690 22542 28702 22545
rect 28754 22542 28766 22594
rect 16718 22530 16770 22542
rect 29934 22530 29986 22542
rect 18622 22482 18674 22494
rect 22206 22482 22258 22494
rect 28590 22482 28642 22494
rect 20738 22430 20750 22482
rect 20802 22430 20814 22482
rect 24210 22430 24222 22482
rect 24274 22430 24286 22482
rect 26002 22430 26014 22482
rect 26066 22430 26078 22482
rect 28130 22430 28142 22482
rect 28194 22430 28206 22482
rect 18622 22418 18674 22430
rect 22206 22418 22258 22430
rect 28590 22418 28642 22430
rect 40014 22482 40066 22494
rect 40014 22418 40066 22430
rect 17838 22370 17890 22382
rect 19742 22370 19794 22382
rect 21870 22370 21922 22382
rect 17266 22318 17278 22370
rect 17330 22318 17342 22370
rect 19282 22318 19294 22370
rect 19346 22318 19358 22370
rect 20626 22318 20638 22370
rect 20690 22318 20702 22370
rect 22530 22318 22542 22370
rect 22594 22318 22606 22370
rect 22978 22318 22990 22370
rect 23042 22318 23054 22370
rect 23538 22318 23550 22370
rect 23602 22318 23614 22370
rect 24658 22318 24670 22370
rect 24722 22318 24734 22370
rect 25330 22318 25342 22370
rect 25394 22318 25406 22370
rect 29362 22318 29374 22370
rect 29426 22318 29438 22370
rect 37650 22318 37662 22370
rect 37714 22318 37726 22370
rect 17838 22306 17890 22318
rect 19742 22306 19794 22318
rect 21870 22306 21922 22318
rect 13582 22258 13634 22270
rect 13582 22194 13634 22206
rect 13694 22258 13746 22270
rect 13694 22194 13746 22206
rect 13918 22258 13970 22270
rect 13918 22194 13970 22206
rect 14142 22258 14194 22270
rect 14142 22194 14194 22206
rect 14254 22258 14306 22270
rect 14254 22194 14306 22206
rect 16830 22258 16882 22270
rect 18510 22258 18562 22270
rect 18162 22206 18174 22258
rect 18226 22206 18238 22258
rect 16830 22194 16882 22206
rect 18510 22194 18562 22206
rect 18734 22258 18786 22270
rect 21422 22258 21474 22270
rect 20290 22206 20302 22258
rect 20354 22206 20366 22258
rect 18734 22194 18786 22206
rect 21422 22194 21474 22206
rect 22094 22258 22146 22270
rect 29822 22258 29874 22270
rect 22642 22206 22654 22258
rect 22706 22206 22718 22258
rect 24546 22206 24558 22258
rect 24610 22206 24622 22258
rect 22094 22194 22146 22206
rect 29822 22194 29874 22206
rect 29934 22258 29986 22270
rect 29934 22194 29986 22206
rect 13358 22146 13410 22158
rect 13358 22082 13410 22094
rect 16718 22146 16770 22158
rect 16718 22082 16770 22094
rect 17502 22146 17554 22158
rect 17502 22082 17554 22094
rect 21646 22146 21698 22158
rect 29138 22094 29150 22146
rect 29202 22094 29214 22146
rect 21646 22082 21698 22094
rect 1344 21978 40656 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 40656 21978
rect 1344 21892 40656 21926
rect 11566 21810 11618 21822
rect 11566 21746 11618 21758
rect 15374 21810 15426 21822
rect 15374 21746 15426 21758
rect 17502 21810 17554 21822
rect 17502 21746 17554 21758
rect 17838 21810 17890 21822
rect 17838 21746 17890 21758
rect 25566 21810 25618 21822
rect 25566 21746 25618 21758
rect 25678 21810 25730 21822
rect 27582 21810 27634 21822
rect 26226 21758 26238 21810
rect 26290 21758 26302 21810
rect 25678 21746 25730 21758
rect 27582 21746 27634 21758
rect 26574 21698 26626 21710
rect 12786 21646 12798 21698
rect 12850 21646 12862 21698
rect 19618 21646 19630 21698
rect 19682 21646 19694 21698
rect 20850 21646 20862 21698
rect 20914 21646 20926 21698
rect 23762 21646 23774 21698
rect 23826 21646 23838 21698
rect 28690 21646 28702 21698
rect 28754 21646 28766 21698
rect 26574 21634 26626 21646
rect 11454 21586 11506 21598
rect 4274 21534 4286 21586
rect 4338 21534 4350 21586
rect 11454 21522 11506 21534
rect 11790 21586 11842 21598
rect 16270 21586 16322 21598
rect 25454 21586 25506 21598
rect 12114 21534 12126 21586
rect 12178 21534 12190 21586
rect 20402 21534 20414 21586
rect 20466 21534 20478 21586
rect 20738 21534 20750 21586
rect 20802 21534 20814 21586
rect 22642 21534 22654 21586
rect 22706 21534 22718 21586
rect 23202 21534 23214 21586
rect 23266 21534 23278 21586
rect 25218 21534 25230 21586
rect 25282 21534 25294 21586
rect 11790 21522 11842 21534
rect 16270 21522 16322 21534
rect 25454 21522 25506 21534
rect 25790 21586 25842 21598
rect 27906 21534 27918 21586
rect 27970 21534 27982 21586
rect 25790 21522 25842 21534
rect 17390 21474 17442 21486
rect 14914 21422 14926 21474
rect 14978 21422 14990 21474
rect 16706 21422 16718 21474
rect 16770 21422 16782 21474
rect 17390 21410 17442 21422
rect 18398 21474 18450 21486
rect 21522 21422 21534 21474
rect 21586 21422 21598 21474
rect 23426 21422 23438 21474
rect 23490 21422 23502 21474
rect 30818 21422 30830 21474
rect 30882 21422 30894 21474
rect 18398 21410 18450 21422
rect 1934 21362 1986 21374
rect 1934 21298 1986 21310
rect 1344 21194 40656 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 40656 21194
rect 1344 21108 40656 21142
rect 14814 20914 14866 20926
rect 40014 20914 40066 20926
rect 9874 20862 9886 20914
rect 9938 20862 9950 20914
rect 12002 20862 12014 20914
rect 12066 20862 12078 20914
rect 13458 20862 13470 20914
rect 13522 20862 13534 20914
rect 16146 20862 16158 20914
rect 16210 20862 16222 20914
rect 27906 20862 27918 20914
rect 27970 20862 27982 20914
rect 14814 20850 14866 20862
rect 40014 20850 40066 20862
rect 14030 20802 14082 20814
rect 12786 20750 12798 20802
rect 12850 20750 12862 20802
rect 13682 20750 13694 20802
rect 13746 20750 13758 20802
rect 14030 20738 14082 20750
rect 14478 20802 14530 20814
rect 29374 20802 29426 20814
rect 20066 20750 20078 20802
rect 20130 20750 20142 20802
rect 21298 20750 21310 20802
rect 21362 20750 21374 20802
rect 22194 20750 22206 20802
rect 22258 20750 22270 20802
rect 22530 20750 22542 20802
rect 22594 20750 22606 20802
rect 23538 20750 23550 20802
rect 23602 20750 23614 20802
rect 37650 20750 37662 20802
rect 37714 20750 37726 20802
rect 14478 20738 14530 20750
rect 29374 20738 29426 20750
rect 13470 20690 13522 20702
rect 21410 20638 21422 20690
rect 21474 20638 21486 20690
rect 22754 20638 22766 20690
rect 22818 20638 22830 20690
rect 13470 20626 13522 20638
rect 29038 20578 29090 20590
rect 29038 20514 29090 20526
rect 29262 20578 29314 20590
rect 29262 20514 29314 20526
rect 1344 20410 40656 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 40656 20410
rect 1344 20324 40656 20358
rect 13906 20190 13918 20242
rect 13970 20190 13982 20242
rect 12574 20130 12626 20142
rect 12574 20066 12626 20078
rect 12686 20130 12738 20142
rect 12686 20066 12738 20078
rect 13582 20130 13634 20142
rect 13582 20066 13634 20078
rect 15598 20130 15650 20142
rect 17502 20130 17554 20142
rect 18174 20130 18226 20142
rect 25454 20130 25506 20142
rect 16818 20078 16830 20130
rect 16882 20078 16894 20130
rect 17826 20078 17838 20130
rect 17890 20078 17902 20130
rect 21858 20078 21870 20130
rect 21922 20078 21934 20130
rect 15598 20066 15650 20078
rect 17502 20066 17554 20078
rect 18174 20066 18226 20078
rect 25454 20066 25506 20078
rect 26686 20130 26738 20142
rect 26686 20066 26738 20078
rect 12910 20018 12962 20030
rect 4274 19966 4286 20018
rect 4338 19966 4350 20018
rect 12910 19954 12962 19966
rect 13358 20018 13410 20030
rect 13358 19954 13410 19966
rect 14254 20018 14306 20030
rect 19070 20018 19122 20030
rect 25230 20018 25282 20030
rect 26238 20018 26290 20030
rect 16594 19966 16606 20018
rect 16658 19966 16670 20018
rect 19394 19966 19406 20018
rect 19458 19966 19470 20018
rect 25666 19966 25678 20018
rect 25730 19966 25742 20018
rect 25890 19966 25902 20018
rect 25954 19966 25966 20018
rect 14254 19954 14306 19966
rect 19070 19954 19122 19966
rect 25230 19954 25282 19966
rect 26238 19954 26290 19966
rect 26910 20018 26962 20030
rect 27906 19966 27918 20018
rect 27970 19966 27982 20018
rect 37650 19966 37662 20018
rect 37714 19966 37726 20018
rect 26910 19954 26962 19966
rect 13134 19906 13186 19918
rect 18510 19906 18562 19918
rect 26462 19906 26514 19918
rect 16706 19854 16718 19906
rect 16770 19854 16782 19906
rect 26002 19854 26014 19906
rect 26066 19854 26078 19906
rect 13134 19842 13186 19854
rect 18510 19842 18562 19854
rect 26462 19842 26514 19854
rect 27582 19906 27634 19918
rect 28690 19854 28702 19906
rect 28754 19854 28766 19906
rect 30818 19854 30830 19906
rect 30882 19854 30894 19906
rect 27582 19842 27634 19854
rect 1934 19794 1986 19806
rect 1934 19730 1986 19742
rect 12574 19794 12626 19806
rect 12574 19730 12626 19742
rect 15486 19794 15538 19806
rect 15486 19730 15538 19742
rect 15822 19794 15874 19806
rect 15822 19730 15874 19742
rect 40014 19794 40066 19806
rect 40014 19730 40066 19742
rect 1344 19626 40656 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 40656 19626
rect 1344 19540 40656 19574
rect 22866 19406 22878 19458
rect 22930 19406 22942 19458
rect 1934 19346 1986 19358
rect 13582 19346 13634 19358
rect 9874 19294 9886 19346
rect 9938 19294 9950 19346
rect 12002 19294 12014 19346
rect 12066 19294 12078 19346
rect 1934 19282 1986 19294
rect 13582 19282 13634 19294
rect 15598 19346 15650 19358
rect 15598 19282 15650 19294
rect 16382 19346 16434 19358
rect 16382 19282 16434 19294
rect 21758 19346 21810 19358
rect 22754 19294 22766 19346
rect 22818 19294 22830 19346
rect 26450 19294 26462 19346
rect 26514 19294 26526 19346
rect 28578 19294 28590 19346
rect 28642 19294 28654 19346
rect 21758 19282 21810 19294
rect 15374 19234 15426 19246
rect 4274 19182 4286 19234
rect 4338 19182 4350 19234
rect 12786 19182 12798 19234
rect 12850 19182 12862 19234
rect 15374 19170 15426 19182
rect 15486 19234 15538 19246
rect 17502 19234 17554 19246
rect 18958 19234 19010 19246
rect 16930 19182 16942 19234
rect 16994 19182 17006 19234
rect 17826 19182 17838 19234
rect 17890 19182 17902 19234
rect 15486 19170 15538 19182
rect 17502 19170 17554 19182
rect 18958 19170 19010 19182
rect 19518 19234 19570 19246
rect 19518 19170 19570 19182
rect 20750 19234 20802 19246
rect 20750 19170 20802 19182
rect 21310 19234 21362 19246
rect 21310 19170 21362 19182
rect 23886 19234 23938 19246
rect 23886 19170 23938 19182
rect 24446 19234 24498 19246
rect 29038 19234 29090 19246
rect 25778 19182 25790 19234
rect 25842 19182 25854 19234
rect 24446 19170 24498 19182
rect 29038 19170 29090 19182
rect 29374 19234 29426 19246
rect 29374 19170 29426 19182
rect 29598 19234 29650 19246
rect 29598 19170 29650 19182
rect 16270 19122 16322 19134
rect 14578 19070 14590 19122
rect 14642 19070 14654 19122
rect 16270 19058 16322 19070
rect 19294 19122 19346 19134
rect 19294 19058 19346 19070
rect 19854 19122 19906 19134
rect 19854 19058 19906 19070
rect 23214 19122 23266 19134
rect 23214 19058 23266 19070
rect 14926 19010 14978 19022
rect 14926 18946 14978 18958
rect 15710 19010 15762 19022
rect 15710 18946 15762 18958
rect 15822 19010 15874 19022
rect 17614 19010 17666 19022
rect 24334 19010 24386 19022
rect 17154 18958 17166 19010
rect 17218 18958 17230 19010
rect 18610 18958 18622 19010
rect 18674 18958 18686 19010
rect 20402 18958 20414 19010
rect 20466 18958 20478 19010
rect 15822 18946 15874 18958
rect 17614 18946 17666 18958
rect 24334 18946 24386 18958
rect 24558 19010 24610 19022
rect 24558 18946 24610 18958
rect 25006 19010 25058 19022
rect 25006 18946 25058 18958
rect 29262 19010 29314 19022
rect 29262 18946 29314 18958
rect 1344 18842 40656 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 40656 18842
rect 1344 18756 40656 18790
rect 19630 18674 19682 18686
rect 22878 18674 22930 18686
rect 12338 18622 12350 18674
rect 12402 18622 12414 18674
rect 22306 18622 22318 18674
rect 22370 18622 22382 18674
rect 19630 18610 19682 18622
rect 22878 18610 22930 18622
rect 23326 18674 23378 18686
rect 23650 18622 23662 18674
rect 23714 18622 23726 18674
rect 23326 18610 23378 18622
rect 17838 18562 17890 18574
rect 17838 18498 17890 18510
rect 18734 18562 18786 18574
rect 18734 18498 18786 18510
rect 18846 18562 18898 18574
rect 18846 18498 18898 18510
rect 20526 18562 20578 18574
rect 20526 18498 20578 18510
rect 22766 18562 22818 18574
rect 22766 18498 22818 18510
rect 23998 18562 24050 18574
rect 23998 18498 24050 18510
rect 18622 18450 18674 18462
rect 12562 18398 12574 18450
rect 12626 18398 12638 18450
rect 13570 18398 13582 18450
rect 13634 18398 13646 18450
rect 14354 18398 14366 18450
rect 14418 18398 14430 18450
rect 18622 18386 18674 18398
rect 21422 18450 21474 18462
rect 21422 18386 21474 18398
rect 21534 18450 21586 18462
rect 21534 18386 21586 18398
rect 21982 18450 22034 18462
rect 21982 18386 22034 18398
rect 24110 18450 24162 18462
rect 24110 18386 24162 18398
rect 24222 18450 24274 18462
rect 24222 18386 24274 18398
rect 24670 18450 24722 18462
rect 24670 18386 24722 18398
rect 18062 18338 18114 18350
rect 16482 18286 16494 18338
rect 16546 18286 16558 18338
rect 17714 18286 17726 18338
rect 17778 18286 17790 18338
rect 18062 18274 18114 18286
rect 20190 18338 20242 18350
rect 20190 18274 20242 18286
rect 22654 18338 22706 18350
rect 22654 18274 22706 18286
rect 28814 18338 28866 18350
rect 28814 18274 28866 18286
rect 20750 18226 20802 18238
rect 19282 18174 19294 18226
rect 19346 18174 19358 18226
rect 20750 18162 20802 18174
rect 21086 18226 21138 18238
rect 21086 18162 21138 18174
rect 1344 18058 40656 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 40656 18058
rect 1344 17972 40656 18006
rect 17390 17890 17442 17902
rect 17390 17826 17442 17838
rect 17726 17890 17778 17902
rect 17726 17826 17778 17838
rect 17614 17778 17666 17790
rect 40014 17778 40066 17790
rect 18610 17726 18622 17778
rect 18674 17726 18686 17778
rect 19506 17726 19518 17778
rect 19570 17726 19582 17778
rect 22642 17726 22654 17778
rect 22706 17726 22718 17778
rect 17614 17714 17666 17726
rect 40014 17714 40066 17726
rect 21198 17666 21250 17678
rect 20514 17614 20526 17666
rect 20578 17614 20590 17666
rect 21198 17602 21250 17614
rect 21646 17666 21698 17678
rect 23886 17666 23938 17678
rect 22530 17614 22542 17666
rect 22594 17614 22606 17666
rect 23426 17614 23438 17666
rect 23490 17614 23502 17666
rect 24210 17614 24222 17666
rect 24274 17614 24286 17666
rect 37650 17614 37662 17666
rect 37714 17614 37726 17666
rect 21646 17602 21698 17614
rect 23886 17602 23938 17614
rect 17278 17554 17330 17566
rect 21870 17554 21922 17566
rect 24446 17554 24498 17566
rect 20738 17502 20750 17554
rect 20802 17502 20814 17554
rect 22866 17502 22878 17554
rect 22930 17502 22942 17554
rect 17278 17490 17330 17502
rect 21870 17490 21922 17502
rect 24446 17490 24498 17502
rect 16718 17442 16770 17454
rect 16718 17378 16770 17390
rect 18174 17442 18226 17454
rect 18174 17378 18226 17390
rect 19070 17442 19122 17454
rect 19070 17378 19122 17390
rect 21758 17442 21810 17454
rect 21758 17378 21810 17390
rect 24558 17442 24610 17454
rect 24558 17378 24610 17390
rect 1344 17274 40656 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 40656 17274
rect 1344 17188 40656 17222
rect 21534 17106 21586 17118
rect 22542 17106 22594 17118
rect 19730 17054 19742 17106
rect 19794 17054 19806 17106
rect 21858 17054 21870 17106
rect 21922 17054 21934 17106
rect 21534 17042 21586 17054
rect 22542 17042 22594 17054
rect 24334 17106 24386 17118
rect 24334 17042 24386 17054
rect 22206 16994 22258 17006
rect 13794 16942 13806 16994
rect 13858 16942 13870 16994
rect 22206 16930 22258 16942
rect 24222 16994 24274 17006
rect 24222 16930 24274 16942
rect 26686 16994 26738 17006
rect 26686 16930 26738 16942
rect 16382 16882 16434 16894
rect 24558 16882 24610 16894
rect 13122 16830 13134 16882
rect 13186 16830 13198 16882
rect 19954 16830 19966 16882
rect 20018 16830 20030 16882
rect 16382 16818 16434 16830
rect 24558 16818 24610 16830
rect 25118 16882 25170 16894
rect 25118 16818 25170 16830
rect 25342 16882 25394 16894
rect 25342 16818 25394 16830
rect 25454 16882 25506 16894
rect 25454 16818 25506 16830
rect 25678 16882 25730 16894
rect 25678 16818 25730 16830
rect 26238 16882 26290 16894
rect 26238 16818 26290 16830
rect 26462 16882 26514 16894
rect 37874 16830 37886 16882
rect 37938 16830 37950 16882
rect 26462 16818 26514 16830
rect 26574 16770 26626 16782
rect 15922 16718 15934 16770
rect 15986 16718 15998 16770
rect 26574 16706 26626 16718
rect 40014 16658 40066 16670
rect 40014 16594 40066 16606
rect 1344 16490 40656 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 40656 16490
rect 1344 16404 40656 16438
rect 27470 16322 27522 16334
rect 27470 16258 27522 16270
rect 24882 16158 24894 16210
rect 24946 16158 24958 16210
rect 27010 16158 27022 16210
rect 27074 16158 27086 16210
rect 21310 16098 21362 16110
rect 24210 16046 24222 16098
rect 24274 16046 24286 16098
rect 21310 16034 21362 16046
rect 27358 15986 27410 15998
rect 27358 15922 27410 15934
rect 27470 15874 27522 15886
rect 21634 15822 21646 15874
rect 21698 15822 21710 15874
rect 27470 15810 27522 15822
rect 28030 15874 28082 15886
rect 28030 15810 28082 15822
rect 1344 15706 40656 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 40656 15706
rect 1344 15620 40656 15654
rect 21310 15538 21362 15550
rect 21310 15474 21362 15486
rect 21534 15538 21586 15550
rect 21534 15474 21586 15486
rect 22318 15538 22370 15550
rect 22318 15474 22370 15486
rect 22542 15538 22594 15550
rect 22542 15474 22594 15486
rect 25454 15538 25506 15550
rect 25454 15474 25506 15486
rect 29486 15538 29538 15550
rect 29486 15474 29538 15486
rect 26898 15374 26910 15426
rect 26962 15374 26974 15426
rect 25230 15314 25282 15326
rect 21746 15262 21758 15314
rect 21810 15262 21822 15314
rect 22082 15262 22094 15314
rect 22146 15262 22158 15314
rect 25230 15250 25282 15262
rect 25566 15314 25618 15326
rect 25566 15250 25618 15262
rect 25790 15314 25842 15326
rect 26114 15262 26126 15314
rect 26178 15262 26190 15314
rect 37650 15262 37662 15314
rect 37714 15262 37726 15314
rect 25790 15250 25842 15262
rect 18398 15202 18450 15214
rect 40014 15202 40066 15214
rect 29026 15150 29038 15202
rect 29090 15150 29102 15202
rect 18398 15138 18450 15150
rect 40014 15138 40066 15150
rect 21646 15090 21698 15102
rect 21646 15026 21698 15038
rect 22654 15090 22706 15102
rect 22654 15026 22706 15038
rect 1344 14922 40656 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 40656 14922
rect 1344 14836 40656 14870
rect 18958 14754 19010 14766
rect 18958 14690 19010 14702
rect 29262 14642 29314 14654
rect 16034 14590 16046 14642
rect 16098 14590 16110 14642
rect 18162 14590 18174 14642
rect 18226 14590 18238 14642
rect 26114 14590 26126 14642
rect 26178 14590 26190 14642
rect 28242 14590 28254 14642
rect 28306 14590 28318 14642
rect 29262 14578 29314 14590
rect 18510 14530 18562 14542
rect 20414 14530 20466 14542
rect 15362 14478 15374 14530
rect 15426 14478 15438 14530
rect 19282 14478 19294 14530
rect 19346 14478 19358 14530
rect 18510 14466 18562 14478
rect 20414 14466 20466 14478
rect 21646 14530 21698 14542
rect 21646 14466 21698 14478
rect 22094 14530 22146 14542
rect 22094 14466 22146 14478
rect 22542 14530 22594 14542
rect 22542 14466 22594 14478
rect 22878 14530 22930 14542
rect 25330 14478 25342 14530
rect 25394 14478 25406 14530
rect 22878 14466 22930 14478
rect 20078 14418 20130 14430
rect 18722 14366 18734 14418
rect 18786 14366 18798 14418
rect 20078 14354 20130 14366
rect 20638 14418 20690 14430
rect 20638 14354 20690 14366
rect 22318 14418 22370 14430
rect 22318 14354 22370 14366
rect 18622 14306 18674 14318
rect 18622 14242 18674 14254
rect 20190 14306 20242 14318
rect 20190 14242 20242 14254
rect 21870 14306 21922 14318
rect 21870 14242 21922 14254
rect 22766 14306 22818 14318
rect 22766 14242 22818 14254
rect 23438 14306 23490 14318
rect 23438 14242 23490 14254
rect 1344 14138 40656 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 40656 14138
rect 1344 14052 40656 14086
rect 17502 13970 17554 13982
rect 17502 13906 17554 13918
rect 18286 13970 18338 13982
rect 18286 13906 18338 13918
rect 18846 13970 18898 13982
rect 18846 13906 18898 13918
rect 19518 13970 19570 13982
rect 19518 13906 19570 13918
rect 20078 13970 20130 13982
rect 20078 13906 20130 13918
rect 26686 13970 26738 13982
rect 26686 13906 26738 13918
rect 26910 13970 26962 13982
rect 26910 13906 26962 13918
rect 19742 13858 19794 13870
rect 14690 13806 14702 13858
rect 14754 13806 14766 13858
rect 19742 13794 19794 13806
rect 19854 13858 19906 13870
rect 25230 13858 25282 13870
rect 21074 13806 21086 13858
rect 21138 13806 21150 13858
rect 19854 13794 19906 13806
rect 25230 13794 25282 13806
rect 27022 13858 27074 13870
rect 27022 13794 27074 13806
rect 23662 13746 23714 13758
rect 14018 13694 14030 13746
rect 14082 13694 14094 13746
rect 20402 13694 20414 13746
rect 20466 13694 20478 13746
rect 23662 13682 23714 13694
rect 23886 13746 23938 13758
rect 25342 13746 25394 13758
rect 24098 13694 24110 13746
rect 24162 13694 24174 13746
rect 25554 13694 25566 13746
rect 25618 13694 25630 13746
rect 23886 13682 23938 13694
rect 25342 13682 25394 13694
rect 18174 13634 18226 13646
rect 16818 13582 16830 13634
rect 16882 13582 16894 13634
rect 17938 13582 17950 13634
rect 18002 13582 18014 13634
rect 23202 13582 23214 13634
rect 23266 13582 23278 13634
rect 17266 13470 17278 13522
rect 17330 13519 17342 13522
rect 17953 13519 17999 13582
rect 18174 13570 18226 13582
rect 17330 13473 17999 13519
rect 23550 13522 23602 13534
rect 17330 13470 17342 13473
rect 23550 13458 23602 13470
rect 1344 13354 40656 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 40656 13354
rect 1344 13268 40656 13302
rect 17614 13074 17666 13086
rect 26126 13074 26178 13086
rect 18610 13022 18622 13074
rect 18674 13022 18686 13074
rect 20738 13022 20750 13074
rect 20802 13022 20814 13074
rect 23426 13022 23438 13074
rect 23490 13022 23502 13074
rect 25554 13022 25566 13074
rect 25618 13022 25630 13074
rect 17614 13010 17666 13022
rect 26126 13010 26178 13022
rect 17826 12910 17838 12962
rect 17890 12910 17902 12962
rect 22642 12910 22654 12962
rect 22706 12910 22718 12962
rect 1344 12570 40656 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 40656 12570
rect 1344 12484 40656 12518
rect 1344 11786 40656 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 40656 11786
rect 1344 11700 40656 11734
rect 1344 11002 40656 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 40656 11002
rect 1344 10916 40656 10950
rect 1344 10218 40656 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 40656 10218
rect 1344 10132 40656 10166
rect 1344 9434 40656 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 40656 9434
rect 1344 9348 40656 9382
rect 40238 9154 40290 9166
rect 40238 9090 40290 9102
rect 1344 8650 40656 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 40656 8650
rect 1344 8564 40656 8598
rect 1344 7866 40656 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 40656 7866
rect 1344 7780 40656 7814
rect 1344 7082 40656 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 40656 7082
rect 1344 6996 40656 7030
rect 1344 6298 40656 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 40656 6298
rect 1344 6212 40656 6246
rect 1344 5514 40656 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 40656 5514
rect 1344 5428 40656 5462
rect 1344 4730 40656 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 40656 4730
rect 1344 4644 40656 4678
rect 25554 4286 25566 4338
rect 25618 4286 25630 4338
rect 26238 4114 26290 4126
rect 26238 4050 26290 4062
rect 1344 3946 40656 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 40656 3946
rect 1344 3860 40656 3894
rect 18622 3666 18674 3678
rect 18622 3602 18674 3614
rect 25566 3666 25618 3678
rect 25566 3602 25618 3614
rect 18050 3502 18062 3554
rect 18114 3502 18126 3554
rect 20738 3502 20750 3554
rect 20802 3502 20814 3554
rect 24546 3502 24558 3554
rect 24610 3502 24622 3554
rect 21758 3330 21810 3342
rect 21758 3266 21810 3278
rect 1344 3162 40656 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 40656 3162
rect 1344 3076 40656 3110
<< via1 >>
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 18622 38222 18674 38274
rect 22094 38222 22146 38274
rect 25566 38222 25618 38274
rect 18062 37998 18114 38050
rect 21310 37998 21362 38050
rect 24558 37998 24610 38050
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 18398 37438 18450 37490
rect 28142 37438 28194 37490
rect 17390 37214 17442 37266
rect 27582 37214 27634 37266
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 17390 36654 17442 36706
rect 16382 36430 16434 36482
rect 40238 36318 40290 36370
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 17614 29262 17666 29314
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 18062 28702 18114 28754
rect 16158 28478 16210 28530
rect 16270 28478 16322 28530
rect 16942 28478 16994 28530
rect 17278 28478 17330 28530
rect 16494 28366 16546 28418
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 17390 27918 17442 27970
rect 13918 27806 13970 27858
rect 17726 27806 17778 27858
rect 17950 27806 18002 27858
rect 18510 27806 18562 27858
rect 25230 27806 25282 27858
rect 14702 27694 14754 27746
rect 16830 27694 16882 27746
rect 17502 27694 17554 27746
rect 19182 27694 19234 27746
rect 21310 27694 21362 27746
rect 26014 27694 26066 27746
rect 28142 27694 28194 27746
rect 28702 27694 28754 27746
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 19630 27246 19682 27298
rect 17166 27134 17218 27186
rect 19070 27134 19122 27186
rect 24222 27134 24274 27186
rect 27694 27134 27746 27186
rect 40014 27134 40066 27186
rect 14366 27022 14418 27074
rect 17390 27022 17442 27074
rect 17950 27022 18002 27074
rect 18286 27022 18338 27074
rect 18622 27022 18674 27074
rect 19630 27022 19682 27074
rect 21422 27022 21474 27074
rect 24782 27022 24834 27074
rect 28142 27022 28194 27074
rect 37662 27022 37714 27074
rect 15038 26910 15090 26962
rect 17614 26910 17666 26962
rect 17838 26910 17890 26962
rect 18510 26910 18562 26962
rect 19966 26910 20018 26962
rect 22094 26910 22146 26962
rect 25566 26910 25618 26962
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 17502 26462 17554 26514
rect 20414 26462 20466 26514
rect 20526 26462 20578 26514
rect 23326 26462 23378 26514
rect 24446 26462 24498 26514
rect 25566 26462 25618 26514
rect 26574 26462 26626 26514
rect 18510 26350 18562 26402
rect 20638 26350 20690 26402
rect 22654 26350 22706 26402
rect 25454 26350 25506 26402
rect 27134 26350 27186 26402
rect 18062 26238 18114 26290
rect 18734 26238 18786 26290
rect 20302 26238 20354 26290
rect 21086 26238 21138 26290
rect 22766 26238 22818 26290
rect 23550 26238 23602 26290
rect 25230 26238 25282 26290
rect 25678 26238 25730 26290
rect 26126 26238 26178 26290
rect 26350 26238 26402 26290
rect 26686 26238 26738 26290
rect 27022 26238 27074 26290
rect 25902 26126 25954 26178
rect 17838 26014 17890 26066
rect 22654 26014 22706 26066
rect 23214 26014 23266 26066
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 23214 25678 23266 25730
rect 25566 25566 25618 25618
rect 40014 25566 40066 25618
rect 21758 25454 21810 25506
rect 22318 25454 22370 25506
rect 22430 25454 22482 25506
rect 23326 25454 23378 25506
rect 23774 25454 23826 25506
rect 25118 25454 25170 25506
rect 25454 25454 25506 25506
rect 25790 25454 25842 25506
rect 37662 25454 37714 25506
rect 21310 25342 21362 25394
rect 29262 25342 29314 25394
rect 29374 25342 29426 25394
rect 29038 25230 29090 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 16382 24894 16434 24946
rect 17278 24894 17330 24946
rect 17502 24894 17554 24946
rect 19854 24894 19906 24946
rect 23214 24894 23266 24946
rect 27358 24894 27410 24946
rect 4286 24670 4338 24722
rect 15934 24670 15986 24722
rect 17614 24670 17666 24722
rect 19742 24670 19794 24722
rect 20750 24670 20802 24722
rect 20974 24670 21026 24722
rect 21646 24670 21698 24722
rect 22878 24670 22930 24722
rect 27694 24670 27746 24722
rect 13022 24558 13074 24610
rect 15150 24558 15202 24610
rect 20862 24558 20914 24610
rect 21310 24558 21362 24610
rect 22654 24558 22706 24610
rect 28478 24558 28530 24610
rect 30606 24558 30658 24610
rect 1934 24446 1986 24498
rect 19854 24446 19906 24498
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 14814 24110 14866 24162
rect 16158 24110 16210 24162
rect 23214 24110 23266 24162
rect 1934 23998 1986 24050
rect 9998 23998 10050 24050
rect 15262 23998 15314 24050
rect 15822 23998 15874 24050
rect 16942 23998 16994 24050
rect 29262 23998 29314 24050
rect 4286 23886 4338 23938
rect 12910 23886 12962 23938
rect 13806 23886 13858 23938
rect 13918 23886 13970 23938
rect 14926 23886 14978 23938
rect 15150 23886 15202 23938
rect 16494 23886 16546 23938
rect 17614 23886 17666 23938
rect 17950 23886 18002 23938
rect 18174 23886 18226 23938
rect 21870 23886 21922 23938
rect 22430 23886 22482 23938
rect 22878 23886 22930 23938
rect 29038 23886 29090 23938
rect 29486 23886 29538 23938
rect 29598 23886 29650 23938
rect 12126 23774 12178 23826
rect 13470 23774 13522 23826
rect 13582 23774 13634 23826
rect 15710 23774 15762 23826
rect 15934 23774 15986 23826
rect 19406 23774 19458 23826
rect 20302 23774 20354 23826
rect 21982 23774 22034 23826
rect 22318 23774 22370 23826
rect 23102 23774 23154 23826
rect 23214 23774 23266 23826
rect 17390 23662 17442 23714
rect 17726 23662 17778 23714
rect 19294 23662 19346 23714
rect 20638 23662 20690 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 12798 23326 12850 23378
rect 13022 23326 13074 23378
rect 13358 23326 13410 23378
rect 15934 23326 15986 23378
rect 18734 23326 18786 23378
rect 22542 23326 22594 23378
rect 24222 23326 24274 23378
rect 25230 23326 25282 23378
rect 26126 23326 26178 23378
rect 28478 23326 28530 23378
rect 15822 23214 15874 23266
rect 16046 23214 16098 23266
rect 18286 23214 18338 23266
rect 18510 23214 18562 23266
rect 19406 23214 19458 23266
rect 19854 23214 19906 23266
rect 20750 23214 20802 23266
rect 21646 23214 21698 23266
rect 21982 23214 22034 23266
rect 23102 23214 23154 23266
rect 23214 23214 23266 23266
rect 23326 23214 23378 23266
rect 23998 23214 24050 23266
rect 26910 23214 26962 23266
rect 12686 23102 12738 23154
rect 18062 23102 18114 23154
rect 19630 23102 19682 23154
rect 20414 23102 20466 23154
rect 22206 23102 22258 23154
rect 22878 23102 22930 23154
rect 22990 23102 23042 23154
rect 25454 23102 25506 23154
rect 26574 23102 26626 23154
rect 28142 23102 28194 23154
rect 28590 23102 28642 23154
rect 28702 23102 28754 23154
rect 37662 23102 37714 23154
rect 19294 22990 19346 23042
rect 21534 22990 21586 23042
rect 24334 22990 24386 23042
rect 26014 22990 26066 23042
rect 25902 22878 25954 22930
rect 40014 22878 40066 22930
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 16718 22542 16770 22594
rect 28366 22542 28418 22594
rect 28702 22542 28754 22594
rect 29934 22542 29986 22594
rect 18622 22430 18674 22482
rect 20750 22430 20802 22482
rect 22206 22430 22258 22482
rect 24222 22430 24274 22482
rect 26014 22430 26066 22482
rect 28142 22430 28194 22482
rect 28590 22430 28642 22482
rect 40014 22430 40066 22482
rect 17278 22318 17330 22370
rect 17838 22318 17890 22370
rect 19294 22318 19346 22370
rect 19742 22318 19794 22370
rect 20638 22318 20690 22370
rect 21870 22318 21922 22370
rect 22542 22318 22594 22370
rect 22990 22318 23042 22370
rect 23550 22318 23602 22370
rect 24670 22318 24722 22370
rect 25342 22318 25394 22370
rect 29374 22318 29426 22370
rect 37662 22318 37714 22370
rect 13582 22206 13634 22258
rect 13694 22206 13746 22258
rect 13918 22206 13970 22258
rect 14142 22206 14194 22258
rect 14254 22206 14306 22258
rect 16830 22206 16882 22258
rect 18174 22206 18226 22258
rect 18510 22206 18562 22258
rect 18734 22206 18786 22258
rect 20302 22206 20354 22258
rect 21422 22206 21474 22258
rect 22094 22206 22146 22258
rect 22654 22206 22706 22258
rect 24558 22206 24610 22258
rect 29822 22206 29874 22258
rect 29934 22206 29986 22258
rect 13358 22094 13410 22146
rect 16718 22094 16770 22146
rect 17502 22094 17554 22146
rect 21646 22094 21698 22146
rect 29150 22094 29202 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 11566 21758 11618 21810
rect 15374 21758 15426 21810
rect 17502 21758 17554 21810
rect 17838 21758 17890 21810
rect 25566 21758 25618 21810
rect 25678 21758 25730 21810
rect 26238 21758 26290 21810
rect 27582 21758 27634 21810
rect 12798 21646 12850 21698
rect 19630 21646 19682 21698
rect 20862 21646 20914 21698
rect 23774 21646 23826 21698
rect 26574 21646 26626 21698
rect 28702 21646 28754 21698
rect 4286 21534 4338 21586
rect 11454 21534 11506 21586
rect 11790 21534 11842 21586
rect 12126 21534 12178 21586
rect 16270 21534 16322 21586
rect 20414 21534 20466 21586
rect 20750 21534 20802 21586
rect 22654 21534 22706 21586
rect 23214 21534 23266 21586
rect 25230 21534 25282 21586
rect 25454 21534 25506 21586
rect 25790 21534 25842 21586
rect 27918 21534 27970 21586
rect 14926 21422 14978 21474
rect 16718 21422 16770 21474
rect 17390 21422 17442 21474
rect 18398 21422 18450 21474
rect 21534 21422 21586 21474
rect 23438 21422 23490 21474
rect 30830 21422 30882 21474
rect 1934 21310 1986 21362
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 9886 20862 9938 20914
rect 12014 20862 12066 20914
rect 13470 20862 13522 20914
rect 14814 20862 14866 20914
rect 16158 20862 16210 20914
rect 27918 20862 27970 20914
rect 40014 20862 40066 20914
rect 12798 20750 12850 20802
rect 13694 20750 13746 20802
rect 14030 20750 14082 20802
rect 14478 20750 14530 20802
rect 20078 20750 20130 20802
rect 21310 20750 21362 20802
rect 22206 20750 22258 20802
rect 22542 20750 22594 20802
rect 23550 20750 23602 20802
rect 29374 20750 29426 20802
rect 37662 20750 37714 20802
rect 13470 20638 13522 20690
rect 21422 20638 21474 20690
rect 22766 20638 22818 20690
rect 29038 20526 29090 20578
rect 29262 20526 29314 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 13918 20190 13970 20242
rect 12574 20078 12626 20130
rect 12686 20078 12738 20130
rect 13582 20078 13634 20130
rect 15598 20078 15650 20130
rect 16830 20078 16882 20130
rect 17502 20078 17554 20130
rect 17838 20078 17890 20130
rect 18174 20078 18226 20130
rect 21870 20078 21922 20130
rect 25454 20078 25506 20130
rect 26686 20078 26738 20130
rect 4286 19966 4338 20018
rect 12910 19966 12962 20018
rect 13358 19966 13410 20018
rect 14254 19966 14306 20018
rect 16606 19966 16658 20018
rect 19070 19966 19122 20018
rect 19406 19966 19458 20018
rect 25230 19966 25282 20018
rect 25678 19966 25730 20018
rect 25902 19966 25954 20018
rect 26238 19966 26290 20018
rect 26910 19966 26962 20018
rect 27918 19966 27970 20018
rect 37662 19966 37714 20018
rect 13134 19854 13186 19906
rect 16718 19854 16770 19906
rect 18510 19854 18562 19906
rect 26014 19854 26066 19906
rect 26462 19854 26514 19906
rect 27582 19854 27634 19906
rect 28702 19854 28754 19906
rect 30830 19854 30882 19906
rect 1934 19742 1986 19794
rect 12574 19742 12626 19794
rect 15486 19742 15538 19794
rect 15822 19742 15874 19794
rect 40014 19742 40066 19794
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 22878 19406 22930 19458
rect 1934 19294 1986 19346
rect 9886 19294 9938 19346
rect 12014 19294 12066 19346
rect 13582 19294 13634 19346
rect 15598 19294 15650 19346
rect 16382 19294 16434 19346
rect 21758 19294 21810 19346
rect 22766 19294 22818 19346
rect 26462 19294 26514 19346
rect 28590 19294 28642 19346
rect 4286 19182 4338 19234
rect 12798 19182 12850 19234
rect 15374 19182 15426 19234
rect 15486 19182 15538 19234
rect 16942 19182 16994 19234
rect 17502 19182 17554 19234
rect 17838 19182 17890 19234
rect 18958 19182 19010 19234
rect 19518 19182 19570 19234
rect 20750 19182 20802 19234
rect 21310 19182 21362 19234
rect 23886 19182 23938 19234
rect 24446 19182 24498 19234
rect 25790 19182 25842 19234
rect 29038 19182 29090 19234
rect 29374 19182 29426 19234
rect 29598 19182 29650 19234
rect 14590 19070 14642 19122
rect 16270 19070 16322 19122
rect 19294 19070 19346 19122
rect 19854 19070 19906 19122
rect 23214 19070 23266 19122
rect 14926 18958 14978 19010
rect 15710 18958 15762 19010
rect 15822 18958 15874 19010
rect 17166 18958 17218 19010
rect 17614 18958 17666 19010
rect 18622 18958 18674 19010
rect 20414 18958 20466 19010
rect 24334 18958 24386 19010
rect 24558 18958 24610 19010
rect 25006 18958 25058 19010
rect 29262 18958 29314 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 12350 18622 12402 18674
rect 19630 18622 19682 18674
rect 22318 18622 22370 18674
rect 22878 18622 22930 18674
rect 23326 18622 23378 18674
rect 23662 18622 23714 18674
rect 17838 18510 17890 18562
rect 18734 18510 18786 18562
rect 18846 18510 18898 18562
rect 20526 18510 20578 18562
rect 22766 18510 22818 18562
rect 23998 18510 24050 18562
rect 12574 18398 12626 18450
rect 13582 18398 13634 18450
rect 14366 18398 14418 18450
rect 18622 18398 18674 18450
rect 21422 18398 21474 18450
rect 21534 18398 21586 18450
rect 21982 18398 22034 18450
rect 24110 18398 24162 18450
rect 24222 18398 24274 18450
rect 24670 18398 24722 18450
rect 16494 18286 16546 18338
rect 17726 18286 17778 18338
rect 18062 18286 18114 18338
rect 20190 18286 20242 18338
rect 22654 18286 22706 18338
rect 28814 18286 28866 18338
rect 19294 18174 19346 18226
rect 20750 18174 20802 18226
rect 21086 18174 21138 18226
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 17390 17838 17442 17890
rect 17726 17838 17778 17890
rect 17614 17726 17666 17778
rect 18622 17726 18674 17778
rect 19518 17726 19570 17778
rect 22654 17726 22706 17778
rect 40014 17726 40066 17778
rect 20526 17614 20578 17666
rect 21198 17614 21250 17666
rect 21646 17614 21698 17666
rect 22542 17614 22594 17666
rect 23438 17614 23490 17666
rect 23886 17614 23938 17666
rect 24222 17614 24274 17666
rect 37662 17614 37714 17666
rect 17278 17502 17330 17554
rect 20750 17502 20802 17554
rect 21870 17502 21922 17554
rect 22878 17502 22930 17554
rect 24446 17502 24498 17554
rect 16718 17390 16770 17442
rect 18174 17390 18226 17442
rect 19070 17390 19122 17442
rect 21758 17390 21810 17442
rect 24558 17390 24610 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 19742 17054 19794 17106
rect 21534 17054 21586 17106
rect 21870 17054 21922 17106
rect 22542 17054 22594 17106
rect 24334 17054 24386 17106
rect 13806 16942 13858 16994
rect 22206 16942 22258 16994
rect 24222 16942 24274 16994
rect 26686 16942 26738 16994
rect 13134 16830 13186 16882
rect 16382 16830 16434 16882
rect 19966 16830 20018 16882
rect 24558 16830 24610 16882
rect 25118 16830 25170 16882
rect 25342 16830 25394 16882
rect 25454 16830 25506 16882
rect 25678 16830 25730 16882
rect 26238 16830 26290 16882
rect 26462 16830 26514 16882
rect 37886 16830 37938 16882
rect 15934 16718 15986 16770
rect 26574 16718 26626 16770
rect 40014 16606 40066 16658
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 27470 16270 27522 16322
rect 24894 16158 24946 16210
rect 27022 16158 27074 16210
rect 21310 16046 21362 16098
rect 24222 16046 24274 16098
rect 27358 15934 27410 15986
rect 21646 15822 21698 15874
rect 27470 15822 27522 15874
rect 28030 15822 28082 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 21310 15486 21362 15538
rect 21534 15486 21586 15538
rect 22318 15486 22370 15538
rect 22542 15486 22594 15538
rect 25454 15486 25506 15538
rect 29486 15486 29538 15538
rect 26910 15374 26962 15426
rect 21758 15262 21810 15314
rect 22094 15262 22146 15314
rect 25230 15262 25282 15314
rect 25566 15262 25618 15314
rect 25790 15262 25842 15314
rect 26126 15262 26178 15314
rect 37662 15262 37714 15314
rect 18398 15150 18450 15202
rect 29038 15150 29090 15202
rect 40014 15150 40066 15202
rect 21646 15038 21698 15090
rect 22654 15038 22706 15090
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 18958 14702 19010 14754
rect 16046 14590 16098 14642
rect 18174 14590 18226 14642
rect 26126 14590 26178 14642
rect 28254 14590 28306 14642
rect 29262 14590 29314 14642
rect 15374 14478 15426 14530
rect 18510 14478 18562 14530
rect 19294 14478 19346 14530
rect 20414 14478 20466 14530
rect 21646 14478 21698 14530
rect 22094 14478 22146 14530
rect 22542 14478 22594 14530
rect 22878 14478 22930 14530
rect 25342 14478 25394 14530
rect 18734 14366 18786 14418
rect 20078 14366 20130 14418
rect 20638 14366 20690 14418
rect 22318 14366 22370 14418
rect 18622 14254 18674 14306
rect 20190 14254 20242 14306
rect 21870 14254 21922 14306
rect 22766 14254 22818 14306
rect 23438 14254 23490 14306
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 17502 13918 17554 13970
rect 18286 13918 18338 13970
rect 18846 13918 18898 13970
rect 19518 13918 19570 13970
rect 20078 13918 20130 13970
rect 26686 13918 26738 13970
rect 26910 13918 26962 13970
rect 14702 13806 14754 13858
rect 19742 13806 19794 13858
rect 19854 13806 19906 13858
rect 21086 13806 21138 13858
rect 25230 13806 25282 13858
rect 27022 13806 27074 13858
rect 14030 13694 14082 13746
rect 20414 13694 20466 13746
rect 23662 13694 23714 13746
rect 23886 13694 23938 13746
rect 24110 13694 24162 13746
rect 25342 13694 25394 13746
rect 25566 13694 25618 13746
rect 16830 13582 16882 13634
rect 17950 13582 18002 13634
rect 18174 13582 18226 13634
rect 23214 13582 23266 13634
rect 17278 13470 17330 13522
rect 23550 13470 23602 13522
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 17614 13022 17666 13074
rect 18622 13022 18674 13074
rect 20750 13022 20802 13074
rect 23438 13022 23490 13074
rect 25566 13022 25618 13074
rect 26126 13022 26178 13074
rect 17838 12910 17890 12962
rect 22654 12910 22706 12962
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 40238 9102 40290 9154
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 25566 4286 25618 4338
rect 26238 4062 26290 4114
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 18622 3614 18674 3666
rect 25566 3614 25618 3666
rect 18062 3502 18114 3554
rect 20750 3502 20802 3554
rect 24558 3502 24610 3554
rect 21758 3278 21810 3330
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
<< metal2 >>
rect 16128 41200 16240 42000
rect 16800 41200 16912 42000
rect 17472 41200 17584 42000
rect 20832 41200 20944 42000
rect 23520 41200 23632 42000
rect 26880 41200 26992 42000
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 16156 36708 16212 41200
rect 16828 37492 16884 41200
rect 17500 38276 17556 41200
rect 17500 38210 17556 38220
rect 18620 38276 18676 38286
rect 18620 38182 18676 38220
rect 20860 38276 20916 41200
rect 20860 38210 20916 38220
rect 22092 38276 22148 38286
rect 22092 38182 22148 38220
rect 23548 38276 23604 41200
rect 23548 38210 23604 38220
rect 25564 38276 25620 38286
rect 25564 38182 25620 38220
rect 16828 37426 16884 37436
rect 18060 38050 18116 38062
rect 18060 37998 18062 38050
rect 18114 37998 18116 38050
rect 17388 37268 17444 37278
rect 16156 36642 16212 36652
rect 17276 37266 17444 37268
rect 17276 37214 17390 37266
rect 17442 37214 17444 37266
rect 17276 37212 17444 37214
rect 16380 36482 16436 36494
rect 16380 36430 16382 36482
rect 16434 36430 16436 36482
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 16380 31948 16436 36430
rect 16268 31892 16436 31948
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 16156 28530 16212 28542
rect 16156 28478 16158 28530
rect 16210 28478 16212 28530
rect 13916 27860 13972 27870
rect 13916 27766 13972 27804
rect 14364 27860 14420 27870
rect 10892 27636 10948 27646
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 4284 24724 4340 24734
rect 4284 24630 4340 24668
rect 1932 24500 1988 24510
rect 1932 24406 1988 24444
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 1932 24050 1988 24062
rect 1932 23998 1934 24050
rect 1986 23998 1988 24050
rect 1932 23604 1988 23998
rect 9996 24052 10052 24062
rect 9996 23958 10052 23996
rect 4284 23940 4340 23950
rect 4284 23846 4340 23884
rect 1932 23538 1988 23548
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 4284 21588 4340 21598
rect 4284 21494 4340 21532
rect 9884 21588 9940 21598
rect 1932 21362 1988 21374
rect 1932 21310 1934 21362
rect 1986 21310 1988 21362
rect 1932 20916 1988 21310
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 1932 20850 1988 20860
rect 9884 20914 9940 21532
rect 9884 20862 9886 20914
rect 9938 20862 9940 20914
rect 9884 20692 9940 20862
rect 9884 20626 9940 20636
rect 10892 20132 10948 27580
rect 12908 27076 12964 27086
rect 12796 24052 12852 24062
rect 12124 23828 12180 23838
rect 12124 23734 12180 23772
rect 12796 23378 12852 23996
rect 12908 23940 12964 27020
rect 14364 27076 14420 27804
rect 14700 27748 14756 27758
rect 14700 27654 14756 27692
rect 16156 27300 16212 28478
rect 16268 28532 16324 31892
rect 16268 28438 16324 28476
rect 16940 28532 16996 28542
rect 16996 28476 17220 28532
rect 16940 28438 16996 28476
rect 16492 28418 16548 28430
rect 16492 28366 16494 28418
rect 16546 28366 16548 28418
rect 16156 27234 16212 27244
rect 16380 27860 16436 27870
rect 14364 26982 14420 27020
rect 15036 26964 15092 26974
rect 15036 26870 15092 26908
rect 16380 24948 16436 27804
rect 16492 27076 16548 28366
rect 16828 27746 16884 27758
rect 16828 27694 16830 27746
rect 16882 27694 16884 27746
rect 16828 27636 16884 27694
rect 16828 27570 16884 27580
rect 17164 27186 17220 28476
rect 17276 28530 17332 37212
rect 17388 37202 17444 37212
rect 17388 36708 17444 36718
rect 17388 36614 17444 36652
rect 18060 31948 18116 37998
rect 21308 38050 21364 38062
rect 21308 37998 21310 38050
rect 21362 37998 21364 38050
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 18396 37492 18452 37502
rect 18396 37398 18452 37436
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 18060 31892 18452 31948
rect 17612 29316 17668 29326
rect 17612 29314 18116 29316
rect 17612 29262 17614 29314
rect 17666 29262 18116 29314
rect 17612 29260 18116 29262
rect 17612 29250 17668 29260
rect 18060 28756 18116 29260
rect 18396 28868 18452 31892
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 18396 28812 18564 28868
rect 18060 28754 18452 28756
rect 18060 28702 18062 28754
rect 18114 28702 18452 28754
rect 18060 28700 18452 28702
rect 18060 28690 18116 28700
rect 17276 28478 17278 28530
rect 17330 28478 17332 28530
rect 17276 28466 17332 28478
rect 17388 28028 18340 28084
rect 17388 27970 17444 28028
rect 17388 27918 17390 27970
rect 17442 27918 17444 27970
rect 17388 27906 17444 27918
rect 17724 27858 17780 27870
rect 17724 27806 17726 27858
rect 17778 27806 17780 27858
rect 17500 27748 17556 27758
rect 17500 27654 17556 27692
rect 17388 27300 17444 27310
rect 17164 27134 17166 27186
rect 17218 27134 17220 27186
rect 17164 27122 17220 27134
rect 17276 27244 17388 27300
rect 16492 27010 16548 27020
rect 15932 24946 16436 24948
rect 15932 24894 16382 24946
rect 16434 24894 16436 24946
rect 15932 24892 16436 24894
rect 15932 24722 15988 24892
rect 15932 24670 15934 24722
rect 15986 24670 15988 24722
rect 15932 24658 15988 24670
rect 13020 24612 13076 24622
rect 15148 24612 15204 24622
rect 13020 24518 13076 24556
rect 14812 24610 15204 24612
rect 14812 24558 15150 24610
rect 15202 24558 15204 24610
rect 14812 24556 15204 24558
rect 14812 24162 14868 24556
rect 15148 24546 15204 24556
rect 16156 24612 16212 24622
rect 14812 24110 14814 24162
rect 14866 24110 14868 24162
rect 14812 24098 14868 24110
rect 16156 24162 16212 24556
rect 16156 24110 16158 24162
rect 16210 24110 16212 24162
rect 16156 24098 16212 24110
rect 13804 24052 13860 24062
rect 12908 23938 13412 23940
rect 12908 23886 12910 23938
rect 12962 23886 13412 23938
rect 12908 23884 13412 23886
rect 12908 23874 12964 23884
rect 12796 23326 12798 23378
rect 12850 23326 12852 23378
rect 12796 23314 12852 23326
rect 13020 23604 13076 23614
rect 13020 23378 13076 23548
rect 13020 23326 13022 23378
rect 13074 23326 13076 23378
rect 13020 23314 13076 23326
rect 13356 23378 13412 23884
rect 13804 23938 13860 23996
rect 15260 24052 15316 24062
rect 15820 24052 15876 24062
rect 15260 24050 15876 24052
rect 15260 23998 15262 24050
rect 15314 23998 15822 24050
rect 15874 23998 15876 24050
rect 15260 23996 15876 23998
rect 15260 23986 15316 23996
rect 15820 23986 15876 23996
rect 13804 23886 13806 23938
rect 13858 23886 13860 23938
rect 13804 23874 13860 23886
rect 13916 23938 13972 23950
rect 13916 23886 13918 23938
rect 13970 23886 13972 23938
rect 13468 23826 13524 23838
rect 13468 23774 13470 23826
rect 13522 23774 13524 23826
rect 13468 23604 13524 23774
rect 13580 23828 13636 23838
rect 13580 23734 13636 23772
rect 13468 23538 13524 23548
rect 13356 23326 13358 23378
rect 13410 23326 13412 23378
rect 13356 23314 13412 23326
rect 13916 23492 13972 23886
rect 14924 23938 14980 23950
rect 14924 23886 14926 23938
rect 14978 23886 14980 23938
rect 14140 23604 14196 23614
rect 12684 23156 12740 23166
rect 12684 23062 12740 23100
rect 13916 22708 13972 23436
rect 13468 22652 13972 22708
rect 14028 23548 14140 23604
rect 11564 22260 11620 22270
rect 11564 21810 11620 22204
rect 13356 22148 13412 22158
rect 11564 21758 11566 21810
rect 11618 21758 11620 21810
rect 11564 21746 11620 21758
rect 12796 22146 13412 22148
rect 12796 22094 13358 22146
rect 13410 22094 13412 22146
rect 12796 22092 13412 22094
rect 12796 21698 12852 22092
rect 13356 22082 13412 22092
rect 13468 21924 13524 22652
rect 14028 22596 14084 23548
rect 14140 23538 14196 23548
rect 14924 23492 14980 23886
rect 15148 23940 15204 23950
rect 15148 23846 15204 23884
rect 14924 23426 14980 23436
rect 15596 23828 15652 23838
rect 13580 22540 14084 22596
rect 14140 23156 14196 23166
rect 13580 22260 13636 22540
rect 13580 22166 13636 22204
rect 13692 22260 13748 22270
rect 13916 22260 13972 22270
rect 14140 22260 14196 23100
rect 15596 22932 15652 23772
rect 15708 23826 15764 23838
rect 15708 23774 15710 23826
rect 15762 23774 15764 23826
rect 15708 23268 15764 23774
rect 15932 23828 15988 23838
rect 15932 23734 15988 23772
rect 15932 23492 15988 23502
rect 15932 23378 15988 23436
rect 15932 23326 15934 23378
rect 15986 23326 15988 23378
rect 15932 23314 15988 23326
rect 16044 23380 16100 23390
rect 15820 23268 15876 23278
rect 15708 23266 15876 23268
rect 15708 23214 15822 23266
rect 15874 23214 15876 23266
rect 15708 23212 15876 23214
rect 15820 23156 15876 23212
rect 16044 23266 16100 23324
rect 16044 23214 16046 23266
rect 16098 23214 16100 23266
rect 16044 23202 16100 23214
rect 15876 23100 15988 23156
rect 15820 23090 15876 23100
rect 15596 22876 15876 22932
rect 13692 22258 13972 22260
rect 13692 22206 13694 22258
rect 13746 22206 13918 22258
rect 13970 22206 13972 22258
rect 13692 22204 13972 22206
rect 13692 22194 13748 22204
rect 13916 22194 13972 22204
rect 14028 22258 14196 22260
rect 14028 22206 14142 22258
rect 14194 22206 14196 22258
rect 14028 22204 14196 22206
rect 13468 21868 13636 21924
rect 12796 21646 12798 21698
rect 12850 21646 12852 21698
rect 12796 21634 12852 21646
rect 11452 21588 11508 21598
rect 11452 21494 11508 21532
rect 11788 21588 11844 21598
rect 11788 21586 12068 21588
rect 11788 21534 11790 21586
rect 11842 21534 12068 21586
rect 11788 21532 12068 21534
rect 11788 21522 11844 21532
rect 12012 20914 12068 21532
rect 12012 20862 12014 20914
rect 12066 20862 12068 20914
rect 12012 20850 12068 20862
rect 12124 21586 12180 21598
rect 12124 21534 12126 21586
rect 12178 21534 12180 21586
rect 12124 20916 12180 21534
rect 13468 21588 13524 21598
rect 12124 20850 12180 20860
rect 12796 20916 12852 20926
rect 12796 20802 12852 20860
rect 12796 20750 12798 20802
rect 12850 20750 12852 20802
rect 12796 20738 12852 20750
rect 13356 20916 13412 20926
rect 13356 20188 13412 20860
rect 13468 20914 13524 21532
rect 13468 20862 13470 20914
rect 13522 20862 13524 20914
rect 13468 20850 13524 20862
rect 13468 20692 13524 20702
rect 13468 20598 13524 20636
rect 10892 20066 10948 20076
rect 12572 20130 12628 20142
rect 12572 20078 12574 20130
rect 12626 20078 12628 20130
rect 4284 20020 4340 20030
rect 4284 19926 4340 19964
rect 9884 20020 9940 20030
rect 1932 19796 1988 19806
rect 1932 19702 1988 19740
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 1932 19346 1988 19358
rect 1932 19294 1934 19346
rect 1986 19294 1988 19346
rect 1932 18900 1988 19294
rect 9884 19346 9940 19964
rect 12460 20020 12516 20030
rect 12572 20020 12628 20078
rect 12516 19964 12628 20020
rect 12684 20130 12740 20142
rect 13356 20132 13524 20188
rect 12684 20078 12686 20130
rect 12738 20078 12740 20130
rect 12684 20020 12740 20078
rect 12348 19908 12404 19918
rect 9884 19294 9886 19346
rect 9938 19294 9940 19346
rect 9884 19282 9940 19294
rect 12012 19852 12348 19908
rect 12012 19346 12068 19852
rect 12348 19842 12404 19852
rect 12012 19294 12014 19346
rect 12066 19294 12068 19346
rect 12012 19282 12068 19294
rect 4284 19236 4340 19246
rect 4284 19142 4340 19180
rect 12348 19236 12404 19246
rect 1932 18834 1988 18844
rect 12348 18674 12404 19180
rect 12348 18622 12350 18674
rect 12402 18622 12404 18674
rect 12348 18610 12404 18622
rect 12460 18452 12516 19964
rect 12684 19954 12740 19964
rect 12908 20018 12964 20030
rect 12908 19966 12910 20018
rect 12962 19966 12964 20018
rect 12572 19796 12628 19806
rect 12908 19796 12964 19966
rect 13356 20018 13412 20030
rect 13356 19966 13358 20018
rect 13410 19966 13412 20018
rect 13132 19908 13188 19918
rect 13132 19814 13188 19852
rect 12572 19794 12964 19796
rect 12572 19742 12574 19794
rect 12626 19742 12964 19794
rect 12572 19740 12964 19742
rect 12572 19730 12628 19740
rect 13356 19572 13412 19966
rect 13356 19506 13412 19516
rect 13468 19348 13524 20132
rect 13580 20130 13636 21868
rect 14028 21252 14084 22204
rect 14140 22194 14196 22204
rect 14252 22258 14308 22270
rect 14252 22206 14254 22258
rect 14306 22206 14308 22258
rect 14252 21924 14308 22206
rect 14252 21858 14308 21868
rect 14924 22148 14980 22158
rect 14924 21474 14980 22092
rect 15372 21812 15428 21822
rect 14924 21422 14926 21474
rect 14978 21422 14980 21474
rect 14924 21410 14980 21422
rect 15036 21756 15372 21812
rect 13580 20078 13582 20130
rect 13634 20078 13636 20130
rect 13580 20066 13636 20078
rect 13692 21196 14084 21252
rect 13692 20802 13748 21196
rect 14812 20916 14868 20926
rect 15036 20916 15092 21756
rect 15372 21718 15428 21756
rect 14868 20860 15092 20916
rect 15148 21588 15204 21598
rect 14812 20822 14868 20860
rect 13692 20750 13694 20802
rect 13746 20750 13748 20802
rect 13692 20188 13748 20750
rect 14028 20804 14084 20814
rect 14476 20804 14532 20814
rect 14028 20802 14532 20804
rect 14028 20750 14030 20802
rect 14082 20750 14478 20802
rect 14530 20750 14532 20802
rect 14028 20748 14532 20750
rect 14028 20738 14084 20748
rect 13916 20244 13972 20254
rect 13804 20242 13972 20244
rect 13804 20190 13918 20242
rect 13970 20190 13972 20242
rect 13804 20188 13972 20190
rect 13692 20132 13860 20188
rect 13916 20178 13972 20188
rect 13692 20020 13748 20132
rect 13692 19954 13748 19964
rect 14252 20020 14308 20030
rect 14252 19926 14308 19964
rect 13580 19348 13636 19358
rect 12796 19346 13636 19348
rect 12796 19294 13582 19346
rect 13634 19294 13636 19346
rect 12796 19292 13636 19294
rect 12796 19234 12852 19292
rect 12796 19182 12798 19234
rect 12850 19182 12852 19234
rect 12796 19170 12852 19182
rect 12572 18452 12628 18462
rect 12460 18450 12628 18452
rect 12460 18398 12574 18450
rect 12626 18398 12628 18450
rect 12460 18396 12628 18398
rect 12572 18386 12628 18396
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 13132 16884 13188 19292
rect 13580 18450 13636 19292
rect 13580 18398 13582 18450
rect 13634 18398 13636 18450
rect 13580 18386 13636 18398
rect 14364 19124 14420 19134
rect 14476 19124 14532 20748
rect 15148 19908 15204 21532
rect 15596 20130 15652 20142
rect 15596 20078 15598 20130
rect 15650 20078 15652 20130
rect 15596 20020 15652 20078
rect 15596 19954 15652 19964
rect 15148 19842 15204 19852
rect 15484 19794 15540 19806
rect 15484 19742 15486 19794
rect 15538 19742 15540 19794
rect 15372 19234 15428 19246
rect 15372 19182 15374 19234
rect 15426 19182 15428 19234
rect 14588 19124 14644 19134
rect 14476 19122 14644 19124
rect 14476 19070 14590 19122
rect 14642 19070 14644 19122
rect 14476 19068 14644 19070
rect 14364 18450 14420 19068
rect 14588 19012 14644 19068
rect 15372 19124 15428 19182
rect 15484 19234 15540 19742
rect 15820 19796 15876 22876
rect 15932 22596 15988 23100
rect 15932 22540 16100 22596
rect 15820 19794 15988 19796
rect 15820 19742 15822 19794
rect 15874 19742 15988 19794
rect 15820 19740 15988 19742
rect 15820 19730 15876 19740
rect 15596 19572 15652 19582
rect 15596 19346 15652 19516
rect 15596 19294 15598 19346
rect 15650 19294 15652 19346
rect 15596 19282 15652 19294
rect 15484 19182 15486 19234
rect 15538 19182 15540 19234
rect 15484 19170 15540 19182
rect 15372 19058 15428 19068
rect 14588 18946 14644 18956
rect 14924 19010 14980 19022
rect 14924 18958 14926 19010
rect 14978 18958 14980 19010
rect 14924 18564 14980 18958
rect 15708 19012 15764 19022
rect 15708 18918 15764 18956
rect 15820 19010 15876 19022
rect 15820 18958 15822 19010
rect 15874 18958 15876 19010
rect 14924 18498 14980 18508
rect 14364 18398 14366 18450
rect 14418 18398 14420 18450
rect 14364 18386 14420 18398
rect 15820 18452 15876 18958
rect 15820 18386 15876 18396
rect 13804 17556 13860 17566
rect 13804 16994 13860 17500
rect 15932 17108 15988 19740
rect 16044 19012 16100 22540
rect 16268 21924 16324 24892
rect 16380 24882 16436 24892
rect 17276 24946 17332 27244
rect 17388 27234 17444 27244
rect 17388 27076 17444 27086
rect 17388 26982 17444 27020
rect 17612 26964 17668 26974
rect 17612 26870 17668 26908
rect 17724 26740 17780 27806
rect 17948 27858 18004 27870
rect 17948 27806 17950 27858
rect 18002 27806 18004 27858
rect 17948 27076 18004 27806
rect 17948 26982 18004 27020
rect 18284 27074 18340 28028
rect 18396 27860 18452 28700
rect 18508 28084 18564 28812
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 18508 28028 18676 28084
rect 18508 27860 18564 27898
rect 18396 27804 18508 27860
rect 18508 27794 18564 27804
rect 18284 27022 18286 27074
rect 18338 27022 18340 27074
rect 18284 27010 18340 27022
rect 18508 27636 18564 27646
rect 18620 27636 18676 28028
rect 18564 27580 18676 27636
rect 19068 27860 19124 27870
rect 17500 26684 17780 26740
rect 17836 26962 17892 26974
rect 17836 26910 17838 26962
rect 17890 26910 17892 26962
rect 17500 26514 17556 26684
rect 17500 26462 17502 26514
rect 17554 26462 17556 26514
rect 17500 26450 17556 26462
rect 17836 26404 17892 26910
rect 18508 26962 18564 27580
rect 18620 27300 18676 27310
rect 18620 27074 18676 27244
rect 19068 27186 19124 27804
rect 19180 27748 19236 27758
rect 21308 27748 21364 37998
rect 24556 38050 24612 38062
rect 24556 37998 24558 38050
rect 24610 37998 24612 38050
rect 24556 31948 24612 37998
rect 26908 37492 26964 41200
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 26908 37426 26964 37436
rect 28140 37492 28196 37502
rect 28140 37398 28196 37436
rect 19180 27746 19684 27748
rect 19180 27694 19182 27746
rect 19234 27694 19684 27746
rect 19180 27692 19684 27694
rect 19180 27682 19236 27692
rect 19628 27298 19684 27692
rect 19628 27246 19630 27298
rect 19682 27246 19684 27298
rect 19628 27234 19684 27246
rect 20524 27746 21364 27748
rect 20524 27694 21310 27746
rect 21362 27694 21364 27746
rect 20524 27692 21364 27694
rect 19068 27134 19070 27186
rect 19122 27134 19124 27186
rect 19068 27122 19124 27134
rect 18620 27022 18622 27074
rect 18674 27022 18676 27074
rect 18620 27010 18676 27022
rect 19628 27076 19684 27086
rect 19628 26982 19684 27020
rect 18508 26910 18510 26962
rect 18562 26910 18564 26962
rect 18508 26898 18564 26910
rect 19964 26962 20020 26974
rect 19964 26910 19966 26962
rect 20018 26910 20020 26962
rect 19964 26852 20020 26910
rect 19964 26796 20468 26852
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 20412 26514 20468 26796
rect 20412 26462 20414 26514
rect 20466 26462 20468 26514
rect 20412 26450 20468 26462
rect 20524 26514 20580 27692
rect 21308 27682 21364 27692
rect 24220 31892 24612 31948
rect 27580 37266 27636 37278
rect 27580 37214 27582 37266
rect 27634 37214 27636 37266
rect 27580 31948 27636 37214
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 40236 36372 40292 36382
rect 40236 36278 40292 36316
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 27580 31892 28196 31948
rect 24220 27188 24276 31892
rect 23772 27186 24276 27188
rect 23772 27134 24222 27186
rect 24274 27134 24276 27186
rect 23772 27132 24276 27134
rect 21420 27076 21476 27086
rect 21420 26982 21476 27020
rect 20524 26462 20526 26514
rect 20578 26462 20580 26514
rect 20524 26450 20580 26462
rect 20860 26964 20916 26974
rect 18060 26404 18116 26414
rect 17836 26348 18060 26404
rect 18060 26290 18116 26348
rect 18508 26404 18564 26414
rect 18508 26310 18564 26348
rect 20636 26402 20692 26414
rect 20636 26350 20638 26402
rect 20690 26350 20692 26402
rect 18060 26238 18062 26290
rect 18114 26238 18116 26290
rect 18060 26226 18116 26238
rect 18732 26290 18788 26302
rect 18732 26238 18734 26290
rect 18786 26238 18788 26290
rect 17836 26068 17892 26078
rect 17836 26066 18228 26068
rect 17836 26014 17838 26066
rect 17890 26014 18228 26066
rect 17836 26012 18228 26014
rect 17836 26002 17892 26012
rect 17276 24894 17278 24946
rect 17330 24894 17332 24946
rect 17276 24882 17332 24894
rect 17500 24948 17556 24958
rect 17500 24946 17892 24948
rect 17500 24894 17502 24946
rect 17554 24894 17892 24946
rect 17500 24892 17892 24894
rect 17500 24882 17556 24892
rect 16940 24724 16996 24734
rect 17612 24724 17668 24734
rect 16940 24052 16996 24668
rect 16940 23958 16996 23996
rect 17500 24722 17668 24724
rect 17500 24670 17614 24722
rect 17666 24670 17668 24722
rect 17500 24668 17668 24670
rect 16492 23938 16548 23950
rect 16492 23886 16494 23938
rect 16546 23886 16548 23938
rect 16492 23828 16548 23886
rect 16492 23762 16548 23772
rect 17388 23714 17444 23726
rect 17388 23662 17390 23714
rect 17442 23662 17444 23714
rect 16716 23380 16772 23390
rect 16716 22594 16772 23324
rect 17388 23380 17444 23662
rect 17500 23716 17556 24668
rect 17612 24658 17668 24668
rect 17612 23940 17668 23950
rect 17612 23846 17668 23884
rect 17836 23828 17892 24892
rect 17948 23940 18004 23950
rect 17948 23846 18004 23884
rect 18172 23938 18228 26012
rect 18172 23886 18174 23938
rect 18226 23886 18228 23938
rect 17500 23650 17556 23660
rect 17724 23716 17780 23726
rect 17836 23716 17892 23772
rect 17836 23660 18004 23716
rect 17724 23622 17780 23660
rect 17388 23314 17444 23324
rect 16716 22542 16718 22594
rect 16770 22542 16772 22594
rect 16716 22530 16772 22542
rect 16716 22372 16772 22382
rect 16156 21868 16324 21924
rect 16604 22260 16660 22270
rect 16156 21812 16212 21868
rect 16156 20914 16212 21756
rect 16380 21812 16436 21822
rect 16156 20862 16158 20914
rect 16210 20862 16212 20914
rect 16156 20850 16212 20862
rect 16268 21586 16324 21598
rect 16268 21534 16270 21586
rect 16322 21534 16324 21586
rect 16268 21476 16324 21534
rect 16268 20188 16324 21420
rect 16044 18946 16100 18956
rect 16156 20132 16324 20188
rect 16044 17108 16100 17118
rect 15932 17052 16044 17108
rect 16044 17042 16100 17052
rect 13804 16942 13806 16994
rect 13858 16942 13860 16994
rect 13804 16930 13860 16942
rect 13132 16790 13188 16828
rect 15372 16884 15428 16894
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 14028 14532 14084 14542
rect 14028 13746 14084 14476
rect 15372 14532 15428 16828
rect 15932 16772 15988 16782
rect 16156 16772 16212 20132
rect 16380 19346 16436 21756
rect 16604 21476 16660 22204
rect 16716 22148 16772 22316
rect 17276 22370 17332 22382
rect 17276 22318 17278 22370
rect 17330 22318 17332 22370
rect 16828 22260 16884 22270
rect 17276 22260 17332 22318
rect 17836 22372 17892 22382
rect 17836 22278 17892 22316
rect 16828 22258 17108 22260
rect 16828 22206 16830 22258
rect 16882 22206 17108 22258
rect 16828 22204 17108 22206
rect 16828 22194 16884 22204
rect 16716 22054 16772 22092
rect 16940 22036 16996 22046
rect 16716 21476 16772 21486
rect 16604 21474 16772 21476
rect 16604 21422 16718 21474
rect 16770 21422 16772 21474
rect 16604 21420 16772 21422
rect 16716 21410 16772 21420
rect 16828 20130 16884 20142
rect 16828 20078 16830 20130
rect 16882 20078 16884 20130
rect 16604 20018 16660 20030
rect 16604 19966 16606 20018
rect 16658 19966 16660 20018
rect 16604 19796 16660 19966
rect 16716 19908 16772 19918
rect 16716 19814 16772 19852
rect 16604 19730 16660 19740
rect 16380 19294 16382 19346
rect 16434 19294 16436 19346
rect 16380 19282 16436 19294
rect 16492 19236 16548 19246
rect 16268 19124 16324 19134
rect 16268 19030 16324 19068
rect 16492 18338 16548 19180
rect 16828 19124 16884 20078
rect 16828 19058 16884 19068
rect 16940 19234 16996 21980
rect 17052 21924 17108 22204
rect 17276 22194 17332 22204
rect 17500 22148 17556 22158
rect 17500 22054 17556 22092
rect 17052 21868 17556 21924
rect 17500 21812 17556 21868
rect 17836 21812 17892 21822
rect 17500 21810 17892 21812
rect 17500 21758 17502 21810
rect 17554 21758 17838 21810
rect 17890 21758 17892 21810
rect 17500 21756 17892 21758
rect 17500 21746 17556 21756
rect 17836 21746 17892 21756
rect 17388 21476 17444 21486
rect 17388 21382 17444 21420
rect 17500 20132 17556 20142
rect 17500 20038 17556 20076
rect 17836 20130 17892 20142
rect 17836 20078 17838 20130
rect 17890 20078 17892 20130
rect 17836 20020 17892 20078
rect 17836 19954 17892 19964
rect 16940 19182 16942 19234
rect 16994 19182 16996 19234
rect 16940 18564 16996 19182
rect 17500 19236 17556 19246
rect 17500 19142 17556 19180
rect 17836 19234 17892 19246
rect 17836 19182 17838 19234
rect 17890 19182 17892 19234
rect 17836 19124 17892 19182
rect 17836 19058 17892 19068
rect 16940 18498 16996 18508
rect 17164 19010 17220 19022
rect 17164 18958 17166 19010
rect 17218 18958 17220 19010
rect 16492 18286 16494 18338
rect 16546 18286 16548 18338
rect 16492 18274 16548 18286
rect 17164 18340 17220 18958
rect 17612 19012 17668 19022
rect 17612 18918 17668 18956
rect 17836 18564 17892 18574
rect 17948 18564 18004 23660
rect 18060 23156 18116 23166
rect 18060 23062 18116 23100
rect 18172 23044 18228 23886
rect 18732 23940 18788 26238
rect 20300 26290 20356 26302
rect 20300 26238 20302 26290
rect 20354 26238 20356 26290
rect 19628 25396 19684 25406
rect 19516 25340 19628 25396
rect 18732 23378 18788 23884
rect 18732 23326 18734 23378
rect 18786 23326 18788 23378
rect 18732 23314 18788 23326
rect 18844 23884 19460 23940
rect 18172 22978 18228 22988
rect 18284 23266 18340 23278
rect 18508 23268 18564 23278
rect 18284 23214 18286 23266
rect 18338 23214 18340 23266
rect 18172 22258 18228 22270
rect 18172 22206 18174 22258
rect 18226 22206 18228 22258
rect 18172 21924 18228 22206
rect 18284 22260 18340 23214
rect 18284 22194 18340 22204
rect 18396 23266 18564 23268
rect 18396 23214 18510 23266
rect 18562 23214 18564 23266
rect 18396 23212 18564 23214
rect 18396 21924 18452 23212
rect 18508 23202 18564 23212
rect 18620 23156 18676 23166
rect 18620 22482 18676 23100
rect 18620 22430 18622 22482
rect 18674 22430 18676 22482
rect 18620 22418 18676 22430
rect 18732 22372 18788 22382
rect 18508 22258 18564 22270
rect 18508 22206 18510 22258
rect 18562 22206 18564 22258
rect 18508 22148 18564 22206
rect 18732 22258 18788 22316
rect 18732 22206 18734 22258
rect 18786 22206 18788 22258
rect 18732 22194 18788 22206
rect 18508 22082 18564 22092
rect 18172 21868 18564 21924
rect 18508 21588 18564 21868
rect 18508 21522 18564 21532
rect 18396 21476 18452 21486
rect 18396 21382 18452 21420
rect 18172 20692 18228 20702
rect 18172 20130 18228 20636
rect 18172 20078 18174 20130
rect 18226 20078 18228 20130
rect 18172 20066 18228 20078
rect 18508 19906 18564 19918
rect 18508 19854 18510 19906
rect 18562 19854 18564 19906
rect 18508 19796 18564 19854
rect 18564 19740 18788 19796
rect 18508 19730 18564 19740
rect 18620 19012 18676 19022
rect 17836 18562 18004 18564
rect 17836 18510 17838 18562
rect 17890 18510 18004 18562
rect 17836 18508 18004 18510
rect 18508 19010 18676 19012
rect 18508 18958 18622 19010
rect 18674 18958 18676 19010
rect 18508 18956 18676 18958
rect 17164 18274 17220 18284
rect 17388 18452 17444 18462
rect 17388 17890 17444 18396
rect 17724 18452 17780 18462
rect 17724 18338 17780 18396
rect 17724 18286 17726 18338
rect 17778 18286 17780 18338
rect 17724 18274 17780 18286
rect 17388 17838 17390 17890
rect 17442 17838 17444 17890
rect 17388 17826 17444 17838
rect 17724 17892 17780 17902
rect 17724 17798 17780 17836
rect 17612 17780 17668 17790
rect 17612 17686 17668 17724
rect 17276 17556 17332 17566
rect 17276 17462 17332 17500
rect 17836 17556 17892 18508
rect 18060 18340 18116 18350
rect 18060 18246 18116 18284
rect 17836 17490 17892 17500
rect 16716 17442 16772 17454
rect 16716 17390 16718 17442
rect 16770 17390 16772 17442
rect 16380 16884 16436 16894
rect 16716 16884 16772 17390
rect 16436 16828 16772 16884
rect 18172 17444 18228 17454
rect 16380 16790 16436 16828
rect 15932 16770 16212 16772
rect 15932 16718 15934 16770
rect 15986 16718 16212 16770
rect 15932 16716 16212 16718
rect 15932 16706 15988 16716
rect 16044 15540 16100 15550
rect 16044 14642 16100 15484
rect 16044 14590 16046 14642
rect 16098 14590 16100 14642
rect 16044 14578 16100 14590
rect 18172 14642 18228 17388
rect 18508 15540 18564 18956
rect 18620 18946 18676 18956
rect 18732 18676 18788 19740
rect 18844 19124 18900 23884
rect 19404 23826 19460 23884
rect 19404 23774 19406 23826
rect 19458 23774 19460 23826
rect 19404 23762 19460 23774
rect 19292 23714 19348 23726
rect 19292 23662 19294 23714
rect 19346 23662 19348 23714
rect 19292 23268 19348 23662
rect 19404 23268 19460 23278
rect 19068 23266 19460 23268
rect 19068 23214 19406 23266
rect 19458 23214 19460 23266
rect 19068 23212 19460 23214
rect 19068 20188 19124 23212
rect 19404 23202 19460 23212
rect 19292 23044 19348 23054
rect 19292 22950 19348 22988
rect 19292 22370 19348 22382
rect 19292 22318 19294 22370
rect 19346 22318 19348 22370
rect 19292 22148 19348 22318
rect 19292 22082 19348 22092
rect 18956 20132 19124 20188
rect 19180 21476 19236 21486
rect 18956 19234 19012 20132
rect 18956 19182 18958 19234
rect 19010 19182 19012 19234
rect 18956 19170 19012 19182
rect 19068 20018 19124 20030
rect 19068 19966 19070 20018
rect 19122 19966 19124 20018
rect 19068 19236 19124 19966
rect 19068 19170 19124 19180
rect 18844 19058 18900 19068
rect 18732 18562 18788 18620
rect 18956 19012 19012 19022
rect 18732 18510 18734 18562
rect 18786 18510 18788 18562
rect 18732 18498 18788 18510
rect 18844 18564 18900 18574
rect 18844 18470 18900 18508
rect 18620 18452 18676 18462
rect 18620 17778 18676 18396
rect 18956 18004 19012 18956
rect 18620 17726 18622 17778
rect 18674 17726 18676 17778
rect 18620 17714 18676 17726
rect 18732 17948 19012 18004
rect 18620 15540 18676 15550
rect 18508 15484 18620 15540
rect 18620 15474 18676 15484
rect 18732 15316 18788 17948
rect 18956 17780 19012 17790
rect 18508 15260 18900 15316
rect 18172 14590 18174 14642
rect 18226 14590 18228 14642
rect 18172 14578 18228 14590
rect 18396 15202 18452 15214
rect 18396 15150 18398 15202
rect 18450 15150 18452 15202
rect 14700 14308 14756 14318
rect 14700 13858 14756 14252
rect 15372 13972 15428 14476
rect 18284 14420 18340 14430
rect 15372 13906 15428 13916
rect 17500 13972 17556 13982
rect 14700 13806 14702 13858
rect 14754 13806 14756 13858
rect 14700 13794 14756 13806
rect 14028 13694 14030 13746
rect 14082 13694 14084 13746
rect 14028 13682 14084 13694
rect 16828 13634 16884 13646
rect 16828 13582 16830 13634
rect 16882 13582 16884 13634
rect 16828 13524 16884 13582
rect 17276 13524 17332 13534
rect 16828 13522 17332 13524
rect 16828 13470 17278 13522
rect 17330 13470 17332 13522
rect 16828 13468 17332 13470
rect 17276 13458 17332 13468
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 17500 13076 17556 13916
rect 18284 13970 18340 14364
rect 18284 13918 18286 13970
rect 18338 13918 18340 13970
rect 18284 13906 18340 13918
rect 18396 13972 18452 15150
rect 18508 14530 18564 15260
rect 18508 14478 18510 14530
rect 18562 14478 18564 14530
rect 18508 14466 18564 14478
rect 18732 14420 18788 14430
rect 18732 14326 18788 14364
rect 18620 14308 18676 14318
rect 18620 14214 18676 14252
rect 18396 13906 18452 13916
rect 18844 13972 18900 15260
rect 18956 14754 19012 17724
rect 19068 17444 19124 17454
rect 19068 17350 19124 17388
rect 19180 16772 19236 21420
rect 19516 20188 19572 25340
rect 19628 25330 19684 25340
rect 20188 25396 20244 25406
rect 19628 25172 19684 25182
rect 19628 24724 19684 25116
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 19852 24948 19908 24958
rect 20188 24948 20244 25340
rect 20300 25284 20356 26238
rect 20300 25218 20356 25228
rect 19852 24946 20244 24948
rect 19852 24894 19854 24946
rect 19906 24894 20244 24946
rect 19852 24892 20244 24894
rect 19852 24882 19908 24892
rect 19740 24724 19796 24734
rect 19628 24722 19796 24724
rect 19628 24670 19742 24722
rect 19794 24670 19796 24722
rect 19628 24668 19796 24670
rect 19628 23380 19684 24668
rect 19740 24658 19796 24668
rect 20188 24612 20244 24622
rect 19852 24500 19908 24510
rect 19852 24406 19908 24444
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 19628 23324 19796 23380
rect 19740 23268 19796 23324
rect 19852 23268 19908 23278
rect 19740 23266 19908 23268
rect 19740 23214 19854 23266
rect 19906 23214 19908 23266
rect 19740 23212 19908 23214
rect 19628 23154 19684 23166
rect 19628 23102 19630 23154
rect 19682 23102 19684 23154
rect 19628 22708 19684 23102
rect 19740 23156 19796 23212
rect 19852 23202 19908 23212
rect 19740 23090 19796 23100
rect 19628 22642 19684 22652
rect 20188 22596 20244 24556
rect 20636 24500 20692 26350
rect 20748 24724 20804 24734
rect 20748 24630 20804 24668
rect 20860 24610 20916 26908
rect 22092 26964 22148 26974
rect 22092 26962 23380 26964
rect 22092 26910 22094 26962
rect 22146 26910 23380 26962
rect 22092 26908 23380 26910
rect 22092 26898 22148 26908
rect 23324 26514 23380 26908
rect 23324 26462 23326 26514
rect 23378 26462 23380 26514
rect 23324 26450 23380 26462
rect 21084 26404 21140 26414
rect 21084 26290 21140 26348
rect 22652 26404 22708 26414
rect 23212 26404 23268 26414
rect 22652 26310 22708 26348
rect 23100 26348 23212 26404
rect 21084 26238 21086 26290
rect 21138 26238 21140 26290
rect 21084 26226 21140 26238
rect 22764 26290 22820 26302
rect 22764 26238 22766 26290
rect 22818 26238 22820 26290
rect 22652 26068 22708 26078
rect 22652 25974 22708 26012
rect 21756 25506 21812 25518
rect 21756 25454 21758 25506
rect 21810 25454 21812 25506
rect 21308 25396 21364 25406
rect 21308 25302 21364 25340
rect 21644 24836 21700 24846
rect 20860 24558 20862 24610
rect 20914 24558 20916 24610
rect 20860 24546 20916 24558
rect 20972 24722 21028 24734
rect 20972 24670 20974 24722
rect 21026 24670 21028 24722
rect 20748 24500 20804 24510
rect 20636 24444 20748 24500
rect 20748 24434 20804 24444
rect 20300 23828 20356 23838
rect 20300 23734 20356 23772
rect 20636 23714 20692 23726
rect 20636 23662 20638 23714
rect 20690 23662 20692 23714
rect 20636 23492 20692 23662
rect 20972 23492 21028 24670
rect 21644 24722 21700 24780
rect 21644 24670 21646 24722
rect 21698 24670 21700 24722
rect 21308 24612 21364 24622
rect 21308 24518 21364 24556
rect 21644 23716 21700 24670
rect 21756 24724 21812 25454
rect 22316 25506 22372 25518
rect 22316 25454 22318 25506
rect 22370 25454 22372 25506
rect 22316 24836 22372 25454
rect 22316 24770 22372 24780
rect 22428 25506 22484 25518
rect 22428 25454 22430 25506
rect 22482 25454 22484 25506
rect 21756 23940 21812 24668
rect 22428 24612 22484 25454
rect 22764 24836 22820 26238
rect 23100 24948 23156 26348
rect 23212 26338 23268 26348
rect 23548 26292 23604 26302
rect 23548 26198 23604 26236
rect 23212 26066 23268 26078
rect 23212 26014 23214 26066
rect 23266 26014 23268 26066
rect 23212 25730 23268 26014
rect 23212 25678 23214 25730
rect 23266 25678 23268 25730
rect 23212 25666 23268 25678
rect 23324 25506 23380 25518
rect 23324 25454 23326 25506
rect 23378 25454 23380 25506
rect 23212 24948 23268 24958
rect 23100 24946 23268 24948
rect 23100 24894 23214 24946
rect 23266 24894 23268 24946
rect 23100 24892 23268 24894
rect 23212 24882 23268 24892
rect 22428 24546 22484 24556
rect 22540 24780 22932 24836
rect 22316 24500 22372 24510
rect 21980 24164 22036 24174
rect 21756 23874 21812 23884
rect 21868 23938 21924 23950
rect 21868 23886 21870 23938
rect 21922 23886 21924 23938
rect 21868 23828 21924 23886
rect 21868 23762 21924 23772
rect 21980 23826 22036 24108
rect 21980 23774 21982 23826
rect 22034 23774 22036 23826
rect 21980 23762 22036 23774
rect 22316 23826 22372 24444
rect 22316 23774 22318 23826
rect 22370 23774 22372 23826
rect 21644 23660 21812 23716
rect 20636 23436 21028 23492
rect 20748 23268 20804 23278
rect 20524 23266 20804 23268
rect 20524 23214 20750 23266
rect 20802 23214 20804 23266
rect 20524 23212 20804 23214
rect 19740 22372 19796 22382
rect 19740 22278 19796 22316
rect 19628 22148 19684 22158
rect 19628 21698 19684 22092
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 20188 21812 20244 22540
rect 20412 23154 20468 23166
rect 20412 23102 20414 23154
rect 20466 23102 20468 23154
rect 20412 22372 20468 23102
rect 20412 22306 20468 22316
rect 20524 22484 20580 23212
rect 20748 23202 20804 23212
rect 20860 23044 20916 23436
rect 21644 23268 21700 23278
rect 21644 23174 21700 23212
rect 21532 23044 21588 23054
rect 20860 23042 21588 23044
rect 20860 22990 21534 23042
rect 21586 22990 21588 23042
rect 20860 22988 21588 22990
rect 20188 21746 20244 21756
rect 20300 22258 20356 22270
rect 20300 22206 20302 22258
rect 20354 22206 20356 22258
rect 20300 22148 20356 22206
rect 19628 21646 19630 21698
rect 19682 21646 19684 21698
rect 19628 21634 19684 21646
rect 20076 20804 20132 20814
rect 20076 20710 20132 20748
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 20300 20188 20356 22092
rect 20412 21588 20468 21598
rect 20412 20356 20468 21532
rect 20524 20692 20580 22428
rect 20748 22820 20804 22830
rect 20748 22482 20804 22764
rect 20748 22430 20750 22482
rect 20802 22430 20804 22482
rect 20748 22418 20804 22430
rect 20636 22370 20692 22382
rect 20636 22318 20638 22370
rect 20690 22318 20692 22370
rect 20636 22260 20692 22318
rect 20636 22194 20692 22204
rect 21420 22260 21476 22270
rect 21420 22166 21476 22204
rect 20860 21700 20916 21710
rect 20860 21698 21364 21700
rect 20860 21646 20862 21698
rect 20914 21646 21364 21698
rect 20860 21644 21364 21646
rect 20860 21634 20916 21644
rect 20524 20626 20580 20636
rect 20748 21586 20804 21598
rect 20748 21534 20750 21586
rect 20802 21534 20804 21586
rect 20748 20580 20804 21534
rect 20412 20290 20468 20300
rect 20636 20524 20804 20580
rect 21308 20802 21364 21644
rect 21532 21474 21588 22988
rect 21756 22820 21812 23660
rect 22316 23604 22372 23774
rect 22316 23538 22372 23548
rect 22428 23938 22484 23950
rect 22428 23886 22430 23938
rect 22482 23886 22484 23938
rect 22428 23380 22484 23886
rect 22540 23940 22596 24780
rect 22876 24724 22932 24780
rect 23324 24724 23380 25454
rect 23772 25506 23828 27132
rect 24220 27122 24276 27132
rect 25228 27858 25284 27870
rect 25228 27806 25230 27858
rect 25282 27806 25284 27858
rect 24444 27076 24500 27086
rect 24444 26514 24500 27020
rect 24780 27076 24836 27086
rect 24780 26982 24836 27020
rect 25228 27076 25284 27806
rect 25228 27010 25284 27020
rect 26012 27746 26068 27758
rect 28140 27748 28196 31892
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 26012 27694 26014 27746
rect 26066 27694 26068 27746
rect 24444 26462 24446 26514
rect 24498 26462 24500 26514
rect 24444 26450 24500 26462
rect 25564 26962 25620 26974
rect 25564 26910 25566 26962
rect 25618 26910 25620 26962
rect 25564 26514 25620 26910
rect 25564 26462 25566 26514
rect 25618 26462 25620 26514
rect 25564 26450 25620 26462
rect 25452 26404 25508 26414
rect 25452 26310 25508 26348
rect 23772 25454 23774 25506
rect 23826 25454 23828 25506
rect 23772 25442 23828 25454
rect 24892 26292 24948 26302
rect 24892 25508 24948 26236
rect 25228 26290 25284 26302
rect 25228 26238 25230 26290
rect 25282 26238 25284 26290
rect 25116 25508 25172 25518
rect 24892 25506 25172 25508
rect 24892 25454 25118 25506
rect 25170 25454 25172 25506
rect 24892 25452 25172 25454
rect 25004 25284 25060 25452
rect 25116 25442 25172 25452
rect 25228 25396 25284 26238
rect 25676 26292 25732 26302
rect 25676 26198 25732 26236
rect 25900 26180 25956 26190
rect 25900 26086 25956 26124
rect 25340 26068 25396 26078
rect 25340 25508 25396 26012
rect 26012 25844 26068 27694
rect 28028 27746 28196 27748
rect 28028 27694 28142 27746
rect 28194 27694 28196 27746
rect 28028 27692 28196 27694
rect 27132 27188 27188 27198
rect 26572 26516 26628 26526
rect 26572 26422 26628 26460
rect 27132 26402 27188 27132
rect 27692 27188 27748 27198
rect 27692 27094 27748 27132
rect 27132 26350 27134 26402
rect 27186 26350 27188 26402
rect 27132 26338 27188 26350
rect 27356 27076 27412 27086
rect 26124 26292 26180 26302
rect 26348 26292 26404 26302
rect 26124 26198 26180 26236
rect 26236 26290 26404 26292
rect 26236 26238 26350 26290
rect 26402 26238 26404 26290
rect 26236 26236 26404 26238
rect 25564 25788 26068 25844
rect 25564 25618 25620 25788
rect 26236 25732 26292 26236
rect 26348 26226 26404 26236
rect 26684 26290 26740 26302
rect 26684 26238 26686 26290
rect 26738 26238 26740 26290
rect 25564 25566 25566 25618
rect 25618 25566 25620 25618
rect 25564 25554 25620 25566
rect 25788 25676 26292 25732
rect 26684 26180 26740 26238
rect 27020 26292 27076 26302
rect 27020 26198 27076 26236
rect 25452 25508 25508 25518
rect 25340 25506 25508 25508
rect 25340 25454 25454 25506
rect 25506 25454 25508 25506
rect 25340 25452 25508 25454
rect 25452 25442 25508 25452
rect 25788 25506 25844 25676
rect 25788 25454 25790 25506
rect 25842 25454 25844 25506
rect 25788 25442 25844 25454
rect 26684 25396 26740 26124
rect 25228 25340 25396 25396
rect 25004 25228 25172 25284
rect 25116 25172 25172 25228
rect 25116 25116 25284 25172
rect 22876 24722 23380 24724
rect 22876 24670 22878 24722
rect 22930 24670 23380 24722
rect 22876 24668 23380 24670
rect 22876 24658 22932 24668
rect 22652 24610 22708 24622
rect 22652 24558 22654 24610
rect 22706 24558 22708 24610
rect 22652 24164 22708 24558
rect 23212 24164 23268 24174
rect 22652 24098 22708 24108
rect 22764 24162 23268 24164
rect 22764 24110 23214 24162
rect 23266 24110 23268 24162
rect 22764 24108 23268 24110
rect 22540 23884 22708 23940
rect 22092 23324 22484 23380
rect 22540 23716 22596 23726
rect 22540 23378 22596 23660
rect 22540 23326 22542 23378
rect 22594 23326 22596 23378
rect 21756 22754 21812 22764
rect 21868 23268 21924 23278
rect 21868 22370 21924 23212
rect 21868 22318 21870 22370
rect 21922 22318 21924 22370
rect 21868 22306 21924 22318
rect 21980 23268 22036 23278
rect 22092 23268 22148 23324
rect 22540 23314 22596 23326
rect 21980 23266 22148 23268
rect 21980 23214 21982 23266
rect 22034 23214 22148 23266
rect 21980 23212 22148 23214
rect 21644 22148 21700 22158
rect 21644 22054 21700 22092
rect 21532 21422 21534 21474
rect 21586 21422 21588 21474
rect 21532 21410 21588 21422
rect 21308 20750 21310 20802
rect 21362 20750 21364 20802
rect 19404 20132 19460 20142
rect 19516 20132 19908 20188
rect 20300 20132 20468 20188
rect 19404 20018 19460 20076
rect 19404 19966 19406 20018
rect 19458 19966 19460 20018
rect 19404 19954 19460 19966
rect 19516 19236 19572 19246
rect 19516 19142 19572 19180
rect 19292 19124 19348 19134
rect 19852 19124 19908 20132
rect 19964 20020 20020 20030
rect 19964 19796 20020 19964
rect 19964 19730 20020 19740
rect 19348 19068 19460 19124
rect 19292 19030 19348 19068
rect 19292 18228 19348 18238
rect 19292 17892 19348 18172
rect 19292 17826 19348 17836
rect 19404 17780 19460 19068
rect 19852 19030 19908 19068
rect 20412 19010 20468 20132
rect 20412 18958 20414 19010
rect 20466 18958 20468 19010
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 19628 18676 19684 18686
rect 19628 18582 19684 18620
rect 20188 18338 20244 18350
rect 20188 18286 20190 18338
rect 20242 18286 20244 18338
rect 20188 18116 20244 18286
rect 20188 18050 20244 18060
rect 19516 17780 19572 17790
rect 19404 17778 19572 17780
rect 19404 17726 19518 17778
rect 19570 17726 19572 17778
rect 19404 17724 19572 17726
rect 19516 17714 19572 17724
rect 20412 17668 20468 18958
rect 20524 20132 20580 20142
rect 20524 19348 20580 20076
rect 20636 20020 20692 20524
rect 20636 19954 20692 19964
rect 20748 20356 20804 20366
rect 20524 18562 20580 19292
rect 20748 19234 20804 20300
rect 21308 20188 21364 20750
rect 21868 20804 21924 20814
rect 21420 20692 21476 20702
rect 21420 20598 21476 20636
rect 20748 19182 20750 19234
rect 20802 19182 20804 19234
rect 20748 19170 20804 19182
rect 21084 20132 21364 20188
rect 21532 20468 21588 20478
rect 20524 18510 20526 18562
rect 20578 18510 20580 18562
rect 20524 18498 20580 18510
rect 21084 18452 21140 20132
rect 21308 19348 21364 19358
rect 21308 19234 21364 19292
rect 21308 19182 21310 19234
rect 21362 19182 21364 19234
rect 21308 19170 21364 19182
rect 21420 19236 21476 19246
rect 21084 18386 21140 18396
rect 21196 18788 21252 18798
rect 20748 18228 20804 18238
rect 20748 18134 20804 18172
rect 21084 18228 21140 18238
rect 21196 18228 21252 18732
rect 21420 18450 21476 19180
rect 21420 18398 21422 18450
rect 21474 18398 21476 18450
rect 21420 18386 21476 18398
rect 21532 18450 21588 20412
rect 21868 20130 21924 20748
rect 21868 20078 21870 20130
rect 21922 20078 21924 20130
rect 21980 20188 22036 23212
rect 22204 23154 22260 23166
rect 22204 23102 22206 23154
rect 22258 23102 22260 23154
rect 22204 22482 22260 23102
rect 22540 22708 22596 22718
rect 22204 22430 22206 22482
rect 22258 22430 22260 22482
rect 22204 22418 22260 22430
rect 22428 22652 22540 22708
rect 22092 22260 22148 22270
rect 22092 22258 22372 22260
rect 22092 22206 22094 22258
rect 22146 22206 22372 22258
rect 22092 22204 22372 22206
rect 22092 22194 22148 22204
rect 22204 21700 22260 21710
rect 22204 20802 22260 21644
rect 22204 20750 22206 20802
rect 22258 20750 22260 20802
rect 22204 20468 22260 20750
rect 22204 20402 22260 20412
rect 21980 20122 22036 20132
rect 21868 20020 21924 20078
rect 21868 19954 21924 19964
rect 21756 19796 21812 19806
rect 21756 19346 21812 19740
rect 21756 19294 21758 19346
rect 21810 19294 21812 19346
rect 21756 19282 21812 19294
rect 22316 18788 22372 22204
rect 22428 20188 22484 22652
rect 22540 22642 22596 22652
rect 22540 22370 22596 22382
rect 22540 22318 22542 22370
rect 22594 22318 22596 22370
rect 22540 22260 22596 22318
rect 22540 21924 22596 22204
rect 22652 22258 22708 23884
rect 22764 22596 22820 24108
rect 23212 24098 23268 24108
rect 22876 23940 22932 23950
rect 22876 23846 22932 23884
rect 23100 23826 23156 23838
rect 23100 23774 23102 23826
rect 23154 23774 23156 23826
rect 23100 23716 23156 23774
rect 23212 23828 23268 23838
rect 23212 23734 23268 23772
rect 22876 23660 23156 23716
rect 22876 23154 22932 23660
rect 23212 23604 23268 23614
rect 23100 23268 23156 23278
rect 23100 23174 23156 23212
rect 23212 23266 23268 23548
rect 23996 23380 24052 23390
rect 24220 23380 24276 23390
rect 23212 23214 23214 23266
rect 23266 23214 23268 23266
rect 23212 23202 23268 23214
rect 23324 23266 23380 23278
rect 23324 23214 23326 23266
rect 23378 23214 23380 23266
rect 22876 23102 22878 23154
rect 22930 23102 22932 23154
rect 22876 22820 22932 23102
rect 22988 23156 23044 23166
rect 22988 23062 23044 23100
rect 22876 22754 22932 22764
rect 22988 22708 23044 22718
rect 22764 22540 22932 22596
rect 22652 22206 22654 22258
rect 22706 22206 22708 22258
rect 22652 22194 22708 22206
rect 22540 21868 22820 21924
rect 22652 21588 22708 21598
rect 22652 21494 22708 21532
rect 22540 21476 22596 21486
rect 22540 20802 22596 21420
rect 22764 21028 22820 21868
rect 22876 21140 22932 22540
rect 22988 22370 23044 22652
rect 22988 22318 22990 22370
rect 23042 22318 23044 22370
rect 22988 22306 23044 22318
rect 23324 21924 23380 23214
rect 23996 23266 24052 23324
rect 23996 23214 23998 23266
rect 24050 23214 24052 23266
rect 23996 23202 24052 23214
rect 24108 23324 24220 23380
rect 23548 22484 23604 22494
rect 23548 22370 23604 22428
rect 23548 22318 23550 22370
rect 23602 22318 23604 22370
rect 23548 21924 23604 22318
rect 22988 21868 23380 21924
rect 23436 21868 23604 21924
rect 22988 21252 23044 21868
rect 23436 21700 23492 21868
rect 23324 21644 23492 21700
rect 23772 21700 23828 21710
rect 23212 21586 23268 21598
rect 23212 21534 23214 21586
rect 23266 21534 23268 21586
rect 23212 21476 23268 21534
rect 23212 21410 23268 21420
rect 22988 21196 23156 21252
rect 22876 21084 23044 21140
rect 22764 20972 22932 21028
rect 22540 20750 22542 20802
rect 22594 20750 22596 20802
rect 22540 20738 22596 20750
rect 22764 20690 22820 20702
rect 22764 20638 22766 20690
rect 22818 20638 22820 20690
rect 22764 20188 22820 20638
rect 22428 20132 22708 20188
rect 22652 19348 22708 20132
rect 22764 20122 22820 20132
rect 22876 19458 22932 20972
rect 22876 19406 22878 19458
rect 22930 19406 22932 19458
rect 22876 19394 22932 19406
rect 22764 19348 22820 19358
rect 22652 19346 22820 19348
rect 22652 19294 22766 19346
rect 22818 19294 22820 19346
rect 22652 19292 22820 19294
rect 22764 18900 22820 19292
rect 22988 19236 23044 21084
rect 23100 19796 23156 21196
rect 23100 19730 23156 19740
rect 22988 19170 23044 19180
rect 23212 19122 23268 19134
rect 23212 19070 23214 19122
rect 23266 19070 23268 19122
rect 22764 18844 23044 18900
rect 22316 18732 22932 18788
rect 22316 18674 22372 18732
rect 22316 18622 22318 18674
rect 22370 18622 22372 18674
rect 22316 18610 22372 18622
rect 22876 18674 22932 18732
rect 22876 18622 22878 18674
rect 22930 18622 22932 18674
rect 22764 18564 22820 18574
rect 22764 18470 22820 18508
rect 21532 18398 21534 18450
rect 21586 18398 21588 18450
rect 21532 18386 21588 18398
rect 21980 18452 22036 18462
rect 21980 18358 22036 18396
rect 22652 18340 22708 18350
rect 22652 18246 22708 18284
rect 21084 18226 21252 18228
rect 21084 18174 21086 18226
rect 21138 18174 21252 18226
rect 21084 18172 21252 18174
rect 21084 18162 21140 18172
rect 21644 18116 21700 18126
rect 21532 18060 21644 18116
rect 20524 17668 20580 17678
rect 20412 17666 20580 17668
rect 20412 17614 20526 17666
rect 20578 17614 20580 17666
rect 20412 17612 20580 17614
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 19740 17108 19796 17118
rect 19740 17014 19796 17052
rect 20524 16996 20580 17612
rect 21196 17666 21252 17678
rect 21196 17614 21198 17666
rect 21250 17614 21252 17666
rect 20748 17556 20804 17566
rect 20748 17462 20804 17500
rect 21196 17108 21252 17614
rect 21196 17042 21252 17052
rect 21532 17106 21588 18060
rect 21644 18050 21700 18060
rect 22652 17780 22708 17790
rect 22652 17686 22708 17724
rect 21532 17054 21534 17106
rect 21586 17054 21588 17106
rect 21532 17042 21588 17054
rect 21644 17668 21700 17678
rect 21644 17108 21700 17612
rect 22540 17668 22596 17678
rect 22540 17574 22596 17612
rect 21868 17556 21924 17566
rect 21868 17462 21924 17500
rect 22876 17556 22932 18622
rect 22988 18116 23044 18844
rect 22988 18050 23044 18060
rect 23100 18788 23156 18798
rect 22876 17462 22932 17500
rect 21756 17444 21812 17454
rect 21756 17350 21812 17388
rect 21868 17108 21924 17118
rect 22540 17108 22596 17118
rect 21644 17106 21924 17108
rect 21644 17054 21870 17106
rect 21922 17054 21924 17106
rect 21644 17052 21924 17054
rect 20524 16930 20580 16940
rect 19180 16706 19236 16716
rect 19964 16882 20020 16894
rect 19964 16830 19966 16882
rect 20018 16830 20020 16882
rect 19964 16772 20020 16830
rect 19964 16706 20020 16716
rect 21308 16772 21364 16782
rect 21308 16098 21364 16716
rect 21644 16100 21700 17052
rect 21868 17042 21924 17052
rect 22428 17052 22540 17108
rect 22204 16996 22260 17006
rect 22204 16902 22260 16940
rect 21308 16046 21310 16098
rect 21362 16046 21364 16098
rect 21308 16034 21364 16046
rect 21532 16044 22372 16100
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 21308 15540 21364 15550
rect 21308 15446 21364 15484
rect 21532 15538 21588 16044
rect 21644 15876 21700 15886
rect 21644 15874 21812 15876
rect 21644 15822 21646 15874
rect 21698 15822 21812 15874
rect 21644 15820 21812 15822
rect 21644 15810 21700 15820
rect 21532 15486 21534 15538
rect 21586 15486 21588 15538
rect 21532 15474 21588 15486
rect 21756 15314 21812 15820
rect 22316 15538 22372 16044
rect 22316 15486 22318 15538
rect 22370 15486 22372 15538
rect 22316 15474 22372 15486
rect 22092 15316 22148 15326
rect 22428 15316 22484 17052
rect 22540 17014 22596 17052
rect 22540 15540 22596 15550
rect 22540 15446 22596 15484
rect 21756 15262 21758 15314
rect 21810 15262 21812 15314
rect 21756 15204 21812 15262
rect 21756 15138 21812 15148
rect 21980 15314 22484 15316
rect 21980 15262 22094 15314
rect 22146 15262 22484 15314
rect 21980 15260 22484 15262
rect 22652 15316 22708 15326
rect 18956 14702 18958 14754
rect 19010 14702 19012 14754
rect 18956 14690 19012 14702
rect 21644 15090 21700 15102
rect 21644 15038 21646 15090
rect 21698 15038 21700 15090
rect 21644 14644 21700 15038
rect 20412 14588 21700 14644
rect 19292 14530 19348 14542
rect 19292 14478 19294 14530
rect 19346 14478 19348 14530
rect 19292 14420 19348 14478
rect 20412 14530 20468 14588
rect 20412 14478 20414 14530
rect 20466 14478 20468 14530
rect 20412 14466 20468 14478
rect 21644 14530 21700 14588
rect 21644 14478 21646 14530
rect 21698 14478 21700 14530
rect 21644 14466 21700 14478
rect 19292 14354 19348 14364
rect 20076 14418 20132 14430
rect 20076 14366 20078 14418
rect 20130 14366 20132 14418
rect 20076 14308 20132 14366
rect 20636 14420 20692 14430
rect 20636 14326 20692 14364
rect 21980 14420 22036 15260
rect 22092 15250 22148 15260
rect 22652 15090 22708 15260
rect 23100 15148 23156 18732
rect 23212 15540 23268 19070
rect 23324 18674 23380 21644
rect 23772 21606 23828 21644
rect 23436 21476 23492 21486
rect 23436 21382 23492 21420
rect 23548 20802 23604 20814
rect 23548 20750 23550 20802
rect 23602 20750 23604 20802
rect 23548 20188 23604 20750
rect 24108 20188 24164 23324
rect 24220 23286 24276 23324
rect 25228 23380 25284 25116
rect 25340 23716 25396 25340
rect 26684 25330 26740 25340
rect 27356 24948 27412 27020
rect 28028 26516 28084 27692
rect 28140 27682 28196 27692
rect 28700 27746 28756 27758
rect 28700 27694 28702 27746
rect 28754 27694 28756 27746
rect 28140 27076 28196 27086
rect 28140 26982 28196 27020
rect 28700 27076 28756 27694
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 40012 27186 40068 27198
rect 40012 27134 40014 27186
rect 40066 27134 40068 27186
rect 28700 27010 28756 27020
rect 37660 27076 37716 27086
rect 37660 26982 37716 27020
rect 40012 26964 40068 27134
rect 40012 26898 40068 26908
rect 28028 26450 28084 26460
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 40012 25618 40068 25630
rect 40012 25566 40014 25618
rect 40066 25566 40068 25618
rect 29260 25508 29316 25518
rect 29260 25394 29316 25452
rect 30604 25508 30660 25518
rect 29260 25342 29262 25394
rect 29314 25342 29316 25394
rect 29260 25330 29316 25342
rect 29372 25396 29428 25406
rect 29036 25282 29092 25294
rect 29036 25230 29038 25282
rect 29090 25230 29092 25282
rect 27356 24946 27748 24948
rect 27356 24894 27358 24946
rect 27410 24894 27748 24946
rect 27356 24892 27748 24894
rect 27356 24882 27412 24892
rect 25340 23650 25396 23660
rect 27692 24722 27748 24892
rect 27692 24670 27694 24722
rect 27746 24670 27748 24722
rect 26124 23380 26180 23390
rect 25228 23378 26180 23380
rect 25228 23326 25230 23378
rect 25282 23326 26126 23378
rect 26178 23326 26180 23378
rect 25228 23324 26180 23326
rect 25228 23314 25284 23324
rect 26124 23314 26180 23324
rect 26236 23380 26292 23390
rect 25452 23154 25508 23166
rect 25452 23102 25454 23154
rect 25506 23102 25508 23154
rect 24332 23044 24388 23054
rect 24332 22950 24388 22988
rect 25452 23044 25508 23102
rect 25452 22978 25508 22988
rect 26012 23042 26068 23054
rect 26012 22990 26014 23042
rect 26066 22990 26068 23042
rect 25900 22932 25956 22942
rect 25564 22930 25956 22932
rect 25564 22878 25902 22930
rect 25954 22878 25956 22930
rect 25564 22876 25956 22878
rect 24220 22596 24276 22606
rect 24220 22482 24276 22540
rect 24220 22430 24222 22482
rect 24274 22430 24276 22482
rect 24220 22418 24276 22430
rect 25340 22484 25396 22494
rect 24668 22370 24724 22382
rect 24668 22318 24670 22370
rect 24722 22318 24724 22370
rect 24556 22258 24612 22270
rect 24556 22206 24558 22258
rect 24610 22206 24612 22258
rect 23436 20132 23604 20188
rect 23772 20132 24164 20188
rect 24444 21588 24500 21598
rect 23436 20020 23492 20132
rect 23436 19954 23492 19964
rect 23324 18622 23326 18674
rect 23378 18622 23380 18674
rect 23324 18610 23380 18622
rect 23660 18900 23716 18910
rect 23660 18674 23716 18844
rect 23660 18622 23662 18674
rect 23714 18622 23716 18674
rect 23660 18610 23716 18622
rect 23548 18452 23604 18462
rect 23436 18340 23492 18350
rect 23436 17666 23492 18284
rect 23436 17614 23438 17666
rect 23490 17614 23492 17666
rect 23436 17602 23492 17614
rect 23212 15474 23268 15484
rect 22652 15038 22654 15090
rect 22706 15038 22708 15090
rect 22652 15026 22708 15038
rect 22876 15092 23156 15148
rect 22092 14588 22484 14644
rect 22092 14530 22148 14588
rect 22092 14478 22094 14530
rect 22146 14478 22148 14530
rect 22092 14466 22148 14478
rect 22428 14532 22484 14588
rect 22540 14532 22596 14542
rect 22428 14530 22596 14532
rect 22428 14478 22542 14530
rect 22594 14478 22596 14530
rect 22428 14476 22596 14478
rect 22540 14466 22596 14476
rect 22876 14530 22932 15092
rect 22876 14478 22878 14530
rect 22930 14478 22932 14530
rect 22876 14466 22932 14478
rect 21980 14354 22036 14364
rect 22316 14420 22372 14430
rect 22316 14326 22372 14364
rect 23548 14420 23604 18396
rect 23772 18004 23828 20132
rect 23884 19234 23940 19246
rect 23884 19182 23886 19234
rect 23938 19182 23940 19234
rect 23884 18340 23940 19182
rect 24444 19234 24500 21532
rect 24556 20020 24612 22206
rect 24556 19348 24612 19964
rect 24556 19282 24612 19292
rect 24668 19908 24724 22318
rect 25340 22370 25396 22428
rect 25340 22318 25342 22370
rect 25394 22318 25396 22370
rect 25340 22306 25396 22318
rect 25564 21810 25620 22876
rect 25900 22866 25956 22876
rect 26012 22482 26068 22990
rect 26012 22430 26014 22482
rect 26066 22430 26068 22482
rect 26012 22418 26068 22430
rect 25564 21758 25566 21810
rect 25618 21758 25620 21810
rect 25564 21746 25620 21758
rect 25676 21812 25732 21822
rect 25676 21718 25732 21756
rect 26236 21810 26292 23324
rect 26908 23268 26964 23278
rect 26908 23174 26964 23212
rect 26572 23154 26628 23166
rect 26572 23102 26574 23154
rect 26626 23102 26628 23154
rect 26572 23044 26628 23102
rect 26572 22978 26628 22988
rect 27692 22484 27748 24670
rect 28476 24612 28532 24622
rect 28476 24518 28532 24556
rect 29036 23938 29092 25230
rect 29372 24836 29428 25340
rect 29036 23886 29038 23938
rect 29090 23886 29092 23938
rect 29036 23874 29092 23886
rect 29148 24780 29428 24836
rect 28476 23378 28532 23390
rect 28476 23326 28478 23378
rect 28530 23326 28532 23378
rect 28140 23156 28196 23166
rect 28140 23062 28196 23100
rect 26236 21758 26238 21810
rect 26290 21758 26292 21810
rect 26236 21746 26292 21758
rect 27580 22428 27692 22484
rect 27580 21812 27636 22428
rect 27692 22418 27748 22428
rect 28140 22596 28196 22606
rect 28140 22482 28196 22540
rect 28140 22430 28142 22482
rect 28194 22430 28196 22482
rect 28140 21812 28196 22430
rect 27580 21810 27972 21812
rect 27580 21758 27582 21810
rect 27634 21758 27972 21810
rect 27580 21756 27972 21758
rect 27580 21746 27636 21756
rect 26572 21700 26628 21710
rect 26572 21606 26628 21644
rect 25228 21588 25284 21598
rect 25452 21588 25508 21598
rect 25228 21494 25284 21532
rect 25340 21586 25508 21588
rect 25340 21534 25454 21586
rect 25506 21534 25508 21586
rect 25340 21532 25508 21534
rect 25340 20244 25396 21532
rect 25452 21522 25508 21532
rect 25788 21586 25844 21598
rect 25788 21534 25790 21586
rect 25842 21534 25844 21586
rect 25788 21476 25844 21534
rect 25788 21410 25844 21420
rect 27916 21586 27972 21756
rect 28140 21746 28196 21756
rect 28364 22594 28420 22606
rect 28364 22542 28366 22594
rect 28418 22542 28420 22594
rect 27916 21534 27918 21586
rect 27970 21534 27972 21586
rect 25228 20188 25396 20244
rect 27916 20914 27972 21534
rect 27916 20862 27918 20914
rect 27970 20862 27972 20914
rect 24444 19182 24446 19234
rect 24498 19182 24500 19234
rect 24444 19170 24500 19182
rect 24668 19124 24724 19852
rect 25116 20132 25284 20188
rect 25116 19796 25172 20132
rect 25452 20130 25508 20142
rect 25452 20078 25454 20130
rect 25506 20078 25508 20130
rect 25228 20020 25284 20030
rect 25228 19926 25284 19964
rect 24556 19068 24724 19124
rect 24892 19740 25116 19796
rect 24332 19010 24388 19022
rect 24332 18958 24334 19010
rect 24386 18958 24388 19010
rect 24332 18900 24388 18958
rect 24556 19010 24612 19068
rect 24556 18958 24558 19010
rect 24610 18958 24612 19010
rect 24556 18946 24612 18958
rect 24332 18834 24388 18844
rect 24444 18788 24500 18798
rect 24108 18676 24164 18686
rect 23996 18564 24052 18574
rect 23996 18470 24052 18508
rect 24108 18450 24164 18620
rect 24444 18564 24500 18732
rect 24108 18398 24110 18450
rect 24162 18398 24164 18450
rect 24108 18386 24164 18398
rect 24220 18508 24500 18564
rect 24220 18450 24276 18508
rect 24220 18398 24222 18450
rect 24274 18398 24276 18450
rect 24220 18386 24276 18398
rect 24668 18452 24724 18462
rect 24892 18452 24948 19740
rect 25116 19730 25172 19740
rect 25004 19012 25060 19022
rect 25452 19012 25508 20078
rect 26684 20132 26740 20142
rect 26684 20038 26740 20076
rect 25676 20018 25732 20030
rect 25676 19966 25678 20018
rect 25730 19966 25732 20018
rect 25676 19348 25732 19966
rect 25900 20018 25956 20030
rect 25900 19966 25902 20018
rect 25954 19966 25956 20018
rect 25900 19460 25956 19966
rect 26236 20018 26292 20030
rect 26236 19966 26238 20018
rect 26290 19966 26292 20018
rect 26012 19908 26068 19918
rect 26236 19908 26292 19966
rect 26908 20020 26964 20030
rect 26908 19926 26964 19964
rect 27916 20018 27972 20862
rect 27916 19966 27918 20018
rect 27970 19966 27972 20018
rect 26012 19906 26292 19908
rect 26012 19854 26014 19906
rect 26066 19854 26292 19906
rect 26012 19852 26292 19854
rect 26460 19906 26516 19918
rect 26460 19854 26462 19906
rect 26514 19854 26516 19906
rect 26012 19842 26068 19852
rect 25900 19404 26068 19460
rect 25676 19282 25732 19292
rect 25060 18956 25508 19012
rect 25788 19236 25844 19246
rect 25004 18918 25060 18956
rect 24668 18450 24948 18452
rect 24668 18398 24670 18450
rect 24722 18398 24948 18450
rect 24668 18396 24948 18398
rect 25676 18452 25732 18462
rect 24668 18386 24724 18396
rect 23884 18274 23940 18284
rect 23772 17948 24276 18004
rect 23548 14354 23604 14364
rect 23660 17780 23716 17790
rect 20076 14242 20132 14252
rect 20188 14306 20244 14318
rect 20188 14254 20190 14306
rect 20242 14254 20244 14306
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 19516 13972 19572 13982
rect 20076 13972 20132 13982
rect 18844 13970 19796 13972
rect 18844 13918 18846 13970
rect 18898 13918 19518 13970
rect 19570 13918 19796 13970
rect 18844 13916 19796 13918
rect 18844 13906 18900 13916
rect 19516 13906 19572 13916
rect 19740 13858 19796 13916
rect 20076 13878 20132 13916
rect 19740 13806 19742 13858
rect 19794 13806 19796 13858
rect 19740 13794 19796 13806
rect 19852 13860 19908 13870
rect 19852 13766 19908 13804
rect 17948 13636 18004 13646
rect 18172 13636 18228 13646
rect 17948 13634 18228 13636
rect 17948 13582 17950 13634
rect 18002 13582 18174 13634
rect 18226 13582 18228 13634
rect 17948 13580 18228 13582
rect 17948 13570 18004 13580
rect 17612 13076 17668 13086
rect 17500 13074 17892 13076
rect 17500 13022 17614 13074
rect 17666 13022 17892 13074
rect 17500 13020 17892 13022
rect 17612 13010 17668 13020
rect 17836 12962 17892 13020
rect 17836 12910 17838 12962
rect 17890 12910 17892 12962
rect 17836 12898 17892 12910
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 18060 3554 18116 13580
rect 18172 13570 18228 13580
rect 18620 13524 18676 13534
rect 18620 13074 18676 13468
rect 20188 13524 20244 14254
rect 21084 14308 21140 14318
rect 20748 13860 20804 13870
rect 20412 13748 20468 13758
rect 20412 13654 20468 13692
rect 20188 13458 20244 13468
rect 18620 13022 18622 13074
rect 18674 13022 18676 13074
rect 18620 13010 18676 13022
rect 20748 13074 20804 13804
rect 21084 13858 21140 14252
rect 21868 14308 21924 14318
rect 21868 14214 21924 14252
rect 22764 14306 22820 14318
rect 22764 14254 22766 14306
rect 22818 14254 22820 14306
rect 21084 13806 21086 13858
rect 21138 13806 21140 13858
rect 21084 13794 21140 13806
rect 20748 13022 20750 13074
rect 20802 13022 20804 13074
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 18060 3502 18062 3554
rect 18114 3502 18116 3554
rect 18060 3490 18116 3502
rect 18620 3666 18676 3678
rect 18620 3614 18622 3666
rect 18674 3614 18676 3666
rect 18620 3388 18676 3614
rect 20748 3554 20804 13022
rect 22652 13748 22708 13758
rect 22652 12962 22708 13692
rect 22764 13636 22820 14254
rect 23436 14308 23492 14318
rect 23436 13748 23492 14252
rect 23436 13682 23492 13692
rect 23660 13746 23716 17724
rect 23884 17666 23940 17678
rect 23884 17614 23886 17666
rect 23938 17614 23940 17666
rect 23884 17108 23940 17614
rect 24220 17666 24276 17948
rect 24220 17614 24222 17666
rect 24274 17614 24276 17666
rect 24220 17602 24276 17614
rect 24444 17556 24500 17566
rect 24444 17462 24500 17500
rect 23884 17042 23940 17052
rect 24220 17444 24276 17454
rect 24220 16994 24276 17388
rect 24556 17444 24612 17454
rect 24556 17350 24612 17388
rect 25452 17444 25508 17454
rect 24332 17108 24388 17118
rect 24332 17014 24388 17052
rect 24220 16942 24222 16994
rect 24274 16942 24276 16994
rect 24220 16930 24276 16942
rect 25452 16996 25508 17388
rect 24556 16884 24612 16894
rect 25116 16884 25172 16894
rect 25340 16884 25396 16894
rect 24556 16882 25172 16884
rect 24556 16830 24558 16882
rect 24610 16830 25118 16882
rect 25170 16830 25172 16882
rect 24556 16828 25172 16830
rect 24556 16818 24612 16828
rect 25116 16818 25172 16828
rect 25228 16882 25396 16884
rect 25228 16830 25342 16882
rect 25394 16830 25396 16882
rect 25228 16828 25396 16830
rect 25228 16660 25284 16828
rect 25340 16818 25396 16828
rect 25452 16882 25508 16940
rect 25452 16830 25454 16882
rect 25506 16830 25508 16882
rect 25452 16818 25508 16830
rect 25676 16882 25732 18396
rect 25676 16830 25678 16882
rect 25730 16830 25732 16882
rect 25676 16818 25732 16830
rect 24892 16604 25284 16660
rect 24892 16210 24948 16604
rect 24892 16158 24894 16210
rect 24946 16158 24948 16210
rect 24892 16146 24948 16158
rect 24220 16098 24276 16110
rect 24220 16046 24222 16098
rect 24274 16046 24276 16098
rect 23660 13694 23662 13746
rect 23714 13694 23716 13746
rect 23660 13682 23716 13694
rect 23884 14420 23940 14430
rect 23884 13746 23940 14364
rect 24220 14308 24276 16046
rect 25788 15876 25844 19180
rect 26012 18900 26068 19404
rect 26460 19346 26516 19854
rect 26460 19294 26462 19346
rect 26514 19294 26516 19346
rect 26460 19282 26516 19294
rect 27580 19908 27636 19918
rect 27916 19908 27972 19966
rect 27580 19906 27972 19908
rect 27580 19854 27582 19906
rect 27634 19854 27972 19906
rect 27580 19852 27972 19854
rect 28364 20020 28420 22542
rect 28476 21700 28532 23326
rect 28700 23268 28756 23278
rect 28588 23156 28644 23166
rect 28588 23062 28644 23100
rect 28700 23154 28756 23212
rect 28700 23102 28702 23154
rect 28754 23102 28756 23154
rect 28700 22594 28756 23102
rect 28700 22542 28702 22594
rect 28754 22542 28756 22594
rect 28700 22530 28756 22542
rect 28588 22484 28644 22494
rect 28588 22390 28644 22428
rect 29148 22146 29204 24780
rect 29260 24612 29316 24622
rect 29260 24050 29316 24556
rect 30604 24610 30660 25452
rect 37660 25508 37716 25518
rect 37660 25414 37716 25452
rect 40012 24948 40068 25566
rect 40012 24882 40068 24892
rect 30604 24558 30606 24610
rect 30658 24558 30660 24610
rect 30604 24546 30660 24558
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 29260 23998 29262 24050
rect 29314 23998 29316 24050
rect 29260 23986 29316 23998
rect 29484 23940 29540 23950
rect 29484 23846 29540 23884
rect 29596 23938 29652 23950
rect 29596 23886 29598 23938
rect 29650 23886 29652 23938
rect 29596 23268 29652 23886
rect 29596 23202 29652 23212
rect 29932 23156 29988 23166
rect 29932 22594 29988 23100
rect 29932 22542 29934 22594
rect 29986 22542 29988 22594
rect 29932 22530 29988 22542
rect 30828 23156 30884 23166
rect 29148 22094 29150 22146
rect 29202 22094 29204 22146
rect 28700 21700 28756 21710
rect 28476 21698 28756 21700
rect 28476 21646 28702 21698
rect 28754 21646 28756 21698
rect 28476 21644 28756 21646
rect 28700 21634 28756 21644
rect 29148 20804 29204 22094
rect 29372 22370 29428 22382
rect 29372 22318 29374 22370
rect 29426 22318 29428 22370
rect 29372 22260 29428 22318
rect 29820 22260 29876 22270
rect 29372 22258 29876 22260
rect 29372 22206 29822 22258
rect 29874 22206 29876 22258
rect 29372 22204 29876 22206
rect 29372 21476 29428 22204
rect 29820 22194 29876 22204
rect 29932 22260 29988 22270
rect 29932 22166 29988 22204
rect 30828 22260 30884 23100
rect 37660 23156 37716 23166
rect 37660 23062 37716 23100
rect 40012 22932 40068 22942
rect 40012 22838 40068 22876
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 40012 22482 40068 22494
rect 40012 22430 40014 22482
rect 40066 22430 40068 22482
rect 37660 22372 37716 22382
rect 37660 22278 37716 22316
rect 29372 21410 29428 21420
rect 30828 21474 30884 22204
rect 40012 22260 40068 22430
rect 40012 22194 40068 22204
rect 30828 21422 30830 21474
rect 30882 21422 30884 21474
rect 30828 21410 30884 21422
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 40012 20914 40068 20926
rect 40012 20862 40014 20914
rect 40066 20862 40068 20914
rect 29372 20804 29428 20814
rect 29148 20802 29428 20804
rect 29148 20750 29374 20802
rect 29426 20750 29428 20802
rect 29148 20748 29428 20750
rect 29372 20738 29428 20748
rect 37660 20804 37716 20814
rect 37660 20710 37716 20748
rect 27580 19236 27636 19852
rect 27580 19170 27636 19180
rect 28364 19236 28420 19964
rect 29036 20578 29092 20590
rect 29036 20526 29038 20578
rect 29090 20526 29092 20578
rect 28700 19906 28756 19918
rect 28700 19854 28702 19906
rect 28754 19854 28756 19906
rect 28588 19348 28644 19358
rect 28588 19254 28644 19292
rect 28364 19170 28420 19180
rect 28700 19012 28756 19854
rect 29036 19234 29092 20526
rect 29260 20580 29316 20590
rect 29260 20486 29316 20524
rect 30828 20580 30884 20590
rect 30828 19906 30884 20524
rect 40012 20244 40068 20862
rect 40012 20178 40068 20188
rect 30828 19854 30830 19906
rect 30882 19854 30884 19906
rect 30828 19842 30884 19854
rect 37660 20018 37716 20030
rect 37660 19966 37662 20018
rect 37714 19966 37716 20018
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 37660 19348 37716 19966
rect 40012 19794 40068 19806
rect 40012 19742 40014 19794
rect 40066 19742 40068 19794
rect 40012 19572 40068 19742
rect 40012 19506 40068 19516
rect 37660 19282 37716 19292
rect 29036 19182 29038 19234
rect 29090 19182 29092 19234
rect 29036 19170 29092 19182
rect 29372 19234 29428 19246
rect 29372 19182 29374 19234
rect 29426 19182 29428 19234
rect 29260 19012 29316 19022
rect 28700 19010 29316 19012
rect 28700 18958 29262 19010
rect 29314 18958 29316 19010
rect 28700 18956 29316 18958
rect 29260 18946 29316 18956
rect 26012 16772 26068 18844
rect 29372 18676 29428 19182
rect 29596 19236 29652 19246
rect 29596 19142 29652 19180
rect 29372 18610 29428 18620
rect 28812 18338 28868 18350
rect 28812 18286 28814 18338
rect 28866 18286 28868 18338
rect 27020 17668 27076 17678
rect 27020 17108 27076 17612
rect 26684 16996 26740 17006
rect 26684 16902 26740 16940
rect 26012 16706 26068 16716
rect 26236 16882 26292 16894
rect 26236 16830 26238 16882
rect 26290 16830 26292 16882
rect 26124 15876 26180 15886
rect 25788 15820 26124 15876
rect 25452 15540 25508 15550
rect 25452 15538 25956 15540
rect 25452 15486 25454 15538
rect 25506 15486 25956 15538
rect 25452 15484 25956 15486
rect 25452 15474 25508 15484
rect 25228 15316 25284 15326
rect 25228 15222 25284 15260
rect 25452 15316 25508 15326
rect 25452 15148 25508 15260
rect 24220 14242 24276 14252
rect 25228 15092 25508 15148
rect 25564 15314 25620 15326
rect 25564 15262 25566 15314
rect 25618 15262 25620 15314
rect 25228 13858 25284 15092
rect 25340 14530 25396 14542
rect 25340 14478 25342 14530
rect 25394 14478 25396 14530
rect 25340 14308 25396 14478
rect 25564 14532 25620 15262
rect 25788 15316 25844 15326
rect 25788 15222 25844 15260
rect 25900 14644 25956 15484
rect 26124 15314 26180 15820
rect 26124 15262 26126 15314
rect 26178 15262 26180 15314
rect 26124 15148 26180 15262
rect 26236 15316 26292 16830
rect 26460 16882 26516 16894
rect 26460 16830 26462 16882
rect 26514 16830 26516 16882
rect 26460 16324 26516 16830
rect 26460 16258 26516 16268
rect 26572 16770 26628 16782
rect 26572 16718 26574 16770
rect 26626 16718 26628 16770
rect 26572 15428 26628 16718
rect 27020 16210 27076 17052
rect 27020 16158 27022 16210
rect 27074 16158 27076 16210
rect 27020 16146 27076 16158
rect 27356 16772 27412 16782
rect 27356 15986 27412 16716
rect 27468 16324 27524 16334
rect 27468 16230 27524 16268
rect 27356 15934 27358 15986
rect 27410 15934 27412 15986
rect 26908 15428 26964 15438
rect 26572 15426 26964 15428
rect 26572 15374 26910 15426
rect 26962 15374 26964 15426
rect 26572 15372 26964 15374
rect 26908 15362 26964 15372
rect 26236 15250 26292 15260
rect 26124 15092 26292 15148
rect 26124 14644 26180 14654
rect 25900 14642 26180 14644
rect 25900 14590 26126 14642
rect 26178 14590 26180 14642
rect 25900 14588 26180 14590
rect 26124 14578 26180 14588
rect 25564 14466 25620 14476
rect 26236 14308 26292 15092
rect 26908 14644 26964 14654
rect 25396 14252 26292 14308
rect 26684 14532 26740 14542
rect 25340 14242 25396 14252
rect 25228 13806 25230 13858
rect 25282 13806 25284 13858
rect 25228 13794 25284 13806
rect 23884 13694 23886 13746
rect 23938 13694 23940 13746
rect 23884 13682 23940 13694
rect 24108 13748 24164 13758
rect 24108 13654 24164 13692
rect 25340 13748 25396 13758
rect 25340 13654 25396 13692
rect 25564 13746 25620 13758
rect 25564 13694 25566 13746
rect 25618 13694 25620 13746
rect 23212 13636 23268 13646
rect 22764 13634 23268 13636
rect 22764 13582 23214 13634
rect 23266 13582 23268 13634
rect 22764 13580 23268 13582
rect 22652 12910 22654 12962
rect 22706 12910 22708 12962
rect 22652 12898 22708 12910
rect 20748 3502 20750 3554
rect 20802 3502 20804 3554
rect 20748 3490 20804 3502
rect 22876 3668 22932 3678
rect 18172 3332 18676 3388
rect 20188 3444 20244 3454
rect 18172 800 18228 3332
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 20188 800 20244 3388
rect 21756 3444 21812 3454
rect 21756 3330 21812 3388
rect 21756 3278 21758 3330
rect 21810 3278 21812 3330
rect 21756 3266 21812 3278
rect 22876 800 22932 3612
rect 23212 3556 23268 13580
rect 23548 13524 23604 13534
rect 23436 13522 23604 13524
rect 23436 13470 23550 13522
rect 23602 13470 23604 13522
rect 23436 13468 23604 13470
rect 23436 13074 23492 13468
rect 23548 13458 23604 13468
rect 23436 13022 23438 13074
rect 23490 13022 23492 13074
rect 23436 13010 23492 13022
rect 25564 13074 25620 13694
rect 25564 13022 25566 13074
rect 25618 13022 25620 13074
rect 25564 4338 25620 13022
rect 26124 13074 26180 14252
rect 26684 13970 26740 14476
rect 26684 13918 26686 13970
rect 26738 13918 26740 13970
rect 26684 13906 26740 13918
rect 26908 13970 26964 14588
rect 26908 13918 26910 13970
rect 26962 13918 26964 13970
rect 26908 13906 26964 13918
rect 27020 13860 27076 13870
rect 27356 13860 27412 15934
rect 27468 15874 27524 15886
rect 27468 15822 27470 15874
rect 27522 15822 27524 15874
rect 27468 15204 27524 15822
rect 28028 15876 28084 15886
rect 28028 15782 28084 15820
rect 28812 15876 28868 18286
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 40012 17778 40068 17790
rect 40012 17726 40014 17778
rect 40066 17726 40068 17778
rect 37660 17668 37716 17678
rect 37660 17574 37716 17612
rect 37884 16882 37940 16894
rect 37884 16830 37886 16882
rect 37938 16830 37940 16882
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 28812 15810 28868 15820
rect 29260 15876 29316 15886
rect 29260 15540 29316 15820
rect 29484 15540 29540 15550
rect 29260 15538 29540 15540
rect 29260 15486 29486 15538
rect 29538 15486 29540 15538
rect 29260 15484 29540 15486
rect 27468 15138 27524 15148
rect 29036 15204 29092 15214
rect 29036 15110 29092 15148
rect 28252 14644 28308 14654
rect 28252 14550 28308 14588
rect 29260 14642 29316 15484
rect 29484 15474 29540 15484
rect 37660 15314 37716 15326
rect 37660 15262 37662 15314
rect 37714 15262 37716 15314
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 29260 14590 29262 14642
rect 29314 14590 29316 14642
rect 29260 14578 29316 14590
rect 37660 14644 37716 15262
rect 37884 15204 37940 16830
rect 40012 16884 40068 17726
rect 40012 16818 40068 16828
rect 40012 16658 40068 16670
rect 40012 16606 40014 16658
rect 40066 16606 40068 16658
rect 40012 16212 40068 16606
rect 40012 16146 40068 16156
rect 37884 15138 37940 15148
rect 40012 15202 40068 15214
rect 40012 15150 40014 15202
rect 40066 15150 40068 15202
rect 40012 14868 40068 15150
rect 40012 14802 40068 14812
rect 37660 14578 37716 14588
rect 27020 13858 27412 13860
rect 27020 13806 27022 13858
rect 27074 13806 27412 13858
rect 27020 13804 27412 13806
rect 27020 13794 27076 13804
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 26124 13022 26126 13074
rect 26178 13022 26180 13074
rect 26124 13010 26180 13022
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 40236 9154 40292 9166
rect 40236 9102 40238 9154
rect 40290 9102 40292 9154
rect 40236 8820 40292 9102
rect 40236 8754 40292 8764
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 25564 4286 25566 4338
rect 25618 4286 25620 4338
rect 25564 4274 25620 4286
rect 24892 4116 24948 4126
rect 23212 3490 23268 3500
rect 24556 3556 24612 3566
rect 24556 3462 24612 3500
rect 24892 800 24948 4060
rect 26236 4116 26292 4126
rect 26236 4022 26292 4060
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 25564 3668 25620 3678
rect 25564 3574 25620 3612
rect 18144 0 18256 800
rect 20160 0 20272 800
rect 22848 0 22960 800
rect 24864 0 24976 800
<< via2 >>
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 17500 38220 17556 38276
rect 18620 38274 18676 38276
rect 18620 38222 18622 38274
rect 18622 38222 18674 38274
rect 18674 38222 18676 38274
rect 18620 38220 18676 38222
rect 20860 38220 20916 38276
rect 22092 38274 22148 38276
rect 22092 38222 22094 38274
rect 22094 38222 22146 38274
rect 22146 38222 22148 38274
rect 22092 38220 22148 38222
rect 23548 38220 23604 38276
rect 25564 38274 25620 38276
rect 25564 38222 25566 38274
rect 25566 38222 25618 38274
rect 25618 38222 25620 38274
rect 25564 38220 25620 38222
rect 16828 37436 16884 37492
rect 16156 36652 16212 36708
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 13916 27858 13972 27860
rect 13916 27806 13918 27858
rect 13918 27806 13970 27858
rect 13970 27806 13972 27858
rect 13916 27804 13972 27806
rect 14364 27804 14420 27860
rect 10892 27580 10948 27636
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 4284 24722 4340 24724
rect 4284 24670 4286 24722
rect 4286 24670 4338 24722
rect 4338 24670 4340 24722
rect 4284 24668 4340 24670
rect 1932 24498 1988 24500
rect 1932 24446 1934 24498
rect 1934 24446 1986 24498
rect 1986 24446 1988 24498
rect 1932 24444 1988 24446
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 9996 24050 10052 24052
rect 9996 23998 9998 24050
rect 9998 23998 10050 24050
rect 10050 23998 10052 24050
rect 9996 23996 10052 23998
rect 4284 23938 4340 23940
rect 4284 23886 4286 23938
rect 4286 23886 4338 23938
rect 4338 23886 4340 23938
rect 4284 23884 4340 23886
rect 1932 23548 1988 23604
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 4284 21586 4340 21588
rect 4284 21534 4286 21586
rect 4286 21534 4338 21586
rect 4338 21534 4340 21586
rect 4284 21532 4340 21534
rect 9884 21532 9940 21588
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 1932 20860 1988 20916
rect 9884 20636 9940 20692
rect 12908 27020 12964 27076
rect 12796 23996 12852 24052
rect 12124 23826 12180 23828
rect 12124 23774 12126 23826
rect 12126 23774 12178 23826
rect 12178 23774 12180 23826
rect 12124 23772 12180 23774
rect 14700 27746 14756 27748
rect 14700 27694 14702 27746
rect 14702 27694 14754 27746
rect 14754 27694 14756 27746
rect 14700 27692 14756 27694
rect 16268 28530 16324 28532
rect 16268 28478 16270 28530
rect 16270 28478 16322 28530
rect 16322 28478 16324 28530
rect 16268 28476 16324 28478
rect 16940 28530 16996 28532
rect 16940 28478 16942 28530
rect 16942 28478 16994 28530
rect 16994 28478 16996 28530
rect 16940 28476 16996 28478
rect 16156 27244 16212 27300
rect 16380 27804 16436 27860
rect 14364 27074 14420 27076
rect 14364 27022 14366 27074
rect 14366 27022 14418 27074
rect 14418 27022 14420 27074
rect 14364 27020 14420 27022
rect 15036 26962 15092 26964
rect 15036 26910 15038 26962
rect 15038 26910 15090 26962
rect 15090 26910 15092 26962
rect 15036 26908 15092 26910
rect 16828 27580 16884 27636
rect 17388 36706 17444 36708
rect 17388 36654 17390 36706
rect 17390 36654 17442 36706
rect 17442 36654 17444 36706
rect 17388 36652 17444 36654
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 18396 37490 18452 37492
rect 18396 37438 18398 37490
rect 18398 37438 18450 37490
rect 18450 37438 18452 37490
rect 18396 37436 18452 37438
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 17500 27746 17556 27748
rect 17500 27694 17502 27746
rect 17502 27694 17554 27746
rect 17554 27694 17556 27746
rect 17500 27692 17556 27694
rect 17388 27244 17444 27300
rect 16492 27020 16548 27076
rect 13020 24610 13076 24612
rect 13020 24558 13022 24610
rect 13022 24558 13074 24610
rect 13074 24558 13076 24610
rect 13020 24556 13076 24558
rect 16156 24556 16212 24612
rect 13804 23996 13860 24052
rect 13020 23548 13076 23604
rect 13580 23826 13636 23828
rect 13580 23774 13582 23826
rect 13582 23774 13634 23826
rect 13634 23774 13636 23826
rect 13580 23772 13636 23774
rect 13468 23548 13524 23604
rect 13916 23436 13972 23492
rect 12684 23154 12740 23156
rect 12684 23102 12686 23154
rect 12686 23102 12738 23154
rect 12738 23102 12740 23154
rect 12684 23100 12740 23102
rect 14140 23548 14196 23604
rect 11564 22204 11620 22260
rect 15148 23938 15204 23940
rect 15148 23886 15150 23938
rect 15150 23886 15202 23938
rect 15202 23886 15204 23938
rect 15148 23884 15204 23886
rect 14924 23436 14980 23492
rect 15596 23772 15652 23828
rect 14140 23100 14196 23156
rect 13580 22258 13636 22260
rect 13580 22206 13582 22258
rect 13582 22206 13634 22258
rect 13634 22206 13636 22258
rect 13580 22204 13636 22206
rect 15932 23826 15988 23828
rect 15932 23774 15934 23826
rect 15934 23774 15986 23826
rect 15986 23774 15988 23826
rect 15932 23772 15988 23774
rect 15932 23436 15988 23492
rect 16044 23324 16100 23380
rect 15820 23100 15876 23156
rect 11452 21586 11508 21588
rect 11452 21534 11454 21586
rect 11454 21534 11506 21586
rect 11506 21534 11508 21586
rect 11452 21532 11508 21534
rect 13468 21532 13524 21588
rect 12124 20860 12180 20916
rect 12796 20860 12852 20916
rect 13356 20860 13412 20916
rect 13468 20690 13524 20692
rect 13468 20638 13470 20690
rect 13470 20638 13522 20690
rect 13522 20638 13524 20690
rect 13468 20636 13524 20638
rect 10892 20076 10948 20132
rect 4284 20018 4340 20020
rect 4284 19966 4286 20018
rect 4286 19966 4338 20018
rect 4338 19966 4340 20018
rect 4284 19964 4340 19966
rect 9884 19964 9940 20020
rect 1932 19794 1988 19796
rect 1932 19742 1934 19794
rect 1934 19742 1986 19794
rect 1986 19742 1988 19794
rect 1932 19740 1988 19742
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 12460 19964 12516 20020
rect 12684 19964 12740 20020
rect 12348 19852 12404 19908
rect 4284 19234 4340 19236
rect 4284 19182 4286 19234
rect 4286 19182 4338 19234
rect 4338 19182 4340 19234
rect 4284 19180 4340 19182
rect 12348 19180 12404 19236
rect 1932 18844 1988 18900
rect 13132 19906 13188 19908
rect 13132 19854 13134 19906
rect 13134 19854 13186 19906
rect 13186 19854 13188 19906
rect 13132 19852 13188 19854
rect 13356 19516 13412 19572
rect 14252 21868 14308 21924
rect 14924 22092 14980 22148
rect 15372 21810 15428 21812
rect 15372 21758 15374 21810
rect 15374 21758 15426 21810
rect 15426 21758 15428 21810
rect 15372 21756 15428 21758
rect 14812 20914 14868 20916
rect 14812 20862 14814 20914
rect 14814 20862 14866 20914
rect 14866 20862 14868 20914
rect 14812 20860 14868 20862
rect 15148 21532 15204 21588
rect 13692 19964 13748 20020
rect 14252 20018 14308 20020
rect 14252 19966 14254 20018
rect 14254 19966 14306 20018
rect 14306 19966 14308 20018
rect 14252 19964 14308 19966
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 14364 19068 14420 19124
rect 15596 19964 15652 20020
rect 15148 19852 15204 19908
rect 15596 19516 15652 19572
rect 15372 19068 15428 19124
rect 14588 18956 14644 19012
rect 15708 19010 15764 19012
rect 15708 18958 15710 19010
rect 15710 18958 15762 19010
rect 15762 18958 15764 19010
rect 15708 18956 15764 18958
rect 14924 18508 14980 18564
rect 15820 18396 15876 18452
rect 13804 17500 13860 17556
rect 17388 27074 17444 27076
rect 17388 27022 17390 27074
rect 17390 27022 17442 27074
rect 17442 27022 17444 27074
rect 17388 27020 17444 27022
rect 17612 26962 17668 26964
rect 17612 26910 17614 26962
rect 17614 26910 17666 26962
rect 17666 26910 17668 26962
rect 17612 26908 17668 26910
rect 17948 27074 18004 27076
rect 17948 27022 17950 27074
rect 17950 27022 18002 27074
rect 18002 27022 18004 27074
rect 17948 27020 18004 27022
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 18508 27858 18564 27860
rect 18508 27806 18510 27858
rect 18510 27806 18562 27858
rect 18562 27806 18564 27858
rect 18508 27804 18564 27806
rect 18508 27580 18564 27636
rect 19068 27804 19124 27860
rect 18620 27244 18676 27300
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 26908 37436 26964 37492
rect 28140 37490 28196 37492
rect 28140 37438 28142 37490
rect 28142 37438 28194 37490
rect 28194 37438 28196 37490
rect 28140 37436 28196 37438
rect 19628 27074 19684 27076
rect 19628 27022 19630 27074
rect 19630 27022 19682 27074
rect 19682 27022 19684 27074
rect 19628 27020 19684 27022
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 40236 36370 40292 36372
rect 40236 36318 40238 36370
rect 40238 36318 40290 36370
rect 40290 36318 40292 36370
rect 40236 36316 40292 36318
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 21420 27074 21476 27076
rect 21420 27022 21422 27074
rect 21422 27022 21474 27074
rect 21474 27022 21476 27074
rect 21420 27020 21476 27022
rect 20860 26908 20916 26964
rect 18060 26348 18116 26404
rect 18508 26402 18564 26404
rect 18508 26350 18510 26402
rect 18510 26350 18562 26402
rect 18562 26350 18564 26402
rect 18508 26348 18564 26350
rect 16940 24668 16996 24724
rect 16940 24050 16996 24052
rect 16940 23998 16942 24050
rect 16942 23998 16994 24050
rect 16994 23998 16996 24050
rect 16940 23996 16996 23998
rect 16492 23772 16548 23828
rect 16716 23324 16772 23380
rect 17612 23938 17668 23940
rect 17612 23886 17614 23938
rect 17614 23886 17666 23938
rect 17666 23886 17668 23938
rect 17612 23884 17668 23886
rect 17948 23938 18004 23940
rect 17948 23886 17950 23938
rect 17950 23886 18002 23938
rect 18002 23886 18004 23938
rect 17948 23884 18004 23886
rect 17836 23772 17892 23828
rect 17500 23660 17556 23716
rect 17724 23714 17780 23716
rect 17724 23662 17726 23714
rect 17726 23662 17778 23714
rect 17778 23662 17780 23714
rect 17724 23660 17780 23662
rect 17388 23324 17444 23380
rect 16716 22316 16772 22372
rect 16604 22204 16660 22260
rect 16156 21756 16212 21812
rect 16380 21756 16436 21812
rect 16268 21420 16324 21476
rect 16044 18956 16100 19012
rect 16044 17052 16100 17108
rect 13132 16882 13188 16884
rect 13132 16830 13134 16882
rect 13134 16830 13186 16882
rect 13186 16830 13188 16882
rect 13132 16828 13188 16830
rect 15372 16828 15428 16884
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 14028 14476 14084 14532
rect 17836 22370 17892 22372
rect 17836 22318 17838 22370
rect 17838 22318 17890 22370
rect 17890 22318 17892 22370
rect 17836 22316 17892 22318
rect 16716 22146 16772 22148
rect 16716 22094 16718 22146
rect 16718 22094 16770 22146
rect 16770 22094 16772 22146
rect 16716 22092 16772 22094
rect 16940 21980 16996 22036
rect 16716 19906 16772 19908
rect 16716 19854 16718 19906
rect 16718 19854 16770 19906
rect 16770 19854 16772 19906
rect 16716 19852 16772 19854
rect 16604 19740 16660 19796
rect 16492 19180 16548 19236
rect 16268 19122 16324 19124
rect 16268 19070 16270 19122
rect 16270 19070 16322 19122
rect 16322 19070 16324 19122
rect 16268 19068 16324 19070
rect 16828 19068 16884 19124
rect 17276 22204 17332 22260
rect 17500 22146 17556 22148
rect 17500 22094 17502 22146
rect 17502 22094 17554 22146
rect 17554 22094 17556 22146
rect 17500 22092 17556 22094
rect 17388 21474 17444 21476
rect 17388 21422 17390 21474
rect 17390 21422 17442 21474
rect 17442 21422 17444 21474
rect 17388 21420 17444 21422
rect 17500 20130 17556 20132
rect 17500 20078 17502 20130
rect 17502 20078 17554 20130
rect 17554 20078 17556 20130
rect 17500 20076 17556 20078
rect 17836 19964 17892 20020
rect 17500 19234 17556 19236
rect 17500 19182 17502 19234
rect 17502 19182 17554 19234
rect 17554 19182 17556 19234
rect 17500 19180 17556 19182
rect 17836 19068 17892 19124
rect 16940 18508 16996 18564
rect 17612 19010 17668 19012
rect 17612 18958 17614 19010
rect 17614 18958 17666 19010
rect 17666 18958 17668 19010
rect 17612 18956 17668 18958
rect 18060 23154 18116 23156
rect 18060 23102 18062 23154
rect 18062 23102 18114 23154
rect 18114 23102 18116 23154
rect 18060 23100 18116 23102
rect 19628 25340 19684 25396
rect 18732 23884 18788 23940
rect 18172 22988 18228 23044
rect 18284 22204 18340 22260
rect 18620 23100 18676 23156
rect 18732 22316 18788 22372
rect 18508 22092 18564 22148
rect 18508 21532 18564 21588
rect 18396 21474 18452 21476
rect 18396 21422 18398 21474
rect 18398 21422 18450 21474
rect 18450 21422 18452 21474
rect 18396 21420 18452 21422
rect 18172 20636 18228 20692
rect 18508 19740 18564 19796
rect 17164 18284 17220 18340
rect 17388 18396 17444 18452
rect 17724 18396 17780 18452
rect 17724 17890 17780 17892
rect 17724 17838 17726 17890
rect 17726 17838 17778 17890
rect 17778 17838 17780 17890
rect 17724 17836 17780 17838
rect 17612 17778 17668 17780
rect 17612 17726 17614 17778
rect 17614 17726 17666 17778
rect 17666 17726 17668 17778
rect 17612 17724 17668 17726
rect 17276 17554 17332 17556
rect 17276 17502 17278 17554
rect 17278 17502 17330 17554
rect 17330 17502 17332 17554
rect 17276 17500 17332 17502
rect 18060 18338 18116 18340
rect 18060 18286 18062 18338
rect 18062 18286 18114 18338
rect 18114 18286 18116 18338
rect 18060 18284 18116 18286
rect 17836 17500 17892 17556
rect 16380 16882 16436 16884
rect 16380 16830 16382 16882
rect 16382 16830 16434 16882
rect 16434 16830 16436 16882
rect 16380 16828 16436 16830
rect 18172 17442 18228 17444
rect 18172 17390 18174 17442
rect 18174 17390 18226 17442
rect 18226 17390 18228 17442
rect 18172 17388 18228 17390
rect 16044 15484 16100 15540
rect 19292 23042 19348 23044
rect 19292 22990 19294 23042
rect 19294 22990 19346 23042
rect 19346 22990 19348 23042
rect 19292 22988 19348 22990
rect 19292 22092 19348 22148
rect 19180 21420 19236 21476
rect 19068 19180 19124 19236
rect 18844 19068 18900 19124
rect 18732 18620 18788 18676
rect 18956 18956 19012 19012
rect 18844 18562 18900 18564
rect 18844 18510 18846 18562
rect 18846 18510 18898 18562
rect 18898 18510 18900 18562
rect 18844 18508 18900 18510
rect 18620 18450 18676 18452
rect 18620 18398 18622 18450
rect 18622 18398 18674 18450
rect 18674 18398 18676 18450
rect 18620 18396 18676 18398
rect 18620 15484 18676 15540
rect 18956 17724 19012 17780
rect 15372 14530 15428 14532
rect 15372 14478 15374 14530
rect 15374 14478 15426 14530
rect 15426 14478 15428 14530
rect 15372 14476 15428 14478
rect 14700 14252 14756 14308
rect 18284 14364 18340 14420
rect 15372 13916 15428 13972
rect 17500 13970 17556 13972
rect 17500 13918 17502 13970
rect 17502 13918 17554 13970
rect 17554 13918 17556 13970
rect 17500 13916 17556 13918
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 18732 14418 18788 14420
rect 18732 14366 18734 14418
rect 18734 14366 18786 14418
rect 18786 14366 18788 14418
rect 18732 14364 18788 14366
rect 18620 14306 18676 14308
rect 18620 14254 18622 14306
rect 18622 14254 18674 14306
rect 18674 14254 18676 14306
rect 18620 14252 18676 14254
rect 18396 13916 18452 13972
rect 19068 17442 19124 17444
rect 19068 17390 19070 17442
rect 19070 17390 19122 17442
rect 19122 17390 19124 17442
rect 19068 17388 19124 17390
rect 20188 25340 20244 25396
rect 19628 25116 19684 25172
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 20300 25228 20356 25284
rect 20188 24556 20244 24612
rect 19852 24498 19908 24500
rect 19852 24446 19854 24498
rect 19854 24446 19906 24498
rect 19906 24446 19908 24498
rect 19852 24444 19908 24446
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 19740 23100 19796 23156
rect 19628 22652 19684 22708
rect 20748 24722 20804 24724
rect 20748 24670 20750 24722
rect 20750 24670 20802 24722
rect 20802 24670 20804 24722
rect 20748 24668 20804 24670
rect 21084 26348 21140 26404
rect 22652 26402 22708 26404
rect 22652 26350 22654 26402
rect 22654 26350 22706 26402
rect 22706 26350 22708 26402
rect 22652 26348 22708 26350
rect 23212 26348 23268 26404
rect 22652 26066 22708 26068
rect 22652 26014 22654 26066
rect 22654 26014 22706 26066
rect 22706 26014 22708 26066
rect 22652 26012 22708 26014
rect 21308 25394 21364 25396
rect 21308 25342 21310 25394
rect 21310 25342 21362 25394
rect 21362 25342 21364 25394
rect 21308 25340 21364 25342
rect 21644 24780 21700 24836
rect 20748 24444 20804 24500
rect 20300 23826 20356 23828
rect 20300 23774 20302 23826
rect 20302 23774 20354 23826
rect 20354 23774 20356 23826
rect 20300 23772 20356 23774
rect 21308 24610 21364 24612
rect 21308 24558 21310 24610
rect 21310 24558 21362 24610
rect 21362 24558 21364 24610
rect 21308 24556 21364 24558
rect 22316 24780 22372 24836
rect 21756 24668 21812 24724
rect 23548 26290 23604 26292
rect 23548 26238 23550 26290
rect 23550 26238 23602 26290
rect 23602 26238 23604 26290
rect 23548 26236 23604 26238
rect 22428 24556 22484 24612
rect 22316 24444 22372 24500
rect 21980 24108 22036 24164
rect 21756 23884 21812 23940
rect 21868 23772 21924 23828
rect 20188 22540 20244 22596
rect 19740 22370 19796 22372
rect 19740 22318 19742 22370
rect 19742 22318 19794 22370
rect 19794 22318 19796 22370
rect 19740 22316 19796 22318
rect 19628 22092 19684 22148
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 20412 22316 20468 22372
rect 21644 23266 21700 23268
rect 21644 23214 21646 23266
rect 21646 23214 21698 23266
rect 21698 23214 21700 23266
rect 21644 23212 21700 23214
rect 20524 22428 20580 22484
rect 20188 21756 20244 21812
rect 20300 22092 20356 22148
rect 20076 20802 20132 20804
rect 20076 20750 20078 20802
rect 20078 20750 20130 20802
rect 20130 20750 20132 20802
rect 20076 20748 20132 20750
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 20412 21586 20468 21588
rect 20412 21534 20414 21586
rect 20414 21534 20466 21586
rect 20466 21534 20468 21586
rect 20412 21532 20468 21534
rect 20748 22764 20804 22820
rect 20636 22204 20692 22260
rect 21420 22258 21476 22260
rect 21420 22206 21422 22258
rect 21422 22206 21474 22258
rect 21474 22206 21476 22258
rect 21420 22204 21476 22206
rect 20524 20636 20580 20692
rect 20412 20300 20468 20356
rect 22316 23548 22372 23604
rect 24444 27020 24500 27076
rect 24780 27074 24836 27076
rect 24780 27022 24782 27074
rect 24782 27022 24834 27074
rect 24834 27022 24836 27074
rect 24780 27020 24836 27022
rect 25228 27020 25284 27076
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 25452 26402 25508 26404
rect 25452 26350 25454 26402
rect 25454 26350 25506 26402
rect 25506 26350 25508 26402
rect 25452 26348 25508 26350
rect 24892 26236 24948 26292
rect 25676 26290 25732 26292
rect 25676 26238 25678 26290
rect 25678 26238 25730 26290
rect 25730 26238 25732 26290
rect 25676 26236 25732 26238
rect 25900 26178 25956 26180
rect 25900 26126 25902 26178
rect 25902 26126 25954 26178
rect 25954 26126 25956 26178
rect 25900 26124 25956 26126
rect 25340 26012 25396 26068
rect 27132 27132 27188 27188
rect 26572 26514 26628 26516
rect 26572 26462 26574 26514
rect 26574 26462 26626 26514
rect 26626 26462 26628 26514
rect 26572 26460 26628 26462
rect 27692 27186 27748 27188
rect 27692 27134 27694 27186
rect 27694 27134 27746 27186
rect 27746 27134 27748 27186
rect 27692 27132 27748 27134
rect 27356 27020 27412 27076
rect 26124 26290 26180 26292
rect 26124 26238 26126 26290
rect 26126 26238 26178 26290
rect 26178 26238 26180 26290
rect 26124 26236 26180 26238
rect 27020 26290 27076 26292
rect 27020 26238 27022 26290
rect 27022 26238 27074 26290
rect 27074 26238 27076 26290
rect 27020 26236 27076 26238
rect 26684 26124 26740 26180
rect 22652 24108 22708 24164
rect 22540 23660 22596 23716
rect 21756 22764 21812 22820
rect 21868 23212 21924 23268
rect 21644 22146 21700 22148
rect 21644 22094 21646 22146
rect 21646 22094 21698 22146
rect 21698 22094 21700 22146
rect 21644 22092 21700 22094
rect 19404 20076 19460 20132
rect 19516 19234 19572 19236
rect 19516 19182 19518 19234
rect 19518 19182 19570 19234
rect 19570 19182 19572 19234
rect 19516 19180 19572 19182
rect 19964 19964 20020 20020
rect 19964 19740 20020 19796
rect 19292 19122 19348 19124
rect 19292 19070 19294 19122
rect 19294 19070 19346 19122
rect 19346 19070 19348 19122
rect 19292 19068 19348 19070
rect 19292 18226 19348 18228
rect 19292 18174 19294 18226
rect 19294 18174 19346 18226
rect 19346 18174 19348 18226
rect 19292 18172 19348 18174
rect 19292 17836 19348 17892
rect 19852 19122 19908 19124
rect 19852 19070 19854 19122
rect 19854 19070 19906 19122
rect 19906 19070 19908 19122
rect 19852 19068 19908 19070
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 19628 18674 19684 18676
rect 19628 18622 19630 18674
rect 19630 18622 19682 18674
rect 19682 18622 19684 18674
rect 19628 18620 19684 18622
rect 20188 18060 20244 18116
rect 20524 20076 20580 20132
rect 20636 19964 20692 20020
rect 20748 20300 20804 20356
rect 20524 19292 20580 19348
rect 21868 20748 21924 20804
rect 21420 20690 21476 20692
rect 21420 20638 21422 20690
rect 21422 20638 21474 20690
rect 21474 20638 21476 20690
rect 21420 20636 21476 20638
rect 21532 20412 21588 20468
rect 21308 19292 21364 19348
rect 21420 19180 21476 19236
rect 21084 18396 21140 18452
rect 21196 18732 21252 18788
rect 20748 18226 20804 18228
rect 20748 18174 20750 18226
rect 20750 18174 20802 18226
rect 20802 18174 20804 18226
rect 20748 18172 20804 18174
rect 22540 22652 22596 22708
rect 22204 21644 22260 21700
rect 22204 20412 22260 20468
rect 21980 20132 22036 20188
rect 21868 19964 21924 20020
rect 21756 19740 21812 19796
rect 22540 22204 22596 22260
rect 22876 23938 22932 23940
rect 22876 23886 22878 23938
rect 22878 23886 22930 23938
rect 22930 23886 22932 23938
rect 22876 23884 22932 23886
rect 23212 23826 23268 23828
rect 23212 23774 23214 23826
rect 23214 23774 23266 23826
rect 23266 23774 23268 23826
rect 23212 23772 23268 23774
rect 23212 23548 23268 23604
rect 23100 23266 23156 23268
rect 23100 23214 23102 23266
rect 23102 23214 23154 23266
rect 23154 23214 23156 23266
rect 23100 23212 23156 23214
rect 23996 23324 24052 23380
rect 22988 23154 23044 23156
rect 22988 23102 22990 23154
rect 22990 23102 23042 23154
rect 23042 23102 23044 23154
rect 22988 23100 23044 23102
rect 22876 22764 22932 22820
rect 22988 22652 23044 22708
rect 22652 21586 22708 21588
rect 22652 21534 22654 21586
rect 22654 21534 22706 21586
rect 22706 21534 22708 21586
rect 22652 21532 22708 21534
rect 22540 21420 22596 21476
rect 24220 23378 24276 23380
rect 24220 23326 24222 23378
rect 24222 23326 24274 23378
rect 24274 23326 24276 23378
rect 24220 23324 24276 23326
rect 23548 22428 23604 22484
rect 23772 21698 23828 21700
rect 23772 21646 23774 21698
rect 23774 21646 23826 21698
rect 23826 21646 23828 21698
rect 23772 21644 23828 21646
rect 23212 21420 23268 21476
rect 22764 20132 22820 20188
rect 23100 19740 23156 19796
rect 22988 19180 23044 19236
rect 22764 18562 22820 18564
rect 22764 18510 22766 18562
rect 22766 18510 22818 18562
rect 22818 18510 22820 18562
rect 22764 18508 22820 18510
rect 21980 18450 22036 18452
rect 21980 18398 21982 18450
rect 21982 18398 22034 18450
rect 22034 18398 22036 18450
rect 21980 18396 22036 18398
rect 22652 18338 22708 18340
rect 22652 18286 22654 18338
rect 22654 18286 22706 18338
rect 22706 18286 22708 18338
rect 22652 18284 22708 18286
rect 21644 18060 21700 18116
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 19740 17106 19796 17108
rect 19740 17054 19742 17106
rect 19742 17054 19794 17106
rect 19794 17054 19796 17106
rect 19740 17052 19796 17054
rect 20748 17554 20804 17556
rect 20748 17502 20750 17554
rect 20750 17502 20802 17554
rect 20802 17502 20804 17554
rect 20748 17500 20804 17502
rect 21196 17052 21252 17108
rect 22652 17778 22708 17780
rect 22652 17726 22654 17778
rect 22654 17726 22706 17778
rect 22706 17726 22708 17778
rect 22652 17724 22708 17726
rect 21644 17666 21700 17668
rect 21644 17614 21646 17666
rect 21646 17614 21698 17666
rect 21698 17614 21700 17666
rect 21644 17612 21700 17614
rect 22540 17666 22596 17668
rect 22540 17614 22542 17666
rect 22542 17614 22594 17666
rect 22594 17614 22596 17666
rect 22540 17612 22596 17614
rect 21868 17554 21924 17556
rect 21868 17502 21870 17554
rect 21870 17502 21922 17554
rect 21922 17502 21924 17554
rect 21868 17500 21924 17502
rect 22988 18060 23044 18116
rect 23100 18732 23156 18788
rect 22876 17554 22932 17556
rect 22876 17502 22878 17554
rect 22878 17502 22930 17554
rect 22930 17502 22932 17554
rect 22876 17500 22932 17502
rect 21756 17442 21812 17444
rect 21756 17390 21758 17442
rect 21758 17390 21810 17442
rect 21810 17390 21812 17442
rect 21756 17388 21812 17390
rect 20524 16940 20580 16996
rect 19180 16716 19236 16772
rect 19964 16716 20020 16772
rect 21308 16716 21364 16772
rect 22540 17106 22596 17108
rect 22540 17054 22542 17106
rect 22542 17054 22594 17106
rect 22594 17054 22596 17106
rect 22540 17052 22596 17054
rect 22204 16994 22260 16996
rect 22204 16942 22206 16994
rect 22206 16942 22258 16994
rect 22258 16942 22260 16994
rect 22204 16940 22260 16942
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 21308 15538 21364 15540
rect 21308 15486 21310 15538
rect 21310 15486 21362 15538
rect 21362 15486 21364 15538
rect 21308 15484 21364 15486
rect 22540 15538 22596 15540
rect 22540 15486 22542 15538
rect 22542 15486 22594 15538
rect 22594 15486 22596 15538
rect 22540 15484 22596 15486
rect 21756 15148 21812 15204
rect 22652 15260 22708 15316
rect 19292 14364 19348 14420
rect 20636 14418 20692 14420
rect 20636 14366 20638 14418
rect 20638 14366 20690 14418
rect 20690 14366 20692 14418
rect 20636 14364 20692 14366
rect 23436 21474 23492 21476
rect 23436 21422 23438 21474
rect 23438 21422 23490 21474
rect 23490 21422 23492 21474
rect 23436 21420 23492 21422
rect 26684 25340 26740 25396
rect 28140 27074 28196 27076
rect 28140 27022 28142 27074
rect 28142 27022 28194 27074
rect 28194 27022 28196 27074
rect 28140 27020 28196 27022
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 28700 27020 28756 27076
rect 37660 27074 37716 27076
rect 37660 27022 37662 27074
rect 37662 27022 37714 27074
rect 37714 27022 37716 27074
rect 37660 27020 37716 27022
rect 40012 26908 40068 26964
rect 28028 26460 28084 26516
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 29260 25452 29316 25508
rect 30604 25452 30660 25508
rect 29372 25394 29428 25396
rect 29372 25342 29374 25394
rect 29374 25342 29426 25394
rect 29426 25342 29428 25394
rect 29372 25340 29428 25342
rect 25340 23660 25396 23716
rect 26236 23324 26292 23380
rect 24332 23042 24388 23044
rect 24332 22990 24334 23042
rect 24334 22990 24386 23042
rect 24386 22990 24388 23042
rect 24332 22988 24388 22990
rect 25452 22988 25508 23044
rect 24220 22540 24276 22596
rect 25340 22428 25396 22484
rect 24444 21532 24500 21588
rect 23436 19964 23492 20020
rect 23660 18844 23716 18900
rect 23548 18396 23604 18452
rect 23436 18284 23492 18340
rect 23212 15484 23268 15540
rect 21980 14364 22036 14420
rect 22316 14418 22372 14420
rect 22316 14366 22318 14418
rect 22318 14366 22370 14418
rect 22370 14366 22372 14418
rect 22316 14364 22372 14366
rect 24556 19964 24612 20020
rect 24556 19292 24612 19348
rect 25676 21810 25732 21812
rect 25676 21758 25678 21810
rect 25678 21758 25730 21810
rect 25730 21758 25732 21810
rect 25676 21756 25732 21758
rect 26908 23266 26964 23268
rect 26908 23214 26910 23266
rect 26910 23214 26962 23266
rect 26962 23214 26964 23266
rect 26908 23212 26964 23214
rect 26572 22988 26628 23044
rect 28476 24610 28532 24612
rect 28476 24558 28478 24610
rect 28478 24558 28530 24610
rect 28530 24558 28532 24610
rect 28476 24556 28532 24558
rect 28140 23154 28196 23156
rect 28140 23102 28142 23154
rect 28142 23102 28194 23154
rect 28194 23102 28196 23154
rect 28140 23100 28196 23102
rect 27692 22428 27748 22484
rect 28140 22540 28196 22596
rect 26572 21698 26628 21700
rect 26572 21646 26574 21698
rect 26574 21646 26626 21698
rect 26626 21646 26628 21698
rect 26572 21644 26628 21646
rect 25228 21586 25284 21588
rect 25228 21534 25230 21586
rect 25230 21534 25282 21586
rect 25282 21534 25284 21586
rect 25228 21532 25284 21534
rect 25788 21420 25844 21476
rect 28140 21756 28196 21812
rect 24668 19852 24724 19908
rect 25228 20018 25284 20020
rect 25228 19966 25230 20018
rect 25230 19966 25282 20018
rect 25282 19966 25284 20018
rect 25228 19964 25284 19966
rect 25116 19740 25172 19796
rect 24332 18844 24388 18900
rect 24444 18732 24500 18788
rect 24108 18620 24164 18676
rect 23996 18562 24052 18564
rect 23996 18510 23998 18562
rect 23998 18510 24050 18562
rect 24050 18510 24052 18562
rect 23996 18508 24052 18510
rect 26684 20130 26740 20132
rect 26684 20078 26686 20130
rect 26686 20078 26738 20130
rect 26738 20078 26740 20130
rect 26684 20076 26740 20078
rect 26908 20018 26964 20020
rect 26908 19966 26910 20018
rect 26910 19966 26962 20018
rect 26962 19966 26964 20018
rect 26908 19964 26964 19966
rect 25676 19292 25732 19348
rect 25004 19010 25060 19012
rect 25004 18958 25006 19010
rect 25006 18958 25058 19010
rect 25058 18958 25060 19010
rect 25004 18956 25060 18958
rect 25788 19234 25844 19236
rect 25788 19182 25790 19234
rect 25790 19182 25842 19234
rect 25842 19182 25844 19234
rect 25788 19180 25844 19182
rect 25676 18396 25732 18452
rect 23884 18284 23940 18340
rect 23548 14364 23604 14420
rect 23660 17724 23716 17780
rect 20076 14252 20132 14308
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 20076 13970 20132 13972
rect 20076 13918 20078 13970
rect 20078 13918 20130 13970
rect 20130 13918 20132 13970
rect 20076 13916 20132 13918
rect 19852 13858 19908 13860
rect 19852 13806 19854 13858
rect 19854 13806 19906 13858
rect 19906 13806 19908 13858
rect 19852 13804 19908 13806
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 18620 13468 18676 13524
rect 21084 14252 21140 14308
rect 20748 13804 20804 13860
rect 20412 13746 20468 13748
rect 20412 13694 20414 13746
rect 20414 13694 20466 13746
rect 20466 13694 20468 13746
rect 20412 13692 20468 13694
rect 20188 13468 20244 13524
rect 21868 14306 21924 14308
rect 21868 14254 21870 14306
rect 21870 14254 21922 14306
rect 21922 14254 21924 14306
rect 21868 14252 21924 14254
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 22652 13692 22708 13748
rect 23436 14306 23492 14308
rect 23436 14254 23438 14306
rect 23438 14254 23490 14306
rect 23490 14254 23492 14306
rect 23436 14252 23492 14254
rect 23436 13692 23492 13748
rect 24444 17554 24500 17556
rect 24444 17502 24446 17554
rect 24446 17502 24498 17554
rect 24498 17502 24500 17554
rect 24444 17500 24500 17502
rect 23884 17052 23940 17108
rect 24220 17388 24276 17444
rect 24556 17442 24612 17444
rect 24556 17390 24558 17442
rect 24558 17390 24610 17442
rect 24610 17390 24612 17442
rect 24556 17388 24612 17390
rect 25452 17388 25508 17444
rect 24332 17106 24388 17108
rect 24332 17054 24334 17106
rect 24334 17054 24386 17106
rect 24386 17054 24388 17106
rect 24332 17052 24388 17054
rect 25452 16940 25508 16996
rect 23884 14364 23940 14420
rect 28700 23212 28756 23268
rect 28588 23154 28644 23156
rect 28588 23102 28590 23154
rect 28590 23102 28642 23154
rect 28642 23102 28644 23154
rect 28588 23100 28644 23102
rect 28588 22482 28644 22484
rect 28588 22430 28590 22482
rect 28590 22430 28642 22482
rect 28642 22430 28644 22482
rect 28588 22428 28644 22430
rect 29260 24556 29316 24612
rect 37660 25506 37716 25508
rect 37660 25454 37662 25506
rect 37662 25454 37714 25506
rect 37714 25454 37716 25506
rect 37660 25452 37716 25454
rect 40012 24892 40068 24948
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 29484 23938 29540 23940
rect 29484 23886 29486 23938
rect 29486 23886 29538 23938
rect 29538 23886 29540 23938
rect 29484 23884 29540 23886
rect 29596 23212 29652 23268
rect 29932 23100 29988 23156
rect 30828 23100 30884 23156
rect 29932 22258 29988 22260
rect 29932 22206 29934 22258
rect 29934 22206 29986 22258
rect 29986 22206 29988 22258
rect 29932 22204 29988 22206
rect 37660 23154 37716 23156
rect 37660 23102 37662 23154
rect 37662 23102 37714 23154
rect 37714 23102 37716 23154
rect 37660 23100 37716 23102
rect 40012 22930 40068 22932
rect 40012 22878 40014 22930
rect 40014 22878 40066 22930
rect 40066 22878 40068 22930
rect 40012 22876 40068 22878
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 37660 22370 37716 22372
rect 37660 22318 37662 22370
rect 37662 22318 37714 22370
rect 37714 22318 37716 22370
rect 37660 22316 37716 22318
rect 30828 22204 30884 22260
rect 29372 21420 29428 21476
rect 40012 22204 40068 22260
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 37660 20802 37716 20804
rect 37660 20750 37662 20802
rect 37662 20750 37714 20802
rect 37714 20750 37716 20802
rect 37660 20748 37716 20750
rect 28364 19964 28420 20020
rect 27580 19180 27636 19236
rect 28588 19346 28644 19348
rect 28588 19294 28590 19346
rect 28590 19294 28642 19346
rect 28642 19294 28644 19346
rect 28588 19292 28644 19294
rect 28364 19180 28420 19236
rect 29260 20578 29316 20580
rect 29260 20526 29262 20578
rect 29262 20526 29314 20578
rect 29314 20526 29316 20578
rect 29260 20524 29316 20526
rect 30828 20524 30884 20580
rect 40012 20188 40068 20244
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 40012 19516 40068 19572
rect 37660 19292 37716 19348
rect 26012 18844 26068 18900
rect 29596 19234 29652 19236
rect 29596 19182 29598 19234
rect 29598 19182 29650 19234
rect 29650 19182 29652 19234
rect 29596 19180 29652 19182
rect 29372 18620 29428 18676
rect 27020 17612 27076 17668
rect 27020 17052 27076 17108
rect 26684 16994 26740 16996
rect 26684 16942 26686 16994
rect 26686 16942 26738 16994
rect 26738 16942 26740 16994
rect 26684 16940 26740 16942
rect 26012 16716 26068 16772
rect 26124 15820 26180 15876
rect 25228 15314 25284 15316
rect 25228 15262 25230 15314
rect 25230 15262 25282 15314
rect 25282 15262 25284 15314
rect 25228 15260 25284 15262
rect 25452 15260 25508 15316
rect 24220 14252 24276 14308
rect 25788 15314 25844 15316
rect 25788 15262 25790 15314
rect 25790 15262 25842 15314
rect 25842 15262 25844 15314
rect 25788 15260 25844 15262
rect 26460 16268 26516 16324
rect 27356 16716 27412 16772
rect 27468 16322 27524 16324
rect 27468 16270 27470 16322
rect 27470 16270 27522 16322
rect 27522 16270 27524 16322
rect 27468 16268 27524 16270
rect 26236 15260 26292 15316
rect 25564 14476 25620 14532
rect 26908 14588 26964 14644
rect 25340 14252 25396 14308
rect 26684 14476 26740 14532
rect 24108 13746 24164 13748
rect 24108 13694 24110 13746
rect 24110 13694 24162 13746
rect 24162 13694 24164 13746
rect 24108 13692 24164 13694
rect 25340 13746 25396 13748
rect 25340 13694 25342 13746
rect 25342 13694 25394 13746
rect 25394 13694 25396 13746
rect 25340 13692 25396 13694
rect 22876 3612 22932 3668
rect 20188 3388 20244 3444
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 21756 3388 21812 3444
rect 28028 15874 28084 15876
rect 28028 15822 28030 15874
rect 28030 15822 28082 15874
rect 28082 15822 28084 15874
rect 28028 15820 28084 15822
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 37660 17666 37716 17668
rect 37660 17614 37662 17666
rect 37662 17614 37714 17666
rect 37714 17614 37716 17666
rect 37660 17612 37716 17614
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 28812 15820 28868 15876
rect 29260 15820 29316 15876
rect 27468 15148 27524 15204
rect 29036 15202 29092 15204
rect 29036 15150 29038 15202
rect 29038 15150 29090 15202
rect 29090 15150 29092 15202
rect 29036 15148 29092 15150
rect 28252 14642 28308 14644
rect 28252 14590 28254 14642
rect 28254 14590 28306 14642
rect 28306 14590 28308 14642
rect 28252 14588 28308 14590
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 40012 16828 40068 16884
rect 40012 16156 40068 16212
rect 37884 15148 37940 15204
rect 40012 14812 40068 14868
rect 37660 14588 37716 14644
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 40236 8764 40292 8820
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 24892 4060 24948 4116
rect 23212 3500 23268 3556
rect 24556 3554 24612 3556
rect 24556 3502 24558 3554
rect 24558 3502 24610 3554
rect 24610 3502 24612 3554
rect 24556 3500 24612 3502
rect 26236 4114 26292 4116
rect 26236 4062 26238 4114
rect 26238 4062 26290 4114
rect 26290 4062 26292 4114
rect 26236 4060 26292 4062
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 25564 3666 25620 3668
rect 25564 3614 25566 3666
rect 25566 3614 25618 3666
rect 25618 3614 25620 3666
rect 25564 3612 25620 3614
<< metal3 >>
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 17490 38220 17500 38276
rect 17556 38220 18620 38276
rect 18676 38220 18686 38276
rect 20850 38220 20860 38276
rect 20916 38220 22092 38276
rect 22148 38220 22158 38276
rect 23538 38220 23548 38276
rect 23604 38220 25564 38276
rect 25620 38220 25630 38276
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 16818 37436 16828 37492
rect 16884 37436 18396 37492
rect 18452 37436 18462 37492
rect 26898 37436 26908 37492
rect 26964 37436 28140 37492
rect 28196 37436 28206 37492
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 16146 36652 16156 36708
rect 16212 36652 17388 36708
rect 17444 36652 17454 36708
rect 41200 36372 42000 36400
rect 40226 36316 40236 36372
rect 40292 36316 42000 36372
rect 41200 36288 42000 36316
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 16258 28476 16268 28532
rect 16324 28476 16940 28532
rect 16996 28476 17006 28532
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 13906 27804 13916 27860
rect 13972 27804 14364 27860
rect 14420 27804 16380 27860
rect 16436 27804 18508 27860
rect 18564 27804 19068 27860
rect 19124 27804 19134 27860
rect 14690 27692 14700 27748
rect 14756 27692 17500 27748
rect 17556 27692 17566 27748
rect 0 27636 800 27664
rect 0 27580 10892 27636
rect 10948 27580 10958 27636
rect 16818 27580 16828 27636
rect 16884 27580 18508 27636
rect 18564 27580 18574 27636
rect 0 27552 800 27580
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 16146 27244 16156 27300
rect 16212 27244 17388 27300
rect 17444 27244 18620 27300
rect 18676 27244 18686 27300
rect 27122 27132 27132 27188
rect 27188 27132 27692 27188
rect 27748 27132 31948 27188
rect 31892 27076 31948 27132
rect 12898 27020 12908 27076
rect 12964 27020 14364 27076
rect 14420 27020 14430 27076
rect 16482 27020 16492 27076
rect 16548 27020 17388 27076
rect 17444 27020 17454 27076
rect 17938 27020 17948 27076
rect 18004 27020 19628 27076
rect 19684 27020 20188 27076
rect 21410 27020 21420 27076
rect 21476 27020 24444 27076
rect 24500 27020 24780 27076
rect 24836 27020 25228 27076
rect 25284 27020 27356 27076
rect 27412 27020 28140 27076
rect 28196 27020 28700 27076
rect 28756 27020 28766 27076
rect 31892 27020 37660 27076
rect 37716 27020 37726 27076
rect 20132 26964 20188 27020
rect 41200 26964 42000 26992
rect 15026 26908 15036 26964
rect 15092 26908 17612 26964
rect 17668 26908 17678 26964
rect 20132 26908 20860 26964
rect 20916 26908 20926 26964
rect 40002 26908 40012 26964
rect 40068 26908 42000 26964
rect 41200 26880 42000 26908
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 26562 26460 26572 26516
rect 26628 26460 28028 26516
rect 28084 26460 28094 26516
rect 18050 26348 18060 26404
rect 18116 26348 18508 26404
rect 18564 26348 21084 26404
rect 21140 26348 22652 26404
rect 22708 26348 22718 26404
rect 23202 26348 23212 26404
rect 23268 26348 25452 26404
rect 25508 26348 25518 26404
rect 23538 26236 23548 26292
rect 23604 26236 24892 26292
rect 24948 26236 25676 26292
rect 25732 26236 25742 26292
rect 26114 26236 26124 26292
rect 26180 26236 27020 26292
rect 27076 26236 27086 26292
rect 25890 26124 25900 26180
rect 25956 26124 26684 26180
rect 26740 26124 26750 26180
rect 22642 26012 22652 26068
rect 22708 26012 25340 26068
rect 25396 26012 25406 26068
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 29250 25452 29260 25508
rect 29316 25452 30604 25508
rect 30660 25452 37660 25508
rect 37716 25452 37726 25508
rect 19618 25340 19628 25396
rect 19684 25340 20188 25396
rect 20244 25340 21308 25396
rect 21364 25340 21374 25396
rect 26674 25340 26684 25396
rect 26740 25340 29372 25396
rect 29428 25340 29438 25396
rect 19628 25228 20300 25284
rect 20356 25228 20366 25284
rect 19628 25172 19684 25228
rect 19618 25116 19628 25172
rect 19684 25116 19694 25172
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 41200 24948 42000 24976
rect 40002 24892 40012 24948
rect 40068 24892 42000 24948
rect 41200 24864 42000 24892
rect 21634 24780 21644 24836
rect 21700 24780 22316 24836
rect 22372 24780 22382 24836
rect 4274 24668 4284 24724
rect 4340 24668 13076 24724
rect 16930 24668 16940 24724
rect 16996 24668 20748 24724
rect 20804 24668 21756 24724
rect 21812 24668 21822 24724
rect 13020 24612 13076 24668
rect 13010 24556 13020 24612
rect 13076 24556 16156 24612
rect 16212 24556 16222 24612
rect 20178 24556 20188 24612
rect 20244 24556 21308 24612
rect 21364 24556 22428 24612
rect 22484 24556 22494 24612
rect 28466 24556 28476 24612
rect 28532 24556 29260 24612
rect 29316 24556 29326 24612
rect 1922 24444 1932 24500
rect 1988 24444 1998 24500
rect 19842 24444 19852 24500
rect 19908 24444 20748 24500
rect 20804 24444 22316 24500
rect 22372 24444 22382 24500
rect 0 24276 800 24304
rect 1932 24276 1988 24444
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 0 24220 1988 24276
rect 0 24192 800 24220
rect 20132 24108 21980 24164
rect 22036 24108 22652 24164
rect 22708 24108 22718 24164
rect 8372 23996 9996 24052
rect 10052 23996 12796 24052
rect 12852 23996 12862 24052
rect 13794 23996 13804 24052
rect 13860 23996 16940 24052
rect 16996 23996 17006 24052
rect 8372 23940 8428 23996
rect 20132 23940 20188 24108
rect 4274 23884 4284 23940
rect 4340 23884 8428 23940
rect 15138 23884 15148 23940
rect 15204 23884 17612 23940
rect 17668 23884 17678 23940
rect 17938 23884 17948 23940
rect 18004 23884 18732 23940
rect 18788 23884 20188 23940
rect 21746 23884 21756 23940
rect 21812 23884 22148 23940
rect 22866 23884 22876 23940
rect 22932 23884 29484 23940
rect 29540 23884 29550 23940
rect 22092 23828 22148 23884
rect 12114 23772 12124 23828
rect 12180 23772 13580 23828
rect 13636 23772 13646 23828
rect 15586 23772 15596 23828
rect 15652 23772 15932 23828
rect 15988 23772 15998 23828
rect 16482 23772 16492 23828
rect 16548 23772 17836 23828
rect 17892 23772 17902 23828
rect 20132 23772 20300 23828
rect 20356 23772 21868 23828
rect 21924 23772 21934 23828
rect 22092 23772 23212 23828
rect 23268 23772 23278 23828
rect 15932 23716 15988 23772
rect 20132 23716 20188 23772
rect 15932 23660 17500 23716
rect 17556 23660 17566 23716
rect 17714 23660 17724 23716
rect 17780 23660 20188 23716
rect 22530 23660 22540 23716
rect 22596 23660 25340 23716
rect 25396 23660 25406 23716
rect 0 23604 800 23632
rect 17724 23604 17780 23660
rect 0 23548 1932 23604
rect 1988 23548 1998 23604
rect 13010 23548 13020 23604
rect 13076 23548 13468 23604
rect 13524 23548 13534 23604
rect 14130 23548 14140 23604
rect 14196 23548 17780 23604
rect 22306 23548 22316 23604
rect 22372 23548 23212 23604
rect 23268 23548 23278 23604
rect 0 23520 800 23548
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 13906 23436 13916 23492
rect 13972 23436 14924 23492
rect 14980 23436 15932 23492
rect 15988 23436 15998 23492
rect 16034 23324 16044 23380
rect 16100 23324 16716 23380
rect 16772 23324 17388 23380
rect 17444 23324 23996 23380
rect 24052 23324 24062 23380
rect 24210 23324 24220 23380
rect 24276 23324 26236 23380
rect 26292 23324 26302 23380
rect 24220 23268 24276 23324
rect 20132 23212 21644 23268
rect 21700 23212 21710 23268
rect 21858 23212 21868 23268
rect 21924 23212 23100 23268
rect 23156 23212 24276 23268
rect 26898 23212 26908 23268
rect 26964 23212 28700 23268
rect 28756 23212 29596 23268
rect 29652 23212 29662 23268
rect 12674 23100 12684 23156
rect 12740 23100 14140 23156
rect 14196 23100 14206 23156
rect 15810 23100 15820 23156
rect 15876 23100 18060 23156
rect 18116 23100 18126 23156
rect 18610 23100 18620 23156
rect 18676 23100 19740 23156
rect 19796 23100 19806 23156
rect 20132 23044 20188 23212
rect 22978 23100 22988 23156
rect 23044 23100 28140 23156
rect 28196 23100 28206 23156
rect 28578 23100 28588 23156
rect 28644 23100 29932 23156
rect 29988 23100 29998 23156
rect 30818 23100 30828 23156
rect 30884 23100 37660 23156
rect 37716 23100 37726 23156
rect 18162 22988 18172 23044
rect 18228 22988 19292 23044
rect 19348 22988 20188 23044
rect 24322 22988 24332 23044
rect 24388 22988 25452 23044
rect 25508 22988 26572 23044
rect 26628 22988 26638 23044
rect 41200 22932 42000 22960
rect 40002 22876 40012 22932
rect 40068 22876 42000 22932
rect 41200 22848 42000 22876
rect 20738 22764 20748 22820
rect 20804 22764 21756 22820
rect 21812 22764 22876 22820
rect 22932 22764 22942 22820
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 19618 22652 19628 22708
rect 19684 22652 22540 22708
rect 22596 22652 22988 22708
rect 23044 22652 23054 22708
rect 20178 22540 20188 22596
rect 20244 22540 24220 22596
rect 24276 22540 24286 22596
rect 28130 22540 28140 22596
rect 28196 22540 31948 22596
rect 18732 22428 20188 22484
rect 20514 22428 20524 22484
rect 20580 22428 23548 22484
rect 23604 22428 23614 22484
rect 25330 22428 25340 22484
rect 25396 22428 27692 22484
rect 27748 22428 28588 22484
rect 28644 22428 28654 22484
rect 18732 22372 18788 22428
rect 20132 22372 20188 22428
rect 31892 22372 31948 22540
rect 16706 22316 16716 22372
rect 16772 22316 17836 22372
rect 17892 22316 18732 22372
rect 18788 22316 18798 22372
rect 19730 22316 19740 22372
rect 19796 22316 19806 22372
rect 20132 22316 20412 22372
rect 20468 22316 20478 22372
rect 31892 22316 37660 22372
rect 37716 22316 37726 22372
rect 19740 22260 19796 22316
rect 41200 22260 42000 22288
rect 11554 22204 11564 22260
rect 11620 22204 13580 22260
rect 13636 22204 13646 22260
rect 16594 22204 16604 22260
rect 16660 22204 17276 22260
rect 17332 22204 18284 22260
rect 18340 22204 19348 22260
rect 19740 22204 20636 22260
rect 20692 22204 21420 22260
rect 21476 22204 22540 22260
rect 22596 22204 22606 22260
rect 29922 22204 29932 22260
rect 29988 22204 30828 22260
rect 30884 22204 30894 22260
rect 40002 22204 40012 22260
rect 40068 22204 42000 22260
rect 19292 22148 19348 22204
rect 41200 22176 42000 22204
rect 14914 22092 14924 22148
rect 14980 22092 16716 22148
rect 16772 22092 16782 22148
rect 17490 22092 17500 22148
rect 17556 22092 18508 22148
rect 18564 22092 18574 22148
rect 19282 22092 19292 22148
rect 19348 22092 19628 22148
rect 19684 22092 19694 22148
rect 20290 22092 20300 22148
rect 20356 22092 21644 22148
rect 21700 22092 21710 22148
rect 17500 22036 17556 22092
rect 16930 21980 16940 22036
rect 16996 21980 17556 22036
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 14242 21868 14252 21924
rect 14308 21868 15204 21924
rect 15148 21588 15204 21868
rect 15362 21756 15372 21812
rect 15428 21756 16156 21812
rect 16212 21756 16222 21812
rect 16370 21756 16380 21812
rect 16436 21756 20188 21812
rect 20244 21756 20254 21812
rect 25666 21756 25676 21812
rect 25732 21756 28140 21812
rect 28196 21756 28206 21812
rect 22194 21644 22204 21700
rect 22260 21644 23772 21700
rect 23828 21644 26572 21700
rect 26628 21644 26638 21700
rect 4274 21532 4284 21588
rect 4340 21532 9884 21588
rect 9940 21532 9950 21588
rect 11442 21532 11452 21588
rect 11508 21532 13468 21588
rect 13524 21532 13534 21588
rect 15138 21532 15148 21588
rect 15204 21532 15214 21588
rect 18498 21532 18508 21588
rect 18564 21532 20412 21588
rect 20468 21532 22652 21588
rect 22708 21532 22718 21588
rect 24434 21532 24444 21588
rect 24500 21532 25228 21588
rect 25284 21532 25294 21588
rect 16258 21420 16268 21476
rect 16324 21420 17388 21476
rect 17444 21420 17454 21476
rect 18386 21420 18396 21476
rect 18452 21420 19180 21476
rect 19236 21420 22540 21476
rect 22596 21420 23212 21476
rect 23268 21420 23278 21476
rect 23426 21420 23436 21476
rect 23492 21420 25788 21476
rect 25844 21420 29372 21476
rect 29428 21420 29438 21476
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 0 20916 800 20944
rect 0 20860 1932 20916
rect 1988 20860 1998 20916
rect 12114 20860 12124 20916
rect 12180 20860 12796 20916
rect 12852 20860 13356 20916
rect 13412 20860 14812 20916
rect 14868 20860 14878 20916
rect 0 20832 800 20860
rect 20066 20748 20076 20804
rect 20132 20748 21868 20804
rect 21924 20748 21934 20804
rect 31892 20748 37660 20804
rect 37716 20748 37726 20804
rect 9874 20636 9884 20692
rect 9940 20636 13468 20692
rect 13524 20636 13534 20692
rect 18162 20636 18172 20692
rect 18228 20636 20524 20692
rect 20580 20636 21420 20692
rect 21476 20636 21486 20692
rect 31892 20580 31948 20748
rect 29250 20524 29260 20580
rect 29316 20524 30828 20580
rect 30884 20524 31948 20580
rect 21522 20412 21532 20468
rect 21588 20412 22204 20468
rect 22260 20412 22270 20468
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 20402 20300 20412 20356
rect 20468 20300 20748 20356
rect 20804 20300 20814 20356
rect 41200 20244 42000 20272
rect 40002 20188 40012 20244
rect 40068 20188 42000 20244
rect 21970 20132 21980 20188
rect 22036 20132 22046 20188
rect 22754 20132 22764 20188
rect 22820 20132 22830 20188
rect 41200 20160 42000 20188
rect 10882 20076 10892 20132
rect 10948 20076 17500 20132
rect 17556 20076 19404 20132
rect 19460 20076 19470 20132
rect 19628 20076 20524 20132
rect 20580 20076 20590 20132
rect 21980 20076 26684 20132
rect 26740 20076 26750 20132
rect 19628 20020 19684 20076
rect 4274 19964 4284 20020
rect 4340 19964 9884 20020
rect 9940 19964 12460 20020
rect 12516 19964 12526 20020
rect 12674 19964 12684 20020
rect 12740 19964 13692 20020
rect 13748 19964 13758 20020
rect 14242 19964 14252 20020
rect 14308 19964 15596 20020
rect 15652 19964 17836 20020
rect 17892 19964 19684 20020
rect 19954 19964 19964 20020
rect 20020 19964 20636 20020
rect 20692 19964 20702 20020
rect 21858 19964 21868 20020
rect 21924 19964 23436 20020
rect 23492 19964 23502 20020
rect 24546 19964 24556 20020
rect 24612 19964 25228 20020
rect 25284 19964 25294 20020
rect 26898 19964 26908 20020
rect 26964 19964 28364 20020
rect 28420 19964 28430 20020
rect 12338 19852 12348 19908
rect 12404 19852 13132 19908
rect 13188 19852 13198 19908
rect 15138 19852 15148 19908
rect 15204 19852 16716 19908
rect 16772 19852 24668 19908
rect 24724 19852 24734 19908
rect 1922 19740 1932 19796
rect 1988 19740 1998 19796
rect 16594 19740 16604 19796
rect 16660 19740 18508 19796
rect 18564 19740 19964 19796
rect 20020 19740 20030 19796
rect 21746 19740 21756 19796
rect 21812 19740 23100 19796
rect 23156 19740 25116 19796
rect 25172 19740 25182 19796
rect 0 19572 800 19600
rect 1932 19572 1988 19740
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 41200 19572 42000 19600
rect 0 19516 1988 19572
rect 13346 19516 13356 19572
rect 13412 19516 15596 19572
rect 15652 19516 15662 19572
rect 40002 19516 40012 19572
rect 40068 19516 42000 19572
rect 0 19488 800 19516
rect 41200 19488 42000 19516
rect 20514 19292 20524 19348
rect 20580 19292 21308 19348
rect 21364 19292 21374 19348
rect 24546 19292 24556 19348
rect 24612 19292 24622 19348
rect 25666 19292 25676 19348
rect 25732 19292 28588 19348
rect 28644 19292 37660 19348
rect 37716 19292 37726 19348
rect 4274 19180 4284 19236
rect 4340 19180 12348 19236
rect 12404 19180 12414 19236
rect 16482 19180 16492 19236
rect 16548 19180 17500 19236
rect 17556 19180 19068 19236
rect 19124 19180 19516 19236
rect 19572 19180 21420 19236
rect 21476 19180 21486 19236
rect 22950 19180 22988 19236
rect 23044 19180 23054 19236
rect 24556 19124 24612 19292
rect 25778 19180 25788 19236
rect 25844 19180 27580 19236
rect 27636 19180 27646 19236
rect 28354 19180 28364 19236
rect 28420 19180 29596 19236
rect 29652 19180 29662 19236
rect 14354 19068 14364 19124
rect 14420 19068 15372 19124
rect 15428 19068 16268 19124
rect 16324 19068 16334 19124
rect 16818 19068 16828 19124
rect 16884 19068 17836 19124
rect 17892 19068 18844 19124
rect 18900 19068 19292 19124
rect 19348 19068 19358 19124
rect 19842 19068 19852 19124
rect 19908 19068 24612 19124
rect 14578 18956 14588 19012
rect 14644 18956 14654 19012
rect 15698 18956 15708 19012
rect 15764 18956 16044 19012
rect 16100 18956 17612 19012
rect 17668 18956 17678 19012
rect 17948 18956 18956 19012
rect 19012 18956 25004 19012
rect 25060 18956 25070 19012
rect 0 18900 800 18928
rect 14588 18900 14644 18956
rect 17948 18900 18004 18956
rect 0 18844 1932 18900
rect 1988 18844 1998 18900
rect 14588 18844 18004 18900
rect 23650 18844 23660 18900
rect 23716 18844 24332 18900
rect 24388 18844 26012 18900
rect 26068 18844 26078 18900
rect 0 18816 800 18844
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 21186 18732 21196 18788
rect 21252 18732 23100 18788
rect 23156 18732 24444 18788
rect 24500 18732 24510 18788
rect 18722 18620 18732 18676
rect 18788 18620 19628 18676
rect 19684 18620 19694 18676
rect 24098 18620 24108 18676
rect 24164 18620 29372 18676
rect 29428 18620 29438 18676
rect 14914 18508 14924 18564
rect 14980 18508 16940 18564
rect 16996 18508 18844 18564
rect 18900 18508 18910 18564
rect 22754 18508 22764 18564
rect 22820 18508 23996 18564
rect 24052 18508 24062 18564
rect 15810 18396 15820 18452
rect 15876 18396 17388 18452
rect 17444 18396 17724 18452
rect 17780 18396 17790 18452
rect 18610 18396 18620 18452
rect 18676 18396 21084 18452
rect 21140 18396 21980 18452
rect 22036 18396 22046 18452
rect 22978 18396 22988 18452
rect 23044 18396 23548 18452
rect 23604 18396 25676 18452
rect 25732 18396 25742 18452
rect 17154 18284 17164 18340
rect 17220 18284 18060 18340
rect 18116 18284 22652 18340
rect 22708 18284 23436 18340
rect 23492 18284 23884 18340
rect 23940 18284 23950 18340
rect 19282 18172 19292 18228
rect 19348 18172 20748 18228
rect 20804 18172 20814 18228
rect 20178 18060 20188 18116
rect 20244 18060 21644 18116
rect 21700 18060 22988 18116
rect 23044 18060 23054 18116
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 17714 17836 17724 17892
rect 17780 17836 19292 17892
rect 19348 17836 19358 17892
rect 17602 17724 17612 17780
rect 17668 17724 18956 17780
rect 19012 17724 22652 17780
rect 22708 17724 23660 17780
rect 23716 17724 23726 17780
rect 21634 17612 21644 17668
rect 21700 17612 22540 17668
rect 22596 17612 22606 17668
rect 27010 17612 27020 17668
rect 27076 17612 37660 17668
rect 37716 17612 37726 17668
rect 13794 17500 13804 17556
rect 13860 17500 17276 17556
rect 17332 17500 17342 17556
rect 17826 17500 17836 17556
rect 17892 17500 20748 17556
rect 20804 17500 21868 17556
rect 21924 17500 21934 17556
rect 22866 17500 22876 17556
rect 22932 17500 24444 17556
rect 24500 17500 24510 17556
rect 18162 17388 18172 17444
rect 18228 17388 19068 17444
rect 19124 17388 19134 17444
rect 21746 17388 21756 17444
rect 21812 17388 24220 17444
rect 24276 17388 24286 17444
rect 24546 17388 24556 17444
rect 24612 17388 25452 17444
rect 25508 17388 25518 17444
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 16034 17052 16044 17108
rect 16100 17052 19740 17108
rect 19796 17052 21196 17108
rect 21252 17052 21262 17108
rect 22530 17052 22540 17108
rect 22596 17052 23884 17108
rect 23940 17052 23950 17108
rect 24322 17052 24332 17108
rect 24388 17052 27020 17108
rect 27076 17052 27086 17108
rect 20514 16940 20524 16996
rect 20580 16940 22204 16996
rect 22260 16940 22270 16996
rect 25442 16940 25452 16996
rect 25508 16940 26684 16996
rect 26740 16940 26750 16996
rect 41200 16884 42000 16912
rect 13122 16828 13132 16884
rect 13188 16828 15372 16884
rect 15428 16828 16380 16884
rect 16436 16828 16446 16884
rect 40002 16828 40012 16884
rect 40068 16828 42000 16884
rect 41200 16800 42000 16828
rect 19170 16716 19180 16772
rect 19236 16716 19964 16772
rect 20020 16716 21308 16772
rect 21364 16716 21374 16772
rect 26002 16716 26012 16772
rect 26068 16716 27356 16772
rect 27412 16716 27422 16772
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 26450 16268 26460 16324
rect 26516 16268 27468 16324
rect 27524 16268 27534 16324
rect 41200 16212 42000 16240
rect 40002 16156 40012 16212
rect 40068 16156 42000 16212
rect 41200 16128 42000 16156
rect 26114 15820 26124 15876
rect 26180 15820 28028 15876
rect 28084 15820 28812 15876
rect 28868 15820 29260 15876
rect 29316 15820 29326 15876
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 16034 15484 16044 15540
rect 16100 15484 18620 15540
rect 18676 15484 21308 15540
rect 21364 15484 22540 15540
rect 22596 15484 23212 15540
rect 23268 15484 23278 15540
rect 22642 15260 22652 15316
rect 22708 15260 25228 15316
rect 25284 15260 25294 15316
rect 25442 15260 25452 15316
rect 25508 15260 25788 15316
rect 25844 15260 26236 15316
rect 26292 15260 26302 15316
rect 25452 15204 25508 15260
rect 21746 15148 21756 15204
rect 21812 15148 25508 15204
rect 27458 15148 27468 15204
rect 27524 15148 29036 15204
rect 29092 15148 37884 15204
rect 37940 15148 37950 15204
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 41200 14868 42000 14896
rect 40002 14812 40012 14868
rect 40068 14812 42000 14868
rect 41200 14784 42000 14812
rect 26898 14588 26908 14644
rect 26964 14588 28252 14644
rect 28308 14588 37660 14644
rect 37716 14588 37726 14644
rect 14018 14476 14028 14532
rect 14084 14476 15372 14532
rect 15428 14476 15438 14532
rect 25554 14476 25564 14532
rect 25620 14476 26684 14532
rect 26740 14476 26750 14532
rect 18274 14364 18284 14420
rect 18340 14364 18732 14420
rect 18788 14364 18798 14420
rect 19282 14364 19292 14420
rect 19348 14364 20636 14420
rect 20692 14364 21980 14420
rect 22036 14364 22046 14420
rect 22306 14364 22316 14420
rect 22372 14364 23548 14420
rect 23604 14364 23884 14420
rect 23940 14364 23950 14420
rect 14690 14252 14700 14308
rect 14756 14252 18620 14308
rect 18676 14252 18686 14308
rect 20066 14252 20076 14308
rect 20132 14252 20244 14308
rect 21074 14252 21084 14308
rect 21140 14252 21868 14308
rect 21924 14252 21934 14308
rect 23426 14252 23436 14308
rect 23492 14252 24220 14308
rect 24276 14252 25340 14308
rect 25396 14252 25406 14308
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 20188 13972 20244 14252
rect 15362 13916 15372 13972
rect 15428 13916 17500 13972
rect 17556 13916 18396 13972
rect 18452 13916 18462 13972
rect 20066 13916 20076 13972
rect 20132 13916 20244 13972
rect 19842 13804 19852 13860
rect 19908 13804 20748 13860
rect 20804 13804 20814 13860
rect 20402 13692 20412 13748
rect 20468 13692 22652 13748
rect 22708 13692 23436 13748
rect 23492 13692 23502 13748
rect 24098 13692 24108 13748
rect 24164 13692 25340 13748
rect 25396 13692 25406 13748
rect 18610 13468 18620 13524
rect 18676 13468 20188 13524
rect 20244 13468 20254 13524
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 41200 8820 42000 8848
rect 40226 8764 40236 8820
rect 40292 8764 42000 8820
rect 41200 8736 42000 8764
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 24882 4060 24892 4116
rect 24948 4060 26236 4116
rect 26292 4060 26302 4116
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 22866 3612 22876 3668
rect 22932 3612 25564 3668
rect 25620 3612 25630 3668
rect 23202 3500 23212 3556
rect 23268 3500 24556 3556
rect 24612 3500 24622 3556
rect 20178 3388 20188 3444
rect 20244 3388 21756 3444
rect 21812 3388 21822 3444
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
<< via3 >>
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 22988 19180 23044 19236
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 22988 18396 23044 18452
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
<< metal4 >>
rect 4448 38444 4768 38476
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 37660 20128 38476
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19808 34524 20128 36036
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 19808 23548 20128 25060
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 19808 21980 20128 23492
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 35168 38444 35488 38476
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 22988 19236 23044 19246
rect 22988 18452 23044 19180
rect 22988 18386 23044 18396
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _122_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17248 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _123_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 17024 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _124_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 17584 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _125_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 20272 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _126_
timestamp 1698175906
transform -1 0 18368 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _127_
timestamp 1698175906
transform -1 0 14448 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _128_
timestamp 1698175906
transform 1 0 12544 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _129_
timestamp 1698175906
transform 1 0 18928 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _130_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17360 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _131_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 16240 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _132_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 13328 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _133_
timestamp 1698175906
transform 1 0 18032 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _134_
timestamp 1698175906
transform -1 0 19264 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _135_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17696 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _136_
timestamp 1698175906
transform 1 0 16128 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _137_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18928 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _138_
timestamp 1698175906
transform -1 0 20832 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _139_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17024 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _140_
timestamp 1698175906
transform -1 0 15120 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _141_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 14112 0 1 20384
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _142_
timestamp 1698175906
transform 1 0 11312 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _143_
timestamp 1698175906
transform -1 0 19600 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _144_
timestamp 1698175906
transform -1 0 19152 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_2  _145_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19152 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _146_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 17024 0 -1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _147_
timestamp 1698175906
transform -1 0 24976 0 1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _148_
timestamp 1698175906
transform -1 0 16576 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _149_
timestamp 1698175906
transform -1 0 20944 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _150_
timestamp 1698175906
transform 1 0 20272 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _151_
timestamp 1698175906
transform 1 0 16688 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _152_
timestamp 1698175906
transform -1 0 18256 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _153_
timestamp 1698175906
transform 1 0 21840 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _154_
timestamp 1698175906
transform 1 0 19488 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _155_
timestamp 1698175906
transform 1 0 21392 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _156_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 23856 0 1 17248
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _157_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18368 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _158_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 18032 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _159_
timestamp 1698175906
transform -1 0 14448 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _160_
timestamp 1698175906
transform -1 0 13888 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _161_
timestamp 1698175906
transform 1 0 23184 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _162_
timestamp 1698175906
transform -1 0 27216 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _163_
timestamp 1698175906
transform 1 0 22064 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _164_
timestamp 1698175906
transform 1 0 21952 0 -1 15680
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _165_
timestamp 1698175906
transform 1 0 17696 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _166_
timestamp 1698175906
transform 1 0 21168 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _167_
timestamp 1698175906
transform 1 0 25088 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _168_
timestamp 1698175906
transform 1 0 27216 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _169_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21280 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _170_
timestamp 1698175906
transform -1 0 26768 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _171_
timestamp 1698175906
transform 1 0 23856 0 1 17248
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _172_
timestamp 1698175906
transform -1 0 26880 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _173_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 19264 0 -1 23520
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _174_
timestamp 1698175906
transform -1 0 19040 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _175_
timestamp 1698175906
transform -1 0 20272 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _176_
timestamp 1698175906
transform -1 0 17808 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _177_
timestamp 1698175906
transform 1 0 16016 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _178_
timestamp 1698175906
transform 1 0 19040 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _179_
timestamp 1698175906
transform 1 0 19936 0 1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _180_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 22176 0 -1 25088
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _181_
timestamp 1698175906
transform 1 0 17360 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _182_
timestamp 1698175906
transform 1 0 22960 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _183_
timestamp 1698175906
transform 1 0 25088 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _184_
timestamp 1698175906
transform -1 0 24304 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _185_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 20384 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _186_
timestamp 1698175906
transform -1 0 23072 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _187_
timestamp 1698175906
transform -1 0 21952 0 -1 15680
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _188_
timestamp 1698175906
transform 1 0 21616 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _189_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 22064 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _190_
timestamp 1698175906
transform 1 0 24080 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _191_
timestamp 1698175906
transform 1 0 25088 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _192_
timestamp 1698175906
transform 1 0 18368 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _193_
timestamp 1698175906
transform 1 0 19600 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _194_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 20160 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _195_
timestamp 1698175906
transform -1 0 20160 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _196_
timestamp 1698175906
transform -1 0 16016 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _197_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 15120 0 1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _198_
timestamp 1698175906
transform -1 0 12880 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _199_
timestamp 1698175906
transform 1 0 12880 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _200_
timestamp 1698175906
transform -1 0 20048 0 -1 23520
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _201_
timestamp 1698175906
transform -1 0 18368 0 1 23520
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _202_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 15568 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _203_
timestamp 1698175906
transform -1 0 15568 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _204_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 18256 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _205_
timestamp 1698175906
transform -1 0 18816 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _206_
timestamp 1698175906
transform 1 0 17248 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _207_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21168 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _208_
timestamp 1698175906
transform 1 0 25088 0 -1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _209_
timestamp 1698175906
transform 1 0 23856 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _210_
timestamp 1698175906
transform 1 0 26432 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _211_
timestamp 1698175906
transform 1 0 26208 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _212_
timestamp 1698175906
transform 1 0 19600 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _213_
timestamp 1698175906
transform 1 0 19936 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _214_
timestamp 1698175906
transform 1 0 18032 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _215_
timestamp 1698175906
transform 1 0 18368 0 1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _216_
timestamp 1698175906
transform 1 0 22512 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _217_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21280 0 1 18816
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _218_
timestamp 1698175906
transform 1 0 23856 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _219_
timestamp 1698175906
transform 1 0 22512 0 -1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _220_
timestamp 1698175906
transform -1 0 29680 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _221_
timestamp 1698175906
transform -1 0 29568 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _222_
timestamp 1698175906
transform 1 0 29008 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _223_
timestamp 1698175906
transform -1 0 25760 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _224_
timestamp 1698175906
transform -1 0 24752 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _225_
timestamp 1698175906
transform 1 0 25088 0 -1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _226_
timestamp 1698175906
transform 1 0 25760 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _227_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 23968 0 1 21952
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai222_2  _228_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 24192 0 1 25088
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _229_
timestamp 1698175906
transform 1 0 23072 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _230_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21728 0 1 23520
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _231_
timestamp 1698175906
transform -1 0 29568 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _232_
timestamp 1698175906
transform 1 0 29008 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _233_
timestamp 1698175906
transform 1 0 29680 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _234_
timestamp 1698175906
transform 1 0 22736 0 -1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _235_
timestamp 1698175906
transform 1 0 28112 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _236_
timestamp 1698175906
transform -1 0 27328 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _237_
timestamp 1698175906
transform 1 0 22512 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _238_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21280 0 1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _239_
timestamp 1698175906
transform 1 0 21392 0 -1 23520
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _240_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 25088 0 -1 26656
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _241_
timestamp 1698175906
transform -1 0 22960 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _242_
timestamp 1698175906
transform -1 0 26880 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _243_
timestamp 1698175906
transform -1 0 25872 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _244_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 13104 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _245_
timestamp 1698175906
transform -1 0 12992 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _246_
timestamp 1698175906
transform 1 0 15120 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _247_
timestamp 1698175906
transform 1 0 13440 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _248_
timestamp 1698175906
transform 1 0 12880 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _249_
timestamp 1698175906
transform 1 0 11872 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _250_
timestamp 1698175906
transform 1 0 25200 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _251_
timestamp 1698175906
transform 1 0 25984 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _252_
timestamp 1698175906
transform 1 0 14112 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _253_
timestamp 1698175906
transform 1 0 22512 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _254_
timestamp 1698175906
transform 1 0 20160 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _255_
timestamp 1698175906
transform 1 0 23968 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _256_
timestamp 1698175906
transform 1 0 18256 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _257_
timestamp 1698175906
transform -1 0 12992 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _258_
timestamp 1698175906
transform -1 0 16128 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _259_
timestamp 1698175906
transform 1 0 13776 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _260_
timestamp 1698175906
transform 1 0 25536 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _261_
timestamp 1698175906
transform 1 0 17696 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _262_
timestamp 1698175906
transform 1 0 13776 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _263_
timestamp 1698175906
transform 1 0 27776 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _264_
timestamp 1698175906
transform 1 0 25088 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _265_
timestamp 1698175906
transform 1 0 21168 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _266_
timestamp 1698175906
transform 1 0 27552 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _267_
timestamp 1698175906
transform 1 0 27776 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _268_
timestamp 1698175906
transform 1 0 24640 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _269_
timestamp 1698175906
transform 1 0 25088 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _272_
timestamp 1698175906
transform -1 0 12880 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _273_
timestamp 1698175906
transform 1 0 16800 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__141__A3 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 14560 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__208__A1
timestamp 1698175906
transform 1 0 24976 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__212__A2
timestamp 1698175906
transform -1 0 19600 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__215__A2
timestamp 1698175906
transform -1 0 18928 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__244__CLK
timestamp 1698175906
transform 1 0 13328 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__245__CLK
timestamp 1698175906
transform 1 0 14784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__246__CLK
timestamp 1698175906
transform 1 0 18368 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__247__CLK
timestamp 1698175906
transform 1 0 16688 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__248__CLK
timestamp 1698175906
transform 1 0 16352 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__249__CLK
timestamp 1698175906
transform 1 0 15344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__250__CLK
timestamp 1698175906
transform 1 0 29232 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__251__CLK
timestamp 1698175906
transform 1 0 29456 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__252__CLK
timestamp 1698175906
transform 1 0 19040 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__253__CLK
timestamp 1698175906
transform -1 0 26208 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__254__CLK
timestamp 1698175906
transform 1 0 23408 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__255__CLK
timestamp 1698175906
transform 1 0 28000 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__256__CLK
timestamp 1698175906
transform 1 0 18032 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__257__CLK
timestamp 1698175906
transform 1 0 13552 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__258__CLK
timestamp 1698175906
transform 1 0 16352 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__259__CLK
timestamp 1698175906
transform -1 0 17696 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__260__CLK
timestamp 1698175906
transform 1 0 28784 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__261__CLK
timestamp 1698175906
transform -1 0 17696 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__262__CLK
timestamp 1698175906
transform 1 0 17472 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__263__CLK
timestamp 1698175906
transform 1 0 27552 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__264__CLK
timestamp 1698175906
transform 1 0 28560 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__265__CLK
timestamp 1698175906
transform 1 0 24416 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__266__CLK
timestamp 1698175906
transform 1 0 27328 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__267__CLK
timestamp 1698175906
transform 1 0 27552 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__268__CLK
timestamp 1698175906
transform 1 0 28112 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__269__CLK
timestamp 1698175906
transform -1 0 28784 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1698175906
transform 1 0 17472 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19264 0 -1 20384
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1698175906
transform -1 0 20944 0 1 20384
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1698175906
transform 1 0 23184 0 1 20384
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1568 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698175906
transform 1 0 5376 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698175906
transform 1 0 9184 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698175906
transform 1 0 12992 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_138 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 16800 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_142 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17248 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_198
timestamp 1698175906
transform 1 0 23520 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_202
timestamp 1698175906
transform 1 0 23968 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_232
timestamp 1698175906
transform 1 0 27328 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_236
timestamp 1698175906
transform 1 0 27776 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_240
timestamp 1698175906
transform 1 0 28224 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_274
timestamp 1698175906
transform 1 0 32032 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_308
timestamp 1698175906
transform 1 0 35840 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_342
timestamp 1698175906
transform 1 0 39648 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_346
timestamp 1698175906
transform 1 0 40096 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_348 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 40320 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1568 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698175906
transform 1 0 8736 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698175906
transform 1 0 9408 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698175906
transform 1 0 16576 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_142
timestamp 1698175906
transform 1 0 17248 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_206
timestamp 1698175906
transform 1 0 24416 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_238
timestamp 1698175906
transform 1 0 28000 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_270 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 31584 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_278
timestamp 1698175906
transform 1 0 32480 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_282
timestamp 1698175906
transform 1 0 32928 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_346
timestamp 1698175906
transform 1 0 40096 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_348
timestamp 1698175906
transform 1 0 40320 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698175906
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698175906
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698175906
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698175906
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_107
timestamp 1698175906
transform 1 0 13328 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_171
timestamp 1698175906
transform 1 0 20496 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_177
timestamp 1698175906
transform 1 0 21168 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_241
timestamp 1698175906
transform 1 0 28336 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698175906
transform 1 0 29008 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698175906
transform 1 0 36176 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_317
timestamp 1698175906
transform 1 0 36848 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698175906
transform 1 0 1568 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698175906
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698175906
transform 1 0 9408 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698175906
transform 1 0 16576 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_142
timestamp 1698175906
transform 1 0 17248 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_206
timestamp 1698175906
transform 1 0 24416 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_212
timestamp 1698175906
transform 1 0 25088 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_276
timestamp 1698175906
transform 1 0 32256 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_282
timestamp 1698175906
transform 1 0 32928 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_346
timestamp 1698175906
transform 1 0 40096 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_348
timestamp 1698175906
transform 1 0 40320 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698175906
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698175906
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698175906
transform 1 0 5488 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698175906
transform 1 0 12656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_107
timestamp 1698175906
transform 1 0 13328 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698175906
transform 1 0 20496 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_177
timestamp 1698175906
transform 1 0 21168 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_241
timestamp 1698175906
transform 1 0 28336 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698175906
transform 1 0 29008 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698175906
transform 1 0 36176 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_317
timestamp 1698175906
transform 1 0 36848 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698175906
transform 1 0 1568 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698175906
transform 1 0 8736 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698175906
transform 1 0 9408 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698175906
transform 1 0 16576 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_142
timestamp 1698175906
transform 1 0 17248 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_206
timestamp 1698175906
transform 1 0 24416 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_212
timestamp 1698175906
transform 1 0 25088 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698175906
transform 1 0 32256 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_282
timestamp 1698175906
transform 1 0 32928 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_346
timestamp 1698175906
transform 1 0 40096 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_348
timestamp 1698175906
transform 1 0 40320 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698175906
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698175906
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698175906
transform 1 0 5488 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698175906
transform 1 0 12656 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_107
timestamp 1698175906
transform 1 0 13328 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_171
timestamp 1698175906
transform 1 0 20496 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_177
timestamp 1698175906
transform 1 0 21168 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_241
timestamp 1698175906
transform 1 0 28336 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_247
timestamp 1698175906
transform 1 0 29008 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_311
timestamp 1698175906
transform 1 0 36176 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_317
timestamp 1698175906
transform 1 0 36848 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698175906
transform 1 0 1568 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698175906
transform 1 0 8736 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_72
timestamp 1698175906
transform 1 0 9408 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698175906
transform 1 0 16576 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_142
timestamp 1698175906
transform 1 0 17248 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_206
timestamp 1698175906
transform 1 0 24416 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_212
timestamp 1698175906
transform 1 0 25088 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_276
timestamp 1698175906
transform 1 0 32256 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_7_282
timestamp 1698175906
transform 1 0 32928 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_314 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 36512 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_330
timestamp 1698175906
transform 1 0 38304 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_338
timestamp 1698175906
transform 1 0 39200 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_342
timestamp 1698175906
transform 1 0 39648 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_344
timestamp 1698175906
transform 1 0 39872 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698175906
transform 1 0 1568 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698175906
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_37
timestamp 1698175906
transform 1 0 5488 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_101
timestamp 1698175906
transform 1 0 12656 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_107
timestamp 1698175906
transform 1 0 13328 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_171
timestamp 1698175906
transform 1 0 20496 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_177
timestamp 1698175906
transform 1 0 21168 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_241
timestamp 1698175906
transform 1 0 28336 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_247
timestamp 1698175906
transform 1 0 29008 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_311
timestamp 1698175906
transform 1 0 36176 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_317
timestamp 1698175906
transform 1 0 36848 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698175906
transform 1 0 1568 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698175906
transform 1 0 8736 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_72
timestamp 1698175906
transform 1 0 9408 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_136
timestamp 1698175906
transform 1 0 16576 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_142
timestamp 1698175906
transform 1 0 17248 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_206
timestamp 1698175906
transform 1 0 24416 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_212
timestamp 1698175906
transform 1 0 25088 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_276
timestamp 1698175906
transform 1 0 32256 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_282
timestamp 1698175906
transform 1 0 32928 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_346
timestamp 1698175906
transform 1 0 40096 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_348
timestamp 1698175906
transform 1 0 40320 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698175906
transform 1 0 1568 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698175906
transform 1 0 5152 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_37
timestamp 1698175906
transform 1 0 5488 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698175906
transform 1 0 12656 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_107
timestamp 1698175906
transform 1 0 13328 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_171
timestamp 1698175906
transform 1 0 20496 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_177
timestamp 1698175906
transform 1 0 21168 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_241
timestamp 1698175906
transform 1 0 28336 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_247
timestamp 1698175906
transform 1 0 29008 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_311
timestamp 1698175906
transform 1 0 36176 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_317
timestamp 1698175906
transform 1 0 36848 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2
timestamp 1698175906
transform 1 0 1568 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698175906
transform 1 0 8736 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_72
timestamp 1698175906
transform 1 0 9408 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698175906
transform 1 0 16576 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_142
timestamp 1698175906
transform 1 0 17248 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_206
timestamp 1698175906
transform 1 0 24416 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_212
timestamp 1698175906
transform 1 0 25088 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_276
timestamp 1698175906
transform 1 0 32256 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_282
timestamp 1698175906
transform 1 0 32928 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_346
timestamp 1698175906
transform 1 0 40096 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_348
timestamp 1698175906
transform 1 0 40320 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698175906
transform 1 0 1568 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698175906
transform 1 0 5152 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_37
timestamp 1698175906
transform 1 0 5488 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698175906
transform 1 0 12656 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_107
timestamp 1698175906
transform 1 0 13328 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_139
timestamp 1698175906
transform 1 0 16912 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_143
timestamp 1698175906
transform 1 0 17360 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_177
timestamp 1698175906
transform 1 0 21168 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_185
timestamp 1698175906
transform 1 0 22064 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_218
timestamp 1698175906
transform 1 0 25760 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_222
timestamp 1698175906
transform 1 0 26208 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_238
timestamp 1698175906
transform 1 0 28000 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_242
timestamp 1698175906
transform 1 0 28448 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_244
timestamp 1698175906
transform 1 0 28672 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_247
timestamp 1698175906
transform 1 0 29008 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_311
timestamp 1698175906
transform 1 0 36176 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_317
timestamp 1698175906
transform 1 0 36848 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_2
timestamp 1698175906
transform 1 0 1568 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_66
timestamp 1698175906
transform 1 0 8736 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_72
timestamp 1698175906
transform 1 0 9408 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_104
timestamp 1698175906
transform 1 0 12992 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_108
timestamp 1698175906
transform 1 0 13440 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_110
timestamp 1698175906
transform 1 0 13664 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_142
timestamp 1698175906
transform 1 0 17248 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_146
timestamp 1698175906
transform 1 0 17696 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_148
timestamp 1698175906
transform 1 0 17920 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_153
timestamp 1698175906
transform 1 0 18480 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_157
timestamp 1698175906
transform 1 0 18928 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_205
timestamp 1698175906
transform 1 0 24304 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_209
timestamp 1698175906
transform 1 0 24752 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_218
timestamp 1698175906
transform 1 0 25760 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_231
timestamp 1698175906
transform 1 0 27216 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_263
timestamp 1698175906
transform 1 0 30800 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_279
timestamp 1698175906
transform 1 0 32592 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_282
timestamp 1698175906
transform 1 0 32928 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_346
timestamp 1698175906
transform 1 0 40096 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_348
timestamp 1698175906
transform 1 0 40320 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698175906
transform 1 0 1568 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698175906
transform 1 0 5152 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_37
timestamp 1698175906
transform 1 0 5488 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_101
timestamp 1698175906
transform 1 0 12656 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_107
timestamp 1698175906
transform 1 0 13328 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_162
timestamp 1698175906
transform 1 0 19488 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_174
timestamp 1698175906
transform 1 0 20832 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_177
timestamp 1698175906
transform 1 0 21168 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_194
timestamp 1698175906
transform 1 0 23072 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_196
timestamp 1698175906
transform 1 0 23296 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_199
timestamp 1698175906
transform 1 0 23632 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_207
timestamp 1698175906
transform 1 0 24528 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_211
timestamp 1698175906
transform 1 0 24976 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_242
timestamp 1698175906
transform 1 0 28448 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_244
timestamp 1698175906
transform 1 0 28672 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_247
timestamp 1698175906
transform 1 0 29008 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_251
timestamp 1698175906
transform 1 0 29456 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_317
timestamp 1698175906
transform 1 0 36848 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_2
timestamp 1698175906
transform 1 0 1568 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_66
timestamp 1698175906
transform 1 0 8736 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_72
timestamp 1698175906
transform 1 0 9408 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_136
timestamp 1698175906
transform 1 0 16576 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_142
timestamp 1698175906
transform 1 0 17248 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_150
timestamp 1698175906
transform 1 0 18144 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_154
timestamp 1698175906
transform 1 0 18592 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_170
timestamp 1698175906
transform 1 0 20384 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_174
timestamp 1698175906
transform 1 0 20832 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_176
timestamp 1698175906
transform 1 0 21056 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_191
timestamp 1698175906
transform 1 0 22736 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_207
timestamp 1698175906
transform 1 0 24528 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_209
timestamp 1698175906
transform 1 0 24752 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_249
timestamp 1698175906
transform 1 0 29232 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_253
timestamp 1698175906
transform 1 0 29680 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_269
timestamp 1698175906
transform 1 0 31472 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_277
timestamp 1698175906
transform 1 0 32368 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_279
timestamp 1698175906
transform 1 0 32592 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_282
timestamp 1698175906
transform 1 0 32928 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_314
timestamp 1698175906
transform 1 0 36512 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_322
timestamp 1698175906
transform 1 0 37408 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_2
timestamp 1698175906
transform 1 0 1568 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698175906
transform 1 0 5152 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_37
timestamp 1698175906
transform 1 0 5488 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_101
timestamp 1698175906
transform 1 0 12656 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_107
timestamp 1698175906
transform 1 0 13328 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_171
timestamp 1698175906
transform 1 0 20496 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_183
timestamp 1698175906
transform 1 0 21840 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_199
timestamp 1698175906
transform 1 0 23632 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_201
timestamp 1698175906
transform 1 0 23856 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_236
timestamp 1698175906
transform 1 0 27776 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_240
timestamp 1698175906
transform 1 0 28224 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_244
timestamp 1698175906
transform 1 0 28672 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_247
timestamp 1698175906
transform 1 0 29008 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_311
timestamp 1698175906
transform 1 0 36176 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_317
timestamp 1698175906
transform 1 0 36848 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_2
timestamp 1698175906
transform 1 0 1568 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_66
timestamp 1698175906
transform 1 0 8736 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_72
timestamp 1698175906
transform 1 0 9408 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_88
timestamp 1698175906
transform 1 0 11200 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_96
timestamp 1698175906
transform 1 0 12096 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_100
timestamp 1698175906
transform 1 0 12544 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_102
timestamp 1698175906
transform 1 0 12768 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_132
timestamp 1698175906
transform 1 0 16128 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_136
timestamp 1698175906
transform 1 0 16576 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_142
timestamp 1698175906
transform 1 0 17248 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_158
timestamp 1698175906
transform 1 0 19040 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_162
timestamp 1698175906
transform 1 0 19488 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_169
timestamp 1698175906
transform 1 0 20272 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_177
timestamp 1698175906
transform 1 0 21168 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_191
timestamp 1698175906
transform 1 0 22736 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_199
timestamp 1698175906
transform 1 0 23632 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_208
timestamp 1698175906
transform 1 0 24640 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_228
timestamp 1698175906
transform 1 0 26880 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_260
timestamp 1698175906
transform 1 0 30464 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_276
timestamp 1698175906
transform 1 0 32256 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_282
timestamp 1698175906
transform 1 0 32928 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_314
timestamp 1698175906
transform 1 0 36512 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_322
timestamp 1698175906
transform 1 0 37408 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_2
timestamp 1698175906
transform 1 0 1568 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698175906
transform 1 0 5152 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_37
timestamp 1698175906
transform 1 0 5488 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_101
timestamp 1698175906
transform 1 0 12656 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_107
timestamp 1698175906
transform 1 0 13328 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_123
timestamp 1698175906
transform 1 0 15120 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_131
timestamp 1698175906
transform 1 0 16016 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_135
timestamp 1698175906
transform 1 0 16464 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_139
timestamp 1698175906
transform 1 0 16912 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_165
timestamp 1698175906
transform 1 0 19824 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_185
timestamp 1698175906
transform 1 0 22064 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_187
timestamp 1698175906
transform 1 0 22288 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_208
timestamp 1698175906
transform 1 0 24640 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_240
timestamp 1698175906
transform 1 0 28224 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_244
timestamp 1698175906
transform 1 0 28672 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_247
timestamp 1698175906
transform 1 0 29008 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_311
timestamp 1698175906
transform 1 0 36176 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_317
timestamp 1698175906
transform 1 0 36848 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_321
timestamp 1698175906
transform 1 0 37296 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_2
timestamp 1698175906
transform 1 0 1568 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_66
timestamp 1698175906
transform 1 0 8736 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_72
timestamp 1698175906
transform 1 0 9408 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_88
timestamp 1698175906
transform 1 0 11200 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_96
timestamp 1698175906
transform 1 0 12096 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_103
timestamp 1698175906
transform 1 0 12880 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_107
timestamp 1698175906
transform 1 0 13328 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_137
timestamp 1698175906
transform 1 0 16688 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_139
timestamp 1698175906
transform 1 0 16912 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_142
timestamp 1698175906
transform 1 0 17248 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_144
timestamp 1698175906
transform 1 0 17472 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_151
timestamp 1698175906
transform 1 0 18256 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_182
timestamp 1698175906
transform 1 0 21728 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_209
timestamp 1698175906
transform 1 0 24752 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_212
timestamp 1698175906
transform 1 0 25088 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_244
timestamp 1698175906
transform 1 0 28672 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_247
timestamp 1698175906
transform 1 0 29008 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_279
timestamp 1698175906
transform 1 0 32592 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_282
timestamp 1698175906
transform 1 0 32928 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_346
timestamp 1698175906
transform 1 0 40096 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_348
timestamp 1698175906
transform 1 0 40320 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_28
timestamp 1698175906
transform 1 0 4480 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_32
timestamp 1698175906
transform 1 0 4928 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698175906
transform 1 0 5152 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_37
timestamp 1698175906
transform 1 0 5488 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_69
timestamp 1698175906
transform 1 0 9072 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_73
timestamp 1698175906
transform 1 0 9520 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_104
timestamp 1698175906
transform 1 0 12992 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_107
timestamp 1698175906
transform 1 0 13328 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_111
timestamp 1698175906
transform 1 0 13776 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_115
timestamp 1698175906
transform 1 0 14224 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_136
timestamp 1698175906
transform 1 0 16576 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_177
timestamp 1698175906
transform 1 0 21168 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_197
timestamp 1698175906
transform 1 0 23408 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_209
timestamp 1698175906
transform 1 0 24752 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_213
timestamp 1698175906
transform 1 0 25200 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_215
timestamp 1698175906
transform 1 0 25424 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_255
timestamp 1698175906
transform 1 0 29904 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_287
timestamp 1698175906
transform 1 0 33488 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_303
timestamp 1698175906
transform 1 0 35280 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_311
timestamp 1698175906
transform 1 0 36176 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_317
timestamp 1698175906
transform 1 0 36848 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_28
timestamp 1698175906
transform 1 0 4480 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_60
timestamp 1698175906
transform 1 0 8064 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_68
timestamp 1698175906
transform 1 0 8960 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_72
timestamp 1698175906
transform 1 0 9408 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_88
timestamp 1698175906
transform 1 0 11200 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_96
timestamp 1698175906
transform 1 0 12096 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_117
timestamp 1698175906
transform 1 0 14448 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_142
timestamp 1698175906
transform 1 0 17248 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_230
timestamp 1698175906
transform 1 0 27104 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_265
timestamp 1698175906
transform 1 0 31024 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_273
timestamp 1698175906
transform 1 0 31920 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_277
timestamp 1698175906
transform 1 0 32368 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_279
timestamp 1698175906
transform 1 0 32592 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_282
timestamp 1698175906
transform 1 0 32928 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_314
timestamp 1698175906
transform 1 0 36512 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_322
timestamp 1698175906
transform 1 0 37408 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_2
timestamp 1698175906
transform 1 0 1568 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698175906
transform 1 0 5152 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_37
timestamp 1698175906
transform 1 0 5488 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_69
timestamp 1698175906
transform 1 0 9072 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_73
timestamp 1698175906
transform 1 0 9520 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_104
timestamp 1698175906
transform 1 0 12992 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_114
timestamp 1698175906
transform 1 0 14112 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_118
timestamp 1698175906
transform 1 0 14560 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_122
timestamp 1698175906
transform 1 0 15008 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_124
timestamp 1698175906
transform 1 0 15232 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_193
timestamp 1698175906
transform 1 0 22960 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_252
timestamp 1698175906
transform 1 0 29568 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_284
timestamp 1698175906
transform 1 0 33152 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_300
timestamp 1698175906
transform 1 0 34944 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_308
timestamp 1698175906
transform 1 0 35840 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_312
timestamp 1698175906
transform 1 0 36288 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_314
timestamp 1698175906
transform 1 0 36512 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_317
timestamp 1698175906
transform 1 0 36848 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_321
timestamp 1698175906
transform 1 0 37296 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_28
timestamp 1698175906
transform 1 0 4480 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_60
timestamp 1698175906
transform 1 0 8064 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_68
timestamp 1698175906
transform 1 0 8960 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_72
timestamp 1698175906
transform 1 0 9408 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_88
timestamp 1698175906
transform 1 0 11200 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_123
timestamp 1698175906
transform 1 0 15120 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_127
timestamp 1698175906
transform 1 0 15568 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_131
timestamp 1698175906
transform 1 0 16016 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_154
timestamp 1698175906
transform 1 0 18592 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_156
timestamp 1698175906
transform 1 0 18816 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_202
timestamp 1698175906
transform 1 0 23968 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_227
timestamp 1698175906
transform 1 0 26768 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_231
timestamp 1698175906
transform 1 0 27216 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_233
timestamp 1698175906
transform 1 0 27440 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_265
timestamp 1698175906
transform 1 0 31024 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_273
timestamp 1698175906
transform 1 0 31920 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_277
timestamp 1698175906
transform 1 0 32368 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_279
timestamp 1698175906
transform 1 0 32592 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_282
timestamp 1698175906
transform 1 0 32928 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_346
timestamp 1698175906
transform 1 0 40096 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_348
timestamp 1698175906
transform 1 0 40320 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_2
timestamp 1698175906
transform 1 0 1568 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698175906
transform 1 0 5152 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_37
timestamp 1698175906
transform 1 0 5488 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_101
timestamp 1698175906
transform 1 0 12656 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_117
timestamp 1698175906
transform 1 0 14448 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_133
timestamp 1698175906
transform 1 0 16240 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_177
timestamp 1698175906
transform 1 0 21168 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_211
timestamp 1698175906
transform 1 0 24976 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_241
timestamp 1698175906
transform 1 0 28336 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_258
timestamp 1698175906
transform 1 0 30240 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_290
timestamp 1698175906
transform 1 0 33824 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_306
timestamp 1698175906
transform 1 0 35616 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_314
timestamp 1698175906
transform 1 0 36512 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_317
timestamp 1698175906
transform 1 0 36848 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_321
timestamp 1698175906
transform 1 0 37296 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_2
timestamp 1698175906
transform 1 0 1568 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_66
timestamp 1698175906
transform 1 0 8736 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_72
timestamp 1698175906
transform 1 0 9408 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_88
timestamp 1698175906
transform 1 0 11200 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_96
timestamp 1698175906
transform 1 0 12096 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_105
timestamp 1698175906
transform 1 0 13104 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_109
timestamp 1698175906
transform 1 0 13552 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_125
timestamp 1698175906
transform 1 0 15344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_133
timestamp 1698175906
transform 1 0 16240 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_137
timestamp 1698175906
transform 1 0 16688 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_139
timestamp 1698175906
transform 1 0 16912 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_142
timestamp 1698175906
transform 1 0 17248 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_146
timestamp 1698175906
transform 1 0 17696 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_167
timestamp 1698175906
transform 1 0 20048 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_175
timestamp 1698175906
transform 1 0 20944 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_190
timestamp 1698175906
transform 1 0 22624 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_207
timestamp 1698175906
transform 1 0 24528 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_209
timestamp 1698175906
transform 1 0 24752 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_230
timestamp 1698175906
transform 1 0 27104 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_238
timestamp 1698175906
transform 1 0 28000 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_247
timestamp 1698175906
transform 1 0 29008 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_279
timestamp 1698175906
transform 1 0 32592 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_282
timestamp 1698175906
transform 1 0 32928 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_314
timestamp 1698175906
transform 1 0 36512 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_322
timestamp 1698175906
transform 1 0 37408 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_28
timestamp 1698175906
transform 1 0 4480 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_32
timestamp 1698175906
transform 1 0 4928 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698175906
transform 1 0 5152 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_37
timestamp 1698175906
transform 1 0 5488 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_69
timestamp 1698175906
transform 1 0 9072 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_73
timestamp 1698175906
transform 1 0 9520 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_75
timestamp 1698175906
transform 1 0 9744 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_115
timestamp 1698175906
transform 1 0 14224 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_152
timestamp 1698175906
transform 1 0 18368 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_156
timestamp 1698175906
transform 1 0 18816 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_158
timestamp 1698175906
transform 1 0 19040 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_163
timestamp 1698175906
transform 1 0 19600 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_167
timestamp 1698175906
transform 1 0 20048 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_174
timestamp 1698175906
transform 1 0 20832 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_177
timestamp 1698175906
transform 1 0 21168 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_181
timestamp 1698175906
transform 1 0 21616 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_198
timestamp 1698175906
transform 1 0 23520 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_230
timestamp 1698175906
transform 1 0 27104 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_238
timestamp 1698175906
transform 1 0 28000 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_242
timestamp 1698175906
transform 1 0 28448 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_244
timestamp 1698175906
transform 1 0 28672 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_255
timestamp 1698175906
transform 1 0 29904 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_287
timestamp 1698175906
transform 1 0 33488 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_303
timestamp 1698175906
transform 1 0 35280 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_311
timestamp 1698175906
transform 1 0 36176 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_317
timestamp 1698175906
transform 1 0 36848 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_28
timestamp 1698175906
transform 1 0 4480 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_60
timestamp 1698175906
transform 1 0 8064 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_68
timestamp 1698175906
transform 1 0 8960 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_72
timestamp 1698175906
transform 1 0 9408 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_88
timestamp 1698175906
transform 1 0 11200 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_96
timestamp 1698175906
transform 1 0 12096 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_100
timestamp 1698175906
transform 1 0 12544 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_102
timestamp 1698175906
transform 1 0 12768 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_132
timestamp 1698175906
transform 1 0 16128 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_136
timestamp 1698175906
transform 1 0 16576 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_147
timestamp 1698175906
transform 1 0 17808 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_186
timestamp 1698175906
transform 1 0 22176 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_188
timestamp 1698175906
transform 1 0 22400 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_197
timestamp 1698175906
transform 1 0 23408 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_205
timestamp 1698175906
transform 1 0 24304 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_209
timestamp 1698175906
transform 1 0 24752 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_212
timestamp 1698175906
transform 1 0 25088 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_228
timestamp 1698175906
transform 1 0 26880 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_263
timestamp 1698175906
transform 1 0 30800 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_279
timestamp 1698175906
transform 1 0 32592 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_282
timestamp 1698175906
transform 1 0 32928 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_346
timestamp 1698175906
transform 1 0 40096 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_348
timestamp 1698175906
transform 1 0 40320 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_2
timestamp 1698175906
transform 1 0 1568 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698175906
transform 1 0 5152 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_37
timestamp 1698175906
transform 1 0 5488 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_101
timestamp 1698175906
transform 1 0 12656 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_107
timestamp 1698175906
transform 1 0 13328 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_171
timestamp 1698175906
transform 1 0 20496 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_204
timestamp 1698175906
transform 1 0 24192 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_208
timestamp 1698175906
transform 1 0 24640 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_210
timestamp 1698175906
transform 1 0 24864 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_219
timestamp 1698175906
transform 1 0 25872 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_235
timestamp 1698175906
transform 1 0 27664 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_243
timestamp 1698175906
transform 1 0 28560 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_252
timestamp 1698175906
transform 1 0 29568 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_284
timestamp 1698175906
transform 1 0 33152 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_300
timestamp 1698175906
transform 1 0 34944 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_308
timestamp 1698175906
transform 1 0 35840 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_312
timestamp 1698175906
transform 1 0 36288 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_314
timestamp 1698175906
transform 1 0 36512 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_317
timestamp 1698175906
transform 1 0 36848 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_321
timestamp 1698175906
transform 1 0 37296 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_2
timestamp 1698175906
transform 1 0 1568 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_66
timestamp 1698175906
transform 1 0 8736 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_72
timestamp 1698175906
transform 1 0 9408 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_136
timestamp 1698175906
transform 1 0 16576 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_142
timestamp 1698175906
transform 1 0 17248 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_151
timestamp 1698175906
transform 1 0 18256 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_158
timestamp 1698175906
transform 1 0 19040 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_166
timestamp 1698175906
transform 1 0 19936 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_178
timestamp 1698175906
transform 1 0 21280 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_186
timestamp 1698175906
transform 1 0 22176 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_193
timestamp 1698175906
transform 1 0 22960 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_200
timestamp 1698175906
transform 1 0 23744 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_204
timestamp 1698175906
transform 1 0 24192 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_208
timestamp 1698175906
transform 1 0 24640 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_232
timestamp 1698175906
transform 1 0 27328 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_264
timestamp 1698175906
transform 1 0 30912 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_282
timestamp 1698175906
transform 1 0 32928 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_346
timestamp 1698175906
transform 1 0 40096 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_348
timestamp 1698175906
transform 1 0 40320 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_2
timestamp 1698175906
transform 1 0 1568 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698175906
transform 1 0 5152 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_37
timestamp 1698175906
transform 1 0 5488 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_101
timestamp 1698175906
transform 1 0 12656 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_107
timestamp 1698175906
transform 1 0 13328 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_111
timestamp 1698175906
transform 1 0 13776 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_113
timestamp 1698175906
transform 1 0 14000 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_156
timestamp 1698175906
transform 1 0 18816 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_160
timestamp 1698175906
transform 1 0 19264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_168
timestamp 1698175906
transform 1 0 20160 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_172
timestamp 1698175906
transform 1 0 20608 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_174
timestamp 1698175906
transform 1 0 20832 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_206
timestamp 1698175906
transform 1 0 24416 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_237
timestamp 1698175906
transform 1 0 27888 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_241
timestamp 1698175906
transform 1 0 28336 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_247
timestamp 1698175906
transform 1 0 29008 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_311
timestamp 1698175906
transform 1 0 36176 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_317
timestamp 1698175906
transform 1 0 36848 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_321
timestamp 1698175906
transform 1 0 37296 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_2
timestamp 1698175906
transform 1 0 1568 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_66
timestamp 1698175906
transform 1 0 8736 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_72
timestamp 1698175906
transform 1 0 9408 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_104
timestamp 1698175906
transform 1 0 12992 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_108
timestamp 1698175906
transform 1 0 13440 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_110
timestamp 1698175906
transform 1 0 13664 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_150
timestamp 1698175906
transform 1 0 18144 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_180
timestamp 1698175906
transform 1 0 21504 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_196
timestamp 1698175906
transform 1 0 23296 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_204
timestamp 1698175906
transform 1 0 24192 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_208
timestamp 1698175906
transform 1 0 24640 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_241
timestamp 1698175906
transform 1 0 28336 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_245
timestamp 1698175906
transform 1 0 28784 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_277
timestamp 1698175906
transform 1 0 32368 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_279
timestamp 1698175906
transform 1 0 32592 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_282
timestamp 1698175906
transform 1 0 32928 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_346
timestamp 1698175906
transform 1 0 40096 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_348
timestamp 1698175906
transform 1 0 40320 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_2
timestamp 1698175906
transform 1 0 1568 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698175906
transform 1 0 5152 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_37
timestamp 1698175906
transform 1 0 5488 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_101
timestamp 1698175906
transform 1 0 12656 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_107
timestamp 1698175906
transform 1 0 13328 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_123
timestamp 1698175906
transform 1 0 15120 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_136
timestamp 1698175906
transform 1 0 16576 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_144
timestamp 1698175906
transform 1 0 17472 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_148
timestamp 1698175906
transform 1 0 17920 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_151
timestamp 1698175906
transform 1 0 18256 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_167
timestamp 1698175906
transform 1 0 20048 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_177
timestamp 1698175906
transform 1 0 21168 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_241
timestamp 1698175906
transform 1 0 28336 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_247
timestamp 1698175906
transform 1 0 29008 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_311
timestamp 1698175906
transform 1 0 36176 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_317
timestamp 1698175906
transform 1 0 36848 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_2
timestamp 1698175906
transform 1 0 1568 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_66
timestamp 1698175906
transform 1 0 8736 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_72
timestamp 1698175906
transform 1 0 9408 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_136
timestamp 1698175906
transform 1 0 16576 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_142
timestamp 1698175906
transform 1 0 17248 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_146
timestamp 1698175906
transform 1 0 17696 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_212
timestamp 1698175906
transform 1 0 25088 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_276
timestamp 1698175906
transform 1 0 32256 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_282
timestamp 1698175906
transform 1 0 32928 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_346
timestamp 1698175906
transform 1 0 40096 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_348
timestamp 1698175906
transform 1 0 40320 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698175906
transform 1 0 1568 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698175906
transform 1 0 5152 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_37
timestamp 1698175906
transform 1 0 5488 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_101
timestamp 1698175906
transform 1 0 12656 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_107
timestamp 1698175906
transform 1 0 13328 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_171
timestamp 1698175906
transform 1 0 20496 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_177
timestamp 1698175906
transform 1 0 21168 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_241
timestamp 1698175906
transform 1 0 28336 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_247
timestamp 1698175906
transform 1 0 29008 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_311
timestamp 1698175906
transform 1 0 36176 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_317
timestamp 1698175906
transform 1 0 36848 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2
timestamp 1698175906
transform 1 0 1568 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_66
timestamp 1698175906
transform 1 0 8736 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_72
timestamp 1698175906
transform 1 0 9408 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_136
timestamp 1698175906
transform 1 0 16576 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_142
timestamp 1698175906
transform 1 0 17248 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_206
timestamp 1698175906
transform 1 0 24416 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_212
timestamp 1698175906
transform 1 0 25088 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_276
timestamp 1698175906
transform 1 0 32256 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_282
timestamp 1698175906
transform 1 0 32928 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_346
timestamp 1698175906
transform 1 0 40096 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_348
timestamp 1698175906
transform 1 0 40320 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_2
timestamp 1698175906
transform 1 0 1568 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698175906
transform 1 0 5152 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_37
timestamp 1698175906
transform 1 0 5488 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_101
timestamp 1698175906
transform 1 0 12656 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_107
timestamp 1698175906
transform 1 0 13328 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_171
timestamp 1698175906
transform 1 0 20496 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_177
timestamp 1698175906
transform 1 0 21168 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_241
timestamp 1698175906
transform 1 0 28336 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_247
timestamp 1698175906
transform 1 0 29008 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_311
timestamp 1698175906
transform 1 0 36176 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_317
timestamp 1698175906
transform 1 0 36848 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2
timestamp 1698175906
transform 1 0 1568 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_66
timestamp 1698175906
transform 1 0 8736 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_72
timestamp 1698175906
transform 1 0 9408 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_136
timestamp 1698175906
transform 1 0 16576 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_142
timestamp 1698175906
transform 1 0 17248 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_206
timestamp 1698175906
transform 1 0 24416 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_212
timestamp 1698175906
transform 1 0 25088 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_276
timestamp 1698175906
transform 1 0 32256 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_282
timestamp 1698175906
transform 1 0 32928 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_346
timestamp 1698175906
transform 1 0 40096 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_348
timestamp 1698175906
transform 1 0 40320 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698175906
transform 1 0 1568 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698175906
transform 1 0 5152 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_37
timestamp 1698175906
transform 1 0 5488 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_101
timestamp 1698175906
transform 1 0 12656 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_107
timestamp 1698175906
transform 1 0 13328 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_171
timestamp 1698175906
transform 1 0 20496 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_177
timestamp 1698175906
transform 1 0 21168 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_241
timestamp 1698175906
transform 1 0 28336 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_247
timestamp 1698175906
transform 1 0 29008 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_311
timestamp 1698175906
transform 1 0 36176 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_317
timestamp 1698175906
transform 1 0 36848 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_2
timestamp 1698175906
transform 1 0 1568 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_66
timestamp 1698175906
transform 1 0 8736 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_72
timestamp 1698175906
transform 1 0 9408 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_136
timestamp 1698175906
transform 1 0 16576 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_142
timestamp 1698175906
transform 1 0 17248 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_206
timestamp 1698175906
transform 1 0 24416 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_212
timestamp 1698175906
transform 1 0 25088 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_276
timestamp 1698175906
transform 1 0 32256 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_282
timestamp 1698175906
transform 1 0 32928 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_346
timestamp 1698175906
transform 1 0 40096 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_348
timestamp 1698175906
transform 1 0 40320 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698175906
transform 1 0 1568 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698175906
transform 1 0 5152 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_37
timestamp 1698175906
transform 1 0 5488 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_101
timestamp 1698175906
transform 1 0 12656 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_107
timestamp 1698175906
transform 1 0 13328 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_171
timestamp 1698175906
transform 1 0 20496 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_177
timestamp 1698175906
transform 1 0 21168 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_241
timestamp 1698175906
transform 1 0 28336 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_247
timestamp 1698175906
transform 1 0 29008 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_311
timestamp 1698175906
transform 1 0 36176 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_317
timestamp 1698175906
transform 1 0 36848 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2
timestamp 1698175906
transform 1 0 1568 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1698175906
transform 1 0 8736 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_72
timestamp 1698175906
transform 1 0 9408 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_136
timestamp 1698175906
transform 1 0 16576 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_142
timestamp 1698175906
transform 1 0 17248 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_206
timestamp 1698175906
transform 1 0 24416 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_212
timestamp 1698175906
transform 1 0 25088 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_276
timestamp 1698175906
transform 1 0 32256 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_282
timestamp 1698175906
transform 1 0 32928 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_346
timestamp 1698175906
transform 1 0 40096 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_348
timestamp 1698175906
transform 1 0 40320 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_2
timestamp 1698175906
transform 1 0 1568 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698175906
transform 1 0 5152 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_37
timestamp 1698175906
transform 1 0 5488 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_101
timestamp 1698175906
transform 1 0 12656 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_107
timestamp 1698175906
transform 1 0 13328 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_123
timestamp 1698175906
transform 1 0 15120 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_131
timestamp 1698175906
transform 1 0 16016 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_159
timestamp 1698175906
transform 1 0 19152 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_177
timestamp 1698175906
transform 1 0 21168 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_241
timestamp 1698175906
transform 1 0 28336 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_247
timestamp 1698175906
transform 1 0 29008 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_311
timestamp 1698175906
transform 1 0 36176 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_317
timestamp 1698175906
transform 1 0 36848 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_333
timestamp 1698175906
transform 1 0 38640 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_341
timestamp 1698175906
transform 1 0 39536 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_2
timestamp 1698175906
transform 1 0 1568 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_66
timestamp 1698175906
transform 1 0 8736 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_72
timestamp 1698175906
transform 1 0 9408 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_136
timestamp 1698175906
transform 1 0 16576 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_168
timestamp 1698175906
transform 1 0 20160 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_200
timestamp 1698175906
transform 1 0 23744 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_208
timestamp 1698175906
transform 1 0 24640 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_212
timestamp 1698175906
transform 1 0 25088 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_228
timestamp 1698175906
transform 1 0 26880 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_255
timestamp 1698175906
transform 1 0 29904 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_271
timestamp 1698175906
transform 1 0 31696 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_279
timestamp 1698175906
transform 1 0 32592 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_282
timestamp 1698175906
transform 1 0 32928 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_346
timestamp 1698175906
transform 1 0 40096 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_348
timestamp 1698175906
transform 1 0 40320 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_2
timestamp 1698175906
transform 1 0 1568 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_36
timestamp 1698175906
transform 1 0 5376 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_70
timestamp 1698175906
transform 1 0 9184 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_104
timestamp 1698175906
transform 1 0 12992 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_138
timestamp 1698175906
transform 1 0 16800 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_142
timestamp 1698175906
transform 1 0 17248 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_172
timestamp 1698175906
transform 1 0 20608 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_174
timestamp 1698175906
transform 1 0 20832 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_201
timestamp 1698175906
transform 1 0 23856 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_203
timestamp 1698175906
transform 1 0 24080 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_232
timestamp 1698175906
transform 1 0 27328 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_236
timestamp 1698175906
transform 1 0 27776 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_240
timestamp 1698175906
transform 1 0 28224 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_274
timestamp 1698175906
transform 1 0 32032 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_308
timestamp 1698175906
transform 1 0 35840 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_342
timestamp 1698175906
transform 1 0 39648 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_346
timestamp 1698175906
transform 1 0 40096 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_348
timestamp 1698175906
transform 1 0 40320 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita49_25 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 39984 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita49_26
timestamp 1698175906
transform 1 0 39984 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 4480 0 -1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output2
timestamp 1698175906
transform 1 0 37520 0 -1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output3
timestamp 1698175906
transform 1 0 37520 0 1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output4
timestamp 1698175906
transform 1 0 26992 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output5
timestamp 1698175906
transform -1 0 4480 0 1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output6
timestamp 1698175906
transform 1 0 17472 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output7
timestamp 1698175906
transform -1 0 4480 0 -1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output8
timestamp 1698175906
transform 1 0 16240 0 1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output9
timestamp 1698175906
transform 1 0 37520 0 1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output10
timestamp 1698175906
transform 1 0 37520 0 1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output11
timestamp 1698175906
transform 1 0 24416 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output12
timestamp 1698175906
transform 1 0 37520 0 1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output13
timestamp 1698175906
transform 1 0 20944 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output14
timestamp 1698175906
transform 1 0 20608 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output15
timestamp 1698175906
transform 1 0 17472 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output16
timestamp 1698175906
transform 1 0 37520 0 1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output17
timestamp 1698175906
transform 1 0 24416 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output18
timestamp 1698175906
transform 1 0 25088 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output19
timestamp 1698175906
transform 1 0 17248 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output20
timestamp 1698175906
transform 1 0 37520 0 -1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output21
timestamp 1698175906
transform 1 0 37520 0 -1 15680
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output22
timestamp 1698175906
transform -1 0 4480 0 -1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output23
timestamp 1698175906
transform -1 0 4480 0 1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output24
timestamp 1698175906
transform 1 0 37520 0 -1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_45 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698175906
transform -1 0 40656 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_46
timestamp 1698175906
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698175906
transform -1 0 40656 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_47
timestamp 1698175906
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698175906
transform -1 0 40656 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_48
timestamp 1698175906
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698175906
transform -1 0 40656 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_49
timestamp 1698175906
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698175906
transform -1 0 40656 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_50
timestamp 1698175906
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698175906
transform -1 0 40656 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_51
timestamp 1698175906
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698175906
transform -1 0 40656 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_52
timestamp 1698175906
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698175906
transform -1 0 40656 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_53
timestamp 1698175906
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698175906
transform -1 0 40656 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_54
timestamp 1698175906
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698175906
transform -1 0 40656 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_55
timestamp 1698175906
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698175906
transform -1 0 40656 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_56
timestamp 1698175906
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698175906
transform -1 0 40656 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_57
timestamp 1698175906
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698175906
transform -1 0 40656 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_58
timestamp 1698175906
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698175906
transform -1 0 40656 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_59
timestamp 1698175906
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698175906
transform -1 0 40656 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_60
timestamp 1698175906
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698175906
transform -1 0 40656 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_61
timestamp 1698175906
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698175906
transform -1 0 40656 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_62
timestamp 1698175906
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698175906
transform -1 0 40656 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_63
timestamp 1698175906
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698175906
transform -1 0 40656 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_64
timestamp 1698175906
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698175906
transform -1 0 40656 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_65
timestamp 1698175906
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698175906
transform -1 0 40656 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_66
timestamp 1698175906
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698175906
transform -1 0 40656 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_67
timestamp 1698175906
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698175906
transform -1 0 40656 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_68
timestamp 1698175906
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698175906
transform -1 0 40656 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_69
timestamp 1698175906
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698175906
transform -1 0 40656 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_70
timestamp 1698175906
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698175906
transform -1 0 40656 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_71
timestamp 1698175906
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698175906
transform -1 0 40656 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_72
timestamp 1698175906
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698175906
transform -1 0 40656 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_73
timestamp 1698175906
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698175906
transform -1 0 40656 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_74
timestamp 1698175906
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698175906
transform -1 0 40656 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_75
timestamp 1698175906
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698175906
transform -1 0 40656 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_76
timestamp 1698175906
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698175906
transform -1 0 40656 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_77
timestamp 1698175906
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698175906
transform -1 0 40656 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_78
timestamp 1698175906
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698175906
transform -1 0 40656 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_79
timestamp 1698175906
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698175906
transform -1 0 40656 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_80
timestamp 1698175906
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698175906
transform -1 0 40656 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_81
timestamp 1698175906
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698175906
transform -1 0 40656 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_82
timestamp 1698175906
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698175906
transform -1 0 40656 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_83
timestamp 1698175906
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698175906
transform -1 0 40656 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_84
timestamp 1698175906
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698175906
transform -1 0 40656 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_85
timestamp 1698175906
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698175906
transform -1 0 40656 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_86
timestamp 1698175906
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698175906
transform -1 0 40656 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_87
timestamp 1698175906
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698175906
transform -1 0 40656 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_88
timestamp 1698175906
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698175906
transform -1 0 40656 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_89
timestamp 1698175906
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698175906
transform -1 0 40656 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_90 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_91
timestamp 1698175906
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_92
timestamp 1698175906
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_93
timestamp 1698175906
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_94
timestamp 1698175906
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_95
timestamp 1698175906
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_96
timestamp 1698175906
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_97
timestamp 1698175906
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_98
timestamp 1698175906
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_99
timestamp 1698175906
transform 1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_100
timestamp 1698175906
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_101
timestamp 1698175906
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_102
timestamp 1698175906
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_103
timestamp 1698175906
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_104
timestamp 1698175906
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_105
timestamp 1698175906
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_106
timestamp 1698175906
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_107
timestamp 1698175906
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_108
timestamp 1698175906
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_109
timestamp 1698175906
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_110
timestamp 1698175906
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_111
timestamp 1698175906
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_112
timestamp 1698175906
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_113
timestamp 1698175906
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_114
timestamp 1698175906
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_115
timestamp 1698175906
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_116
timestamp 1698175906
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_117
timestamp 1698175906
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_118
timestamp 1698175906
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_119
timestamp 1698175906
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_120
timestamp 1698175906
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_121
timestamp 1698175906
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_122
timestamp 1698175906
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_123
timestamp 1698175906
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_124
timestamp 1698175906
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_125
timestamp 1698175906
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_126
timestamp 1698175906
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_127
timestamp 1698175906
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_128
timestamp 1698175906
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_129
timestamp 1698175906
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_130
timestamp 1698175906
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_131
timestamp 1698175906
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_132
timestamp 1698175906
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_133
timestamp 1698175906
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_134
timestamp 1698175906
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_135
timestamp 1698175906
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_136
timestamp 1698175906
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_137
timestamp 1698175906
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_138
timestamp 1698175906
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_139
timestamp 1698175906
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_140
timestamp 1698175906
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_141
timestamp 1698175906
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_142
timestamp 1698175906
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_143
timestamp 1698175906
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_144
timestamp 1698175906
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_145
timestamp 1698175906
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_146
timestamp 1698175906
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_147
timestamp 1698175906
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_148
timestamp 1698175906
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_149
timestamp 1698175906
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_150
timestamp 1698175906
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_151
timestamp 1698175906
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_152
timestamp 1698175906
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_153
timestamp 1698175906
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_154
timestamp 1698175906
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_155
timestamp 1698175906
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_156
timestamp 1698175906
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_157
timestamp 1698175906
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_158
timestamp 1698175906
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_159
timestamp 1698175906
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_160
timestamp 1698175906
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_161
timestamp 1698175906
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_162
timestamp 1698175906
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_163
timestamp 1698175906
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_164
timestamp 1698175906
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_165
timestamp 1698175906
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_166
timestamp 1698175906
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_167
timestamp 1698175906
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_168
timestamp 1698175906
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_169
timestamp 1698175906
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_170
timestamp 1698175906
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_171
timestamp 1698175906
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_172
timestamp 1698175906
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_173
timestamp 1698175906
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_174
timestamp 1698175906
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_175
timestamp 1698175906
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_176
timestamp 1698175906
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_177
timestamp 1698175906
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_178
timestamp 1698175906
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_179
timestamp 1698175906
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_180
timestamp 1698175906
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_181
timestamp 1698175906
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_182
timestamp 1698175906
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_183
timestamp 1698175906
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_184
timestamp 1698175906
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_185
timestamp 1698175906
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_186
timestamp 1698175906
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_187
timestamp 1698175906
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_188
timestamp 1698175906
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_189
timestamp 1698175906
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_190
timestamp 1698175906
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_191
timestamp 1698175906
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_192
timestamp 1698175906
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_193
timestamp 1698175906
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_194
timestamp 1698175906
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_195
timestamp 1698175906
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_196
timestamp 1698175906
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_197
timestamp 1698175906
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_198
timestamp 1698175906
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_199
timestamp 1698175906
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_200
timestamp 1698175906
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_201
timestamp 1698175906
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_202
timestamp 1698175906
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_203
timestamp 1698175906
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_204
timestamp 1698175906
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_205
timestamp 1698175906
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_206
timestamp 1698175906
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_207
timestamp 1698175906
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_208
timestamp 1698175906
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_209
timestamp 1698175906
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_210
timestamp 1698175906
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_211
timestamp 1698175906
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_212
timestamp 1698175906
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_213
timestamp 1698175906
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_214
timestamp 1698175906
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_215
timestamp 1698175906
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_216
timestamp 1698175906
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_217
timestamp 1698175906
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_218
timestamp 1698175906
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_219
timestamp 1698175906
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_220
timestamp 1698175906
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_221
timestamp 1698175906
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_222
timestamp 1698175906
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_223
timestamp 1698175906
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_224
timestamp 1698175906
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_225
timestamp 1698175906
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_226
timestamp 1698175906
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_227
timestamp 1698175906
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_228
timestamp 1698175906
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_229
timestamp 1698175906
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_230
timestamp 1698175906
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_231
timestamp 1698175906
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_232
timestamp 1698175906
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_233
timestamp 1698175906
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_234
timestamp 1698175906
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_235
timestamp 1698175906
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_236
timestamp 1698175906
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_237
timestamp 1698175906
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_238
timestamp 1698175906
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_239
timestamp 1698175906
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_240
timestamp 1698175906
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_241
timestamp 1698175906
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_242
timestamp 1698175906
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_243
timestamp 1698175906
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_244
timestamp 1698175906
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_245
timestamp 1698175906
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_246
timestamp 1698175906
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_247
timestamp 1698175906
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_248
timestamp 1698175906
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_249
timestamp 1698175906
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_250
timestamp 1698175906
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_251
timestamp 1698175906
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_252
timestamp 1698175906
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_253
timestamp 1698175906
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_254
timestamp 1698175906
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_255
timestamp 1698175906
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_256
timestamp 1698175906
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_257
timestamp 1698175906
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_258
timestamp 1698175906
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_259
timestamp 1698175906
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_260
timestamp 1698175906
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_261
timestamp 1698175906
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_262
timestamp 1698175906
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_263
timestamp 1698175906
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_264
timestamp 1698175906
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_265
timestamp 1698175906
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_266
timestamp 1698175906
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_267
timestamp 1698175906
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_268
timestamp 1698175906
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_269
timestamp 1698175906
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_270
timestamp 1698175906
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_271
timestamp 1698175906
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_272
timestamp 1698175906
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_273
timestamp 1698175906
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_274
timestamp 1698175906
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_275
timestamp 1698175906
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_276
timestamp 1698175906
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_277
timestamp 1698175906
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_278
timestamp 1698175906
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_279
timestamp 1698175906
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_280
timestamp 1698175906
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_281
timestamp 1698175906
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_282
timestamp 1698175906
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_283
timestamp 1698175906
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_284
timestamp 1698175906
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_285
timestamp 1698175906
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_286
timestamp 1698175906
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_287
timestamp 1698175906
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_288
timestamp 1698175906
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_289
timestamp 1698175906
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_290
timestamp 1698175906
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_291
timestamp 1698175906
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_292
timestamp 1698175906
transform 1 0 32704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_293
timestamp 1698175906
transform 1 0 5152 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_294
timestamp 1698175906
transform 1 0 8960 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_295
timestamp 1698175906
transform 1 0 12768 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_296
timestamp 1698175906
transform 1 0 16576 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_297
timestamp 1698175906
transform 1 0 20384 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_298
timestamp 1698175906
transform 1 0 24192 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_299
timestamp 1698175906
transform 1 0 28000 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_300
timestamp 1698175906
transform 1 0 31808 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_301
timestamp 1698175906
transform 1 0 35616 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_302
timestamp 1698175906
transform 1 0 39424 0 1 37632
box -86 -86 310 870
<< labels >>
flabel metal3 s 0 27552 800 27664 0 FreeSans 448 0 0 0 clk
port 0 nsew signal input
flabel metal3 s 41200 36288 42000 36400 0 FreeSans 448 0 0 0 segm[0]
port 1 nsew signal tristate
flabel metal3 s 0 24192 800 24304 0 FreeSans 448 0 0 0 segm[10]
port 2 nsew signal tristate
flabel metal3 s 41200 22848 42000 22960 0 FreeSans 448 0 0 0 segm[11]
port 3 nsew signal tristate
flabel metal3 s 41200 26880 42000 26992 0 FreeSans 448 0 0 0 segm[12]
port 4 nsew signal tristate
flabel metal2 s 26880 41200 26992 42000 0 FreeSans 448 90 0 0 segm[13]
port 5 nsew signal tristate
flabel metal3 s 0 18816 800 18928 0 FreeSans 448 0 0 0 segm[1]
port 6 nsew signal tristate
flabel metal2 s 17472 41200 17584 42000 0 FreeSans 448 90 0 0 segm[2]
port 7 nsew signal tristate
flabel metal3 s 41200 8736 42000 8848 0 FreeSans 448 0 0 0 segm[3]
port 8 nsew signal tristate
flabel metal3 s 0 19488 800 19600 0 FreeSans 448 0 0 0 segm[4]
port 9 nsew signal tristate
flabel metal2 s 16128 41200 16240 42000 0 FreeSans 448 90 0 0 segm[5]
port 10 nsew signal tristate
flabel metal3 s 41200 20160 42000 20272 0 FreeSans 448 0 0 0 segm[6]
port 11 nsew signal tristate
flabel metal3 s 41200 22176 42000 22288 0 FreeSans 448 0 0 0 segm[7]
port 12 nsew signal tristate
flabel metal2 s 23520 41200 23632 42000 0 FreeSans 448 90 0 0 segm[8]
port 13 nsew signal tristate
flabel metal3 s 41200 24864 42000 24976 0 FreeSans 448 0 0 0 segm[9]
port 14 nsew signal tristate
flabel metal2 s 20832 41200 20944 42000 0 FreeSans 448 90 0 0 sel[0]
port 15 nsew signal tristate
flabel metal2 s 20160 0 20272 800 0 FreeSans 448 90 0 0 sel[10]
port 16 nsew signal tristate
flabel metal2 s 18144 0 18256 800 0 FreeSans 448 90 0 0 sel[11]
port 17 nsew signal tristate
flabel metal3 s 41200 16800 42000 16912 0 FreeSans 448 0 0 0 sel[1]
port 18 nsew signal tristate
flabel metal2 s 22848 0 22960 800 0 FreeSans 448 90 0 0 sel[2]
port 19 nsew signal tristate
flabel metal2 s 24864 0 24976 800 0 FreeSans 448 90 0 0 sel[3]
port 20 nsew signal tristate
flabel metal2 s 16800 41200 16912 42000 0 FreeSans 448 90 0 0 sel[4]
port 21 nsew signal tristate
flabel metal3 s 41200 16128 42000 16240 0 FreeSans 448 0 0 0 sel[5]
port 22 nsew signal tristate
flabel metal3 s 41200 14784 42000 14896 0 FreeSans 448 0 0 0 sel[6]
port 23 nsew signal tristate
flabel metal3 s 0 20832 800 20944 0 FreeSans 448 0 0 0 sel[7]
port 24 nsew signal tristate
flabel metal3 s 0 23520 800 23632 0 FreeSans 448 0 0 0 sel[8]
port 25 nsew signal tristate
flabel metal3 s 41200 19488 42000 19600 0 FreeSans 448 0 0 0 sel[9]
port 26 nsew signal tristate
flabel metal4 s 4448 3076 4768 38476 0 FreeSans 1280 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 35168 3076 35488 38476 0 FreeSans 1280 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 19808 3076 20128 38476 0 FreeSans 1280 90 0 0 vss
port 28 nsew ground bidirectional
rlabel metal1 21000 38416 21000 38416 0 vdd
rlabel metal1 21000 37632 21000 37632 0 vss
rlabel metal2 25704 15512 25704 15512 0 _000_
rlabel metal2 26768 15400 26768 15400 0 _001_
rlabel metal3 16352 26936 16352 26936 0 _002_
rlabel metal2 23464 13272 23464 13272 0 _003_
rlabel metal2 21112 14056 21112 14056 0 _004_
rlabel metal2 24920 16408 24920 16408 0 _005_
rlabel metal2 19656 27496 19656 27496 0 _006_
rlabel metal2 12040 19600 12040 19600 0 _007_
rlabel metal2 14840 24360 14840 24360 0 _008_
rlabel metal3 16128 27720 16128 27720 0 _009_
rlabel metal2 26488 19600 26488 19600 0 _010_
rlabel metal2 18648 13272 18648 13272 0 _011_
rlabel metal2 14728 14056 14728 14056 0 _012_
rlabel metal2 29008 18984 29008 18984 0 _013_
rlabel metal2 26040 22736 26040 22736 0 _014_
rlabel metal2 23352 26712 23352 26712 0 _015_
rlabel metal2 29288 24304 29288 24304 0 _016_
rlabel metal2 28616 21672 28616 21672 0 _017_
rlabel metal2 25592 26712 25592 26712 0 _018_
rlabel metal2 25592 25704 25592 25704 0 _019_
rlabel metal3 12880 23800 12880 23800 0 _020_
rlabel metal2 12040 21224 12040 21224 0 _021_
rlabel metal3 22904 15512 22904 15512 0 _022_
rlabel metal2 15400 19152 15400 19152 0 _023_
rlabel metal2 13832 17248 13832 17248 0 _024_
rlabel metal2 12824 21896 12824 21896 0 _025_
rlabel metal3 25200 21672 25200 21672 0 _026_
rlabel metal3 25256 23352 25256 23352 0 _027_
rlabel metal2 25480 17136 25480 17136 0 _028_
rlabel metal2 22008 23968 22008 23968 0 _029_
rlabel metal2 21112 26320 21112 26320 0 _030_
rlabel metal2 21224 17360 21224 17360 0 _031_
rlabel metal2 18648 27160 18648 27160 0 _032_
rlabel metal3 16968 27048 16968 27048 0 _033_
rlabel metal2 22568 22120 22568 22120 0 _034_
rlabel metal2 22904 22960 22904 22960 0 _035_
rlabel metal2 20888 25760 20888 25760 0 _036_
rlabel metal2 22960 21112 22960 21112 0 _037_
rlabel metal3 24752 13720 24752 13720 0 _038_
rlabel metal2 24248 18480 24248 18480 0 _039_
rlabel metal2 22120 14560 22120 14560 0 _040_
rlabel metal2 21672 14784 21672 14784 0 _041_
rlabel metal2 24248 17192 24248 17192 0 _042_
rlabel metal2 24864 16856 24864 16856 0 _043_
rlabel metal2 20328 25760 20328 25760 0 _044_
rlabel metal2 22344 23688 22344 23688 0 _045_
rlabel metal2 20440 26656 20440 26656 0 _046_
rlabel metal2 15512 19488 15512 19488 0 _047_
rlabel metal2 15624 19432 15624 19432 0 _048_
rlabel metal2 12936 19880 12936 19880 0 _049_
rlabel metal3 20916 23240 20916 23240 0 _050_
rlabel metal3 16408 23912 16408 23912 0 _051_
rlabel metal2 15568 24024 15568 24024 0 _052_
rlabel metal2 17528 26600 17528 26600 0 _053_
rlabel metal2 18312 27552 18312 27552 0 _054_
rlabel metal2 22456 23632 22456 23632 0 _055_
rlabel metal2 26264 19936 26264 19936 0 _056_
rlabel metal2 25480 23072 25480 23072 0 _057_
rlabel metal2 28728 22848 28728 22848 0 _058_
rlabel metal3 20160 13944 20160 13944 0 _059_
rlabel metal2 18312 14168 18312 14168 0 _060_
rlabel metal3 23408 18536 23408 18536 0 _061_
rlabel metal2 25312 20216 25312 20216 0 _062_
rlabel metal2 24136 18536 24136 18536 0 _063_
rlabel metal2 25816 21504 25816 21504 0 _064_
rlabel metal2 29176 21448 29176 21448 0 _065_
rlabel metal2 29064 19880 29064 19880 0 _066_
rlabel metal3 24640 26264 24640 26264 0 _067_
rlabel metal3 24864 21560 24864 21560 0 _068_
rlabel metal2 25592 22344 25592 22344 0 _069_
rlabel metal2 22904 24752 22904 24752 0 _070_
rlabel metal2 23240 25872 23240 25872 0 _071_
rlabel metal3 26208 23912 26208 23912 0 _072_
rlabel metal2 29064 24584 29064 24584 0 _073_
rlabel metal2 29960 22848 29960 22848 0 _074_
rlabel metal3 25592 23128 25592 23128 0 _075_
rlabel metal3 26600 26264 26600 26264 0 _076_
rlabel metal2 23184 24920 23184 24920 0 _077_
rlabel metal2 22232 22792 22232 22792 0 _078_
rlabel metal2 22568 23520 22568 23520 0 _079_
rlabel metal2 25424 25480 25424 25480 0 _080_
rlabel metal2 25816 25592 25816 25592 0 _081_
rlabel metal2 17528 21840 17528 21840 0 _082_
rlabel metal2 24024 23296 24024 23296 0 _083_
rlabel via2 21784 24696 21784 24696 0 _084_
rlabel metal2 20552 21952 20552 21952 0 _085_
rlabel via2 20552 19320 20552 19320 0 _086_
rlabel metal2 14168 22680 14168 22680 0 _087_
rlabel metal2 13048 23464 13048 23464 0 _088_
rlabel metal2 19152 23912 19152 23912 0 _089_
rlabel metal2 15848 23184 15848 23184 0 _090_
rlabel metal2 13944 23296 13944 23296 0 _091_
rlabel metal2 21336 21224 21336 21224 0 _092_
rlabel metal2 20720 20552 20720 20552 0 _093_
rlabel metal3 20608 20328 20608 20328 0 _094_
rlabel metal2 19320 22232 19320 22232 0 _095_
rlabel metal2 21560 22232 21560 22232 0 _096_
rlabel metal2 21896 23856 21896 23856 0 _097_
rlabel metal3 17528 22064 17528 22064 0 _098_
rlabel metal2 25480 19544 25480 19544 0 _099_
rlabel metal2 13496 21224 13496 21224 0 _100_
rlabel metal2 19264 23240 19264 23240 0 _101_
rlabel metal2 20216 25144 20216 25144 0 _102_
rlabel metal2 24584 19040 24584 19040 0 _103_
rlabel metal3 20776 24584 20776 24584 0 _104_
rlabel metal3 21000 22120 21000 22120 0 _105_
rlabel metal3 21336 17528 21336 17528 0 _106_
rlabel metal2 23464 17976 23464 17976 0 _107_
rlabel metal2 17752 18368 17752 18368 0 _108_
rlabel metal2 22232 22232 22232 22232 0 _109_
rlabel metal2 23016 22512 23016 22512 0 _110_
rlabel metal3 22120 17640 22120 17640 0 _111_
rlabel metal3 23184 17752 23184 17752 0 _112_
rlabel metal2 19320 18032 19320 18032 0 _113_
rlabel metal2 13832 22232 13832 22232 0 _114_
rlabel metal2 27384 14896 27384 14896 0 _115_
rlabel metal2 26712 14224 26712 14224 0 _116_
rlabel metal3 23240 17080 23240 17080 0 _117_
rlabel metal3 23968 15288 23968 15288 0 _118_
rlabel metal2 22568 21112 22568 21112 0 _119_
rlabel metal3 26040 15288 26040 15288 0 _120_
rlabel metal3 26992 16296 26992 16296 0 _121_
rlabel metal3 5838 27608 5838 27608 0 clk
rlabel metal2 23576 20468 23576 20468 0 clknet_0_clk
rlabel metal2 18088 29008 18088 29008 0 clknet_1_0__leaf_clk
rlabel metal3 23128 27048 23128 27048 0 clknet_1_1__leaf_clk
rlabel metal3 18648 17416 18648 17416 0 dut49.count\[0\]
rlabel metal2 21448 18816 21448 18816 0 dut49.count\[1\]
rlabel metal3 16856 21448 16856 21448 0 dut49.count\[2\]
rlabel metal2 20440 22736 20440 22736 0 dut49.count\[3\]
rlabel metal3 13048 24640 13048 24640 0 net1
rlabel metal2 28168 22512 28168 22512 0 net10
rlabel metal2 23800 26320 23800 26320 0 net11
rlabel metal2 30632 25032 30632 25032 0 net12
rlabel metal2 20552 27104 20552 27104 0 net13
rlabel metal2 20776 8288 20776 8288 0 net14
rlabel metal2 18144 13608 18144 13608 0 net15
rlabel metal2 27048 16912 27048 16912 0 net16
rlabel metal2 23240 8568 23240 8568 0 net17
rlabel metal2 25592 8680 25592 8680 0 net18
rlabel metal2 17360 37240 17360 37240 0 net19
rlabel metal2 30856 22288 30856 22288 0 net2
rlabel metal2 27496 15512 27496 15512 0 net20
rlabel metal2 26936 14280 26936 14280 0 net21
rlabel metal2 9912 20776 9912 20776 0 net22
rlabel metal3 6356 23912 6356 23912 0 net23
rlabel metal2 25704 19656 25704 19656 0 net24
rlabel metal3 40754 36344 40754 36344 0 net25
rlabel metal2 40264 8960 40264 8960 0 net26
rlabel metal2 27160 26768 27160 26768 0 net3
rlabel metal3 27328 26488 27328 26488 0 net4
rlabel metal2 12376 18928 12376 18928 0 net5
rlabel metal2 18536 27272 18536 27272 0 net6
rlabel metal2 9912 19656 9912 19656 0 net7
rlabel metal3 16632 28504 16632 28504 0 net8
rlabel metal3 30072 20552 30072 20552 0 net9
rlabel metal3 1358 24248 1358 24248 0 segm[10]
rlabel metal3 40642 22904 40642 22904 0 segm[11]
rlabel metal2 40040 27048 40040 27048 0 segm[12]
rlabel metal2 26936 39354 26936 39354 0 segm[13]
rlabel metal3 1358 18872 1358 18872 0 segm[1]
rlabel metal2 17528 39746 17528 39746 0 segm[2]
rlabel metal3 1358 19544 1358 19544 0 segm[4]
rlabel metal2 16184 38962 16184 38962 0 segm[5]
rlabel metal2 40040 20552 40040 20552 0 segm[6]
rlabel metal2 40040 22344 40040 22344 0 segm[7]
rlabel metal2 23576 39746 23576 39746 0 segm[8]
rlabel metal2 40040 25256 40040 25256 0 segm[9]
rlabel metal2 20888 39746 20888 39746 0 sel[0]
rlabel metal3 21000 3416 21000 3416 0 sel[10]
rlabel metal2 18200 2058 18200 2058 0 sel[11]
rlabel metal2 40040 17304 40040 17304 0 sel[1]
rlabel metal3 24248 3640 24248 3640 0 sel[2]
rlabel metal3 25592 4088 25592 4088 0 sel[3]
rlabel metal2 16856 39354 16856 39354 0 sel[4]
rlabel metal2 40040 16408 40040 16408 0 sel[5]
rlabel metal2 40040 15008 40040 15008 0 sel[6]
rlabel metal3 1358 20888 1358 20888 0 sel[7]
rlabel metal3 1358 23576 1358 23576 0 sel[8]
rlabel metal2 40040 19656 40040 19656 0 sel[9]
<< properties >>
string FIXED_BBOX 0 0 42000 42000
<< end >>
