magic
tech gf180mcuD
magscale 1 10
timestamp 1699642162
<< metal1 >>
rect 18722 38558 18734 38610
rect 18786 38607 18798 38610
rect 19730 38607 19742 38610
rect 18786 38561 19742 38607
rect 18786 38558 18798 38561
rect 19730 38558 19742 38561
rect 19794 38558 19806 38610
rect 1344 38442 40656 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 40656 38442
rect 1344 38356 40656 38390
rect 21758 38274 21810 38286
rect 21758 38210 21810 38222
rect 25566 38274 25618 38286
rect 25566 38210 25618 38222
rect 18162 38110 18174 38162
rect 18226 38110 18238 38162
rect 19730 37998 19742 38050
rect 19794 37998 19806 38050
rect 20738 37998 20750 38050
rect 20802 37998 20814 38050
rect 24546 37998 24558 38050
rect 24610 37998 24622 38050
rect 1344 37658 40656 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 40656 37658
rect 1344 37572 40656 37606
rect 20078 37490 20130 37502
rect 20078 37426 20130 37438
rect 26238 37490 26290 37502
rect 26238 37426 26290 37438
rect 19506 37214 19518 37266
rect 19570 37214 19582 37266
rect 25218 37214 25230 37266
rect 25282 37214 25294 37266
rect 1344 36874 40656 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 40656 36874
rect 1344 36788 40656 36822
rect 19742 36370 19794 36382
rect 19742 36306 19794 36318
rect 1344 36090 40656 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 40656 36090
rect 1344 36004 40656 36038
rect 1344 35306 40656 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 40656 35306
rect 1344 35220 40656 35254
rect 1344 34522 40656 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 40656 34522
rect 1344 34436 40656 34470
rect 1344 33738 40656 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 40656 33738
rect 1344 33652 40656 33686
rect 1344 32954 40656 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 40656 32954
rect 1344 32868 40656 32902
rect 1344 32170 40656 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 40656 32170
rect 1344 32084 40656 32118
rect 1344 31386 40656 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 40656 31386
rect 1344 31300 40656 31334
rect 1344 30602 40656 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 40656 30602
rect 1344 30516 40656 30550
rect 1344 29818 40656 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 40656 29818
rect 1344 29732 40656 29766
rect 1344 29034 40656 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 40656 29034
rect 1344 28948 40656 28982
rect 1344 28250 40656 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 40656 28250
rect 1344 28164 40656 28198
rect 4274 27806 4286 27858
rect 4338 27806 4350 27858
rect 1934 27634 1986 27646
rect 1934 27570 1986 27582
rect 1344 27466 40656 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 40656 27466
rect 1344 27380 40656 27414
rect 2034 27134 2046 27186
rect 2098 27134 2110 27186
rect 17266 27134 17278 27186
rect 17330 27134 17342 27186
rect 4274 27022 4286 27074
rect 4338 27022 4350 27074
rect 14354 27022 14366 27074
rect 14418 27022 14430 27074
rect 20178 27022 20190 27074
rect 20242 27022 20254 27074
rect 20638 26962 20690 26974
rect 14130 26910 14142 26962
rect 14194 26910 14206 26962
rect 19394 26910 19406 26962
rect 19458 26910 19470 26962
rect 20638 26898 20690 26910
rect 1344 26682 40656 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 40656 26682
rect 1344 26596 40656 26630
rect 19518 26514 19570 26526
rect 15026 26462 15038 26514
rect 15090 26462 15102 26514
rect 19842 26462 19854 26514
rect 19906 26462 19918 26514
rect 19518 26450 19570 26462
rect 18846 26402 18898 26414
rect 18846 26338 18898 26350
rect 4274 26238 4286 26290
rect 4338 26238 4350 26290
rect 14578 26238 14590 26290
rect 14642 26238 14654 26290
rect 15250 26238 15262 26290
rect 15314 26238 15326 26290
rect 37874 26238 37886 26290
rect 37938 26238 37950 26290
rect 15934 26178 15986 26190
rect 11778 26126 11790 26178
rect 11842 26126 11854 26178
rect 13906 26126 13918 26178
rect 13970 26126 13982 26178
rect 15934 26114 15986 26126
rect 18958 26178 19010 26190
rect 18958 26114 19010 26126
rect 25342 26178 25394 26190
rect 39890 26126 39902 26178
rect 39954 26126 39966 26178
rect 25342 26114 25394 26126
rect 1934 26066 1986 26078
rect 1934 26002 1986 26014
rect 1344 25898 40656 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 40656 25898
rect 1344 25812 40656 25846
rect 13582 25730 13634 25742
rect 13582 25666 13634 25678
rect 13470 25618 13522 25630
rect 2034 25566 2046 25618
rect 2098 25566 2110 25618
rect 13470 25554 13522 25566
rect 14702 25618 14754 25630
rect 19182 25618 19234 25630
rect 40014 25618 40066 25630
rect 18722 25566 18734 25618
rect 18786 25566 18798 25618
rect 24770 25566 24782 25618
rect 24834 25566 24846 25618
rect 28018 25566 28030 25618
rect 28082 25566 28094 25618
rect 14702 25554 14754 25566
rect 19182 25554 19234 25566
rect 40014 25554 40066 25566
rect 19294 25506 19346 25518
rect 4274 25454 4286 25506
rect 4338 25454 4350 25506
rect 14354 25454 14366 25506
rect 14418 25454 14430 25506
rect 15026 25454 15038 25506
rect 15090 25454 15102 25506
rect 15810 25454 15822 25506
rect 15874 25454 15886 25506
rect 19294 25442 19346 25454
rect 19518 25506 19570 25518
rect 19518 25442 19570 25454
rect 19630 25506 19682 25518
rect 21858 25454 21870 25506
rect 21922 25454 21934 25506
rect 25218 25454 25230 25506
rect 25282 25454 25294 25506
rect 37650 25454 37662 25506
rect 37714 25454 37726 25506
rect 19630 25442 19682 25454
rect 19070 25394 19122 25406
rect 16594 25342 16606 25394
rect 16658 25342 16670 25394
rect 19070 25330 19122 25342
rect 19966 25394 20018 25406
rect 22642 25342 22654 25394
rect 22706 25342 22718 25394
rect 25890 25342 25902 25394
rect 25954 25342 25966 25394
rect 19966 25330 20018 25342
rect 14590 25282 14642 25294
rect 14590 25218 14642 25230
rect 14814 25282 14866 25294
rect 14814 25218 14866 25230
rect 28478 25282 28530 25294
rect 28478 25218 28530 25230
rect 1344 25114 40656 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 40656 25114
rect 1344 25028 40656 25062
rect 17278 24946 17330 24958
rect 17278 24882 17330 24894
rect 18510 24946 18562 24958
rect 18510 24882 18562 24894
rect 23774 24946 23826 24958
rect 23774 24882 23826 24894
rect 25790 24946 25842 24958
rect 25790 24882 25842 24894
rect 26350 24946 26402 24958
rect 26350 24882 26402 24894
rect 17502 24834 17554 24846
rect 17502 24770 17554 24782
rect 18734 24834 18786 24846
rect 18734 24770 18786 24782
rect 25566 24834 25618 24846
rect 28030 24834 28082 24846
rect 27570 24782 27582 24834
rect 27634 24782 27646 24834
rect 25566 24770 25618 24782
rect 28030 24770 28082 24782
rect 14478 24722 14530 24734
rect 13906 24670 13918 24722
rect 13970 24670 13982 24722
rect 14242 24670 14254 24722
rect 14306 24670 14318 24722
rect 14478 24658 14530 24670
rect 14702 24722 14754 24734
rect 17614 24722 17666 24734
rect 14914 24670 14926 24722
rect 14978 24670 14990 24722
rect 14702 24658 14754 24670
rect 17614 24658 17666 24670
rect 18398 24722 18450 24734
rect 25454 24722 25506 24734
rect 20514 24670 20526 24722
rect 20578 24670 20590 24722
rect 18398 24658 18450 24670
rect 25454 24658 25506 24670
rect 26126 24722 26178 24734
rect 26126 24658 26178 24670
rect 26462 24722 26514 24734
rect 27918 24722 27970 24734
rect 27346 24670 27358 24722
rect 27410 24670 27422 24722
rect 37650 24670 37662 24722
rect 37714 24670 37726 24722
rect 26462 24658 26514 24670
rect 27918 24658 27970 24670
rect 14590 24610 14642 24622
rect 10994 24558 11006 24610
rect 11058 24558 11070 24610
rect 13122 24558 13134 24610
rect 13186 24558 13198 24610
rect 14590 24546 14642 24558
rect 19070 24610 19122 24622
rect 21186 24558 21198 24610
rect 21250 24558 21262 24610
rect 23314 24558 23326 24610
rect 23378 24558 23390 24610
rect 19070 24546 19122 24558
rect 28030 24498 28082 24510
rect 28030 24434 28082 24446
rect 40014 24498 40066 24510
rect 40014 24434 40066 24446
rect 1344 24330 40656 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 40656 24330
rect 1344 24244 40656 24278
rect 12910 24162 12962 24174
rect 12910 24098 12962 24110
rect 12798 24050 12850 24062
rect 12798 23986 12850 23998
rect 20414 24050 20466 24062
rect 20414 23986 20466 23998
rect 21646 24050 21698 24062
rect 29262 24050 29314 24062
rect 22642 23998 22654 24050
rect 22706 23998 22718 24050
rect 28578 23998 28590 24050
rect 28642 23998 28654 24050
rect 21646 23986 21698 23998
rect 29262 23986 29314 23998
rect 20638 23938 20690 23950
rect 18610 23886 18622 23938
rect 18674 23886 18686 23938
rect 20178 23886 20190 23938
rect 20242 23886 20254 23938
rect 20638 23874 20690 23886
rect 20750 23938 20802 23950
rect 20750 23874 20802 23886
rect 21422 23938 21474 23950
rect 23886 23938 23938 23950
rect 22530 23886 22542 23938
rect 22594 23886 22606 23938
rect 25666 23886 25678 23938
rect 25730 23886 25742 23938
rect 21422 23874 21474 23886
rect 23886 23874 23938 23886
rect 21982 23826 22034 23838
rect 21982 23762 22034 23774
rect 22206 23826 22258 23838
rect 22206 23762 22258 23774
rect 22878 23826 22930 23838
rect 22878 23762 22930 23774
rect 23438 23826 23490 23838
rect 23438 23762 23490 23774
rect 23774 23826 23826 23838
rect 26450 23774 26462 23826
rect 26514 23774 26526 23826
rect 23774 23762 23826 23774
rect 14142 23714 14194 23726
rect 15934 23714 15986 23726
rect 21310 23714 21362 23726
rect 15586 23662 15598 23714
rect 15650 23662 15662 23714
rect 18834 23662 18846 23714
rect 18898 23662 18910 23714
rect 14142 23650 14194 23662
rect 15934 23650 15986 23662
rect 21310 23650 21362 23662
rect 23662 23714 23714 23726
rect 23662 23650 23714 23662
rect 23998 23714 24050 23726
rect 23998 23650 24050 23662
rect 1344 23546 40656 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 40656 23546
rect 1344 23460 40656 23494
rect 17502 23378 17554 23390
rect 17502 23314 17554 23326
rect 17950 23378 18002 23390
rect 17950 23314 18002 23326
rect 18062 23378 18114 23390
rect 18062 23314 18114 23326
rect 22318 23378 22370 23390
rect 22318 23314 22370 23326
rect 22430 23378 22482 23390
rect 22430 23314 22482 23326
rect 22542 23378 22594 23390
rect 22542 23314 22594 23326
rect 26462 23378 26514 23390
rect 26462 23314 26514 23326
rect 26126 23266 26178 23278
rect 19282 23214 19294 23266
rect 19346 23214 19358 23266
rect 26126 23202 26178 23214
rect 26238 23266 26290 23278
rect 26238 23202 26290 23214
rect 18174 23154 18226 23166
rect 4274 23102 4286 23154
rect 4338 23102 4350 23154
rect 16818 23102 16830 23154
rect 16882 23102 16894 23154
rect 18174 23090 18226 23102
rect 18622 23154 18674 23166
rect 22206 23154 22258 23166
rect 19058 23102 19070 23154
rect 19122 23102 19134 23154
rect 22754 23102 22766 23154
rect 22818 23102 22830 23154
rect 18622 23090 18674 23102
rect 22206 23090 22258 23102
rect 18398 23042 18450 23054
rect 13906 22990 13918 23042
rect 13970 22990 13982 23042
rect 16034 22990 16046 23042
rect 16098 22990 16110 23042
rect 18398 22978 18450 22990
rect 1934 22930 1986 22942
rect 1934 22866 1986 22878
rect 1344 22762 40656 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 40656 22762
rect 1344 22676 40656 22710
rect 13582 22594 13634 22606
rect 13582 22530 13634 22542
rect 18734 22594 18786 22606
rect 18734 22530 18786 22542
rect 26574 22594 26626 22606
rect 26574 22530 26626 22542
rect 1934 22482 1986 22494
rect 16158 22482 16210 22494
rect 25230 22482 25282 22494
rect 9986 22430 9998 22482
rect 10050 22430 10062 22482
rect 24770 22430 24782 22482
rect 24834 22430 24846 22482
rect 1934 22418 1986 22430
rect 16158 22418 16210 22430
rect 25230 22418 25282 22430
rect 40014 22482 40066 22494
rect 40014 22418 40066 22430
rect 13694 22370 13746 22382
rect 17166 22370 17218 22382
rect 4274 22318 4286 22370
rect 4338 22318 4350 22370
rect 12898 22318 12910 22370
rect 12962 22318 12974 22370
rect 16930 22318 16942 22370
rect 16994 22318 17006 22370
rect 13694 22306 13746 22318
rect 17166 22306 17218 22318
rect 17390 22370 17442 22382
rect 26462 22370 26514 22382
rect 17602 22318 17614 22370
rect 17666 22318 17678 22370
rect 18722 22318 18734 22370
rect 18786 22318 18798 22370
rect 17390 22306 17442 22318
rect 21858 22306 21870 22358
rect 21922 22306 21934 22358
rect 37650 22318 37662 22370
rect 37714 22318 37726 22370
rect 26462 22306 26514 22318
rect 13582 22258 13634 22270
rect 12114 22206 12126 22258
rect 12178 22206 12190 22258
rect 13582 22194 13634 22206
rect 16046 22258 16098 22270
rect 16046 22194 16098 22206
rect 16382 22258 16434 22270
rect 16382 22194 16434 22206
rect 16606 22258 16658 22270
rect 16606 22194 16658 22206
rect 17278 22258 17330 22270
rect 19070 22258 19122 22270
rect 27358 22258 27410 22270
rect 18050 22206 18062 22258
rect 18114 22206 18126 22258
rect 22642 22206 22654 22258
rect 22706 22206 22718 22258
rect 17278 22194 17330 22206
rect 19070 22194 19122 22206
rect 27358 22194 27410 22206
rect 14142 22146 14194 22158
rect 14142 22082 14194 22094
rect 18398 22146 18450 22158
rect 18398 22082 18450 22094
rect 26574 22146 26626 22158
rect 26574 22082 26626 22094
rect 27470 22146 27522 22158
rect 27470 22082 27522 22094
rect 27694 22146 27746 22158
rect 27694 22082 27746 22094
rect 1344 21978 40656 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 40656 21978
rect 1344 21892 40656 21926
rect 13134 21810 13186 21822
rect 21982 21810 22034 21822
rect 18386 21758 18398 21810
rect 18450 21758 18462 21810
rect 13134 21746 13186 21758
rect 21982 21746 22034 21758
rect 23886 21810 23938 21822
rect 23886 21746 23938 21758
rect 24334 21810 24386 21822
rect 24334 21746 24386 21758
rect 24558 21810 24610 21822
rect 24558 21746 24610 21758
rect 26350 21810 26402 21822
rect 26350 21746 26402 21758
rect 14030 21698 14082 21710
rect 14030 21634 14082 21646
rect 20750 21698 20802 21710
rect 20750 21634 20802 21646
rect 23438 21698 23490 21710
rect 23438 21634 23490 21646
rect 13918 21586 13970 21598
rect 20638 21586 20690 21598
rect 18162 21534 18174 21586
rect 18226 21534 18238 21586
rect 13918 21522 13970 21534
rect 20638 21522 20690 21534
rect 20974 21586 21026 21598
rect 20974 21522 21026 21534
rect 21870 21586 21922 21598
rect 21870 21522 21922 21534
rect 22094 21586 22146 21598
rect 22094 21522 22146 21534
rect 22542 21586 22594 21598
rect 24222 21586 24274 21598
rect 23650 21534 23662 21586
rect 23714 21534 23726 21586
rect 25890 21534 25902 21586
rect 25954 21534 25966 21586
rect 29474 21534 29486 21586
rect 29538 21534 29550 21586
rect 37874 21534 37886 21586
rect 37938 21534 37950 21586
rect 22542 21522 22594 21534
rect 24222 21522 24274 21534
rect 23550 21474 23602 21486
rect 40014 21474 40066 21486
rect 26674 21422 26686 21474
rect 26738 21422 26750 21474
rect 28802 21422 28814 21474
rect 28866 21422 28878 21474
rect 23550 21410 23602 21422
rect 40014 21410 40066 21422
rect 13246 21362 13298 21374
rect 13246 21298 13298 21310
rect 13470 21362 13522 21374
rect 13470 21298 13522 21310
rect 25566 21362 25618 21374
rect 25566 21298 25618 21310
rect 25902 21362 25954 21374
rect 25902 21298 25954 21310
rect 1344 21194 40656 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 40656 21194
rect 1344 21108 40656 21142
rect 28590 21026 28642 21038
rect 28590 20962 28642 20974
rect 40014 20914 40066 20926
rect 16818 20862 16830 20914
rect 16882 20862 16894 20914
rect 25218 20862 25230 20914
rect 25282 20862 25294 20914
rect 40014 20850 40066 20862
rect 29934 20802 29986 20814
rect 13682 20750 13694 20802
rect 13746 20750 13758 20802
rect 20738 20750 20750 20802
rect 20802 20750 20814 20802
rect 22642 20750 22654 20802
rect 22706 20750 22718 20802
rect 28578 20750 28590 20802
rect 28642 20750 28654 20802
rect 29362 20750 29374 20802
rect 29426 20750 29438 20802
rect 37650 20750 37662 20802
rect 37714 20750 37726 20802
rect 29934 20738 29986 20750
rect 14366 20690 14418 20702
rect 28254 20690 28306 20702
rect 21298 20638 21310 20690
rect 21362 20638 21374 20690
rect 14366 20626 14418 20638
rect 28254 20626 28306 20638
rect 13470 20578 13522 20590
rect 13470 20514 13522 20526
rect 14702 20578 14754 20590
rect 14702 20514 14754 20526
rect 21646 20578 21698 20590
rect 29586 20526 29598 20578
rect 29650 20526 29662 20578
rect 30258 20526 30270 20578
rect 30322 20526 30334 20578
rect 21646 20514 21698 20526
rect 1344 20410 40656 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 40656 20410
rect 1344 20324 40656 20358
rect 14366 20242 14418 20254
rect 14366 20178 14418 20190
rect 17726 20130 17778 20142
rect 11442 20078 11454 20130
rect 11506 20078 11518 20130
rect 14690 20078 14702 20130
rect 14754 20078 14766 20130
rect 16370 20078 16382 20130
rect 16434 20078 16446 20130
rect 17726 20066 17778 20078
rect 18958 20130 19010 20142
rect 21858 20078 21870 20130
rect 21922 20078 21934 20130
rect 18958 20066 19010 20078
rect 15150 20018 15202 20030
rect 16046 20018 16098 20030
rect 10770 19966 10782 20018
rect 10834 19966 10846 20018
rect 15362 19966 15374 20018
rect 15426 19966 15438 20018
rect 19282 19966 19294 20018
rect 19346 19966 19358 20018
rect 25666 19966 25678 20018
rect 25730 19966 25742 20018
rect 37874 19966 37886 20018
rect 37938 19966 37950 20018
rect 15150 19954 15202 19966
rect 16046 19954 16098 19966
rect 14030 19906 14082 19918
rect 13570 19854 13582 19906
rect 13634 19854 13646 19906
rect 14030 19842 14082 19854
rect 15038 19906 15090 19918
rect 29038 19906 29090 19918
rect 17602 19854 17614 19906
rect 17666 19854 17678 19906
rect 26450 19854 26462 19906
rect 26514 19854 26526 19906
rect 28578 19854 28590 19906
rect 28642 19854 28654 19906
rect 15038 19842 15090 19854
rect 29038 19842 29090 19854
rect 40014 19906 40066 19918
rect 40014 19842 40066 19854
rect 17950 19794 18002 19806
rect 17950 19730 18002 19742
rect 1344 19626 40656 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 40656 19626
rect 1344 19540 40656 19574
rect 14702 19458 14754 19470
rect 14702 19394 14754 19406
rect 15262 19458 15314 19470
rect 15262 19394 15314 19406
rect 19294 19458 19346 19470
rect 22654 19458 22706 19470
rect 19618 19406 19630 19458
rect 19682 19406 19694 19458
rect 19294 19394 19346 19406
rect 22654 19394 22706 19406
rect 22990 19458 23042 19470
rect 22990 19394 23042 19406
rect 40014 19458 40066 19470
rect 40014 19394 40066 19406
rect 21534 19346 21586 19358
rect 12898 19294 12910 19346
rect 12962 19294 12974 19346
rect 16146 19294 16158 19346
rect 16210 19294 16222 19346
rect 21534 19282 21586 19294
rect 21870 19346 21922 19358
rect 21870 19282 21922 19294
rect 22430 19346 22482 19358
rect 22430 19282 22482 19294
rect 24110 19346 24162 19358
rect 24110 19282 24162 19294
rect 25790 19346 25842 19358
rect 26226 19294 26238 19346
rect 26290 19343 26302 19346
rect 26450 19343 26462 19346
rect 26290 19297 26462 19343
rect 26290 19294 26302 19297
rect 26450 19294 26462 19297
rect 26514 19294 26526 19346
rect 25790 19282 25842 19294
rect 15038 19234 15090 19246
rect 17390 19234 17442 19246
rect 20190 19234 20242 19246
rect 10098 19182 10110 19234
rect 10162 19182 10174 19234
rect 13794 19182 13806 19234
rect 13858 19182 13870 19234
rect 16482 19182 16494 19234
rect 16546 19182 16558 19234
rect 17042 19182 17054 19234
rect 17106 19182 17118 19234
rect 19282 19182 19294 19234
rect 19346 19182 19358 19234
rect 15038 19170 15090 19182
rect 17390 19170 17442 19182
rect 20190 19170 20242 19182
rect 21310 19234 21362 19246
rect 21310 19170 21362 19182
rect 21982 19234 22034 19246
rect 21982 19170 22034 19182
rect 24670 19234 24722 19246
rect 24670 19170 24722 19182
rect 24894 19234 24946 19246
rect 24894 19170 24946 19182
rect 26350 19234 26402 19246
rect 26350 19170 26402 19182
rect 26798 19234 26850 19246
rect 26798 19170 26850 19182
rect 27022 19234 27074 19246
rect 27022 19170 27074 19182
rect 27358 19234 27410 19246
rect 37650 19182 37662 19234
rect 37714 19182 37726 19234
rect 27358 19170 27410 19182
rect 14478 19122 14530 19134
rect 18958 19122 19010 19134
rect 10770 19070 10782 19122
rect 10834 19070 10846 19122
rect 14018 19070 14030 19122
rect 14082 19070 14094 19122
rect 16034 19070 16046 19122
rect 16098 19070 16110 19122
rect 14478 19058 14530 19070
rect 18958 19058 19010 19070
rect 20078 19122 20130 19134
rect 20078 19058 20130 19070
rect 20302 19122 20354 19134
rect 20302 19058 20354 19070
rect 23326 19122 23378 19134
rect 23326 19058 23378 19070
rect 24334 19122 24386 19134
rect 24334 19058 24386 19070
rect 25902 19122 25954 19134
rect 25902 19058 25954 19070
rect 14590 19010 14642 19022
rect 21758 19010 21810 19022
rect 15586 18958 15598 19010
rect 15650 18958 15662 19010
rect 17714 18958 17726 19010
rect 17778 18958 17790 19010
rect 14590 18946 14642 18958
rect 21758 18946 21810 18958
rect 23438 19010 23490 19022
rect 25678 19010 25730 19022
rect 23762 18958 23774 19010
rect 23826 18958 23838 19010
rect 25218 18958 25230 19010
rect 25282 18958 25294 19010
rect 23438 18946 23490 18958
rect 25678 18946 25730 18958
rect 27246 19010 27298 19022
rect 27246 18946 27298 18958
rect 1344 18842 40656 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 40656 18842
rect 1344 18756 40656 18790
rect 15486 18674 15538 18686
rect 15486 18610 15538 18622
rect 20638 18674 20690 18686
rect 20638 18610 20690 18622
rect 15038 18562 15090 18574
rect 15038 18498 15090 18510
rect 16270 18562 16322 18574
rect 16270 18498 16322 18510
rect 19742 18562 19794 18574
rect 23998 18562 24050 18574
rect 22754 18510 22766 18562
rect 22818 18510 22830 18562
rect 19742 18498 19794 18510
rect 23998 18498 24050 18510
rect 24110 18562 24162 18574
rect 24110 18498 24162 18510
rect 16382 18450 16434 18462
rect 17614 18450 17666 18462
rect 15698 18398 15710 18450
rect 15762 18398 15774 18450
rect 16034 18398 16046 18450
rect 16098 18398 16110 18450
rect 17378 18398 17390 18450
rect 17442 18398 17454 18450
rect 16382 18386 16434 18398
rect 17614 18386 17666 18398
rect 18622 18450 18674 18462
rect 18622 18386 18674 18398
rect 18846 18450 18898 18462
rect 21534 18450 21586 18462
rect 19954 18398 19966 18450
rect 20018 18398 20030 18450
rect 20402 18398 20414 18450
rect 20466 18398 20478 18450
rect 18846 18386 18898 18398
rect 21534 18386 21586 18398
rect 21758 18450 21810 18462
rect 21758 18386 21810 18398
rect 22430 18450 22482 18462
rect 22430 18386 22482 18398
rect 25230 18450 25282 18462
rect 25230 18386 25282 18398
rect 13134 18338 13186 18350
rect 13134 18274 13186 18286
rect 14926 18338 14978 18350
rect 14926 18274 14978 18286
rect 21310 18338 21362 18350
rect 21310 18274 21362 18286
rect 15374 18226 15426 18238
rect 17838 18226 17890 18238
rect 16818 18174 16830 18226
rect 16882 18174 16894 18226
rect 15374 18162 15426 18174
rect 17838 18162 17890 18174
rect 17950 18226 18002 18238
rect 20750 18226 20802 18238
rect 19170 18174 19182 18226
rect 19234 18174 19246 18226
rect 17950 18162 18002 18174
rect 20750 18162 20802 18174
rect 22206 18226 22258 18238
rect 22206 18162 22258 18174
rect 24110 18226 24162 18238
rect 24110 18162 24162 18174
rect 25454 18226 25506 18238
rect 25778 18174 25790 18226
rect 25842 18174 25854 18226
rect 25454 18162 25506 18174
rect 1344 18058 40656 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 40656 18058
rect 1344 17972 40656 18006
rect 17166 17890 17218 17902
rect 17166 17826 17218 17838
rect 18846 17890 18898 17902
rect 18846 17826 18898 17838
rect 19182 17890 19234 17902
rect 19182 17826 19234 17838
rect 1934 17778 1986 17790
rect 1934 17714 1986 17726
rect 17390 17778 17442 17790
rect 17390 17714 17442 17726
rect 16606 17666 16658 17678
rect 4274 17614 4286 17666
rect 4338 17614 4350 17666
rect 16606 17602 16658 17614
rect 17054 17666 17106 17678
rect 17054 17602 17106 17614
rect 17614 17666 17666 17678
rect 21646 17666 21698 17678
rect 18834 17614 18846 17666
rect 18898 17614 18910 17666
rect 20514 17614 20526 17666
rect 20578 17614 20590 17666
rect 17614 17602 17666 17614
rect 21646 17602 21698 17614
rect 21870 17666 21922 17678
rect 21870 17602 21922 17614
rect 22542 17666 22594 17678
rect 25230 17666 25282 17678
rect 24770 17614 24782 17666
rect 24834 17614 24846 17666
rect 22542 17602 22594 17614
rect 25230 17602 25282 17614
rect 25902 17666 25954 17678
rect 25902 17602 25954 17614
rect 26238 17666 26290 17678
rect 26238 17602 26290 17614
rect 26910 17666 26962 17678
rect 26910 17602 26962 17614
rect 25678 17554 25730 17566
rect 18162 17502 18174 17554
rect 18226 17502 18238 17554
rect 19842 17502 19854 17554
rect 19906 17502 19918 17554
rect 22194 17502 22206 17554
rect 22258 17502 22270 17554
rect 24994 17502 25006 17554
rect 25058 17502 25070 17554
rect 25678 17490 25730 17502
rect 27246 17554 27298 17566
rect 27246 17490 27298 17502
rect 17726 17442 17778 17454
rect 17726 17378 17778 17390
rect 18510 17442 18562 17454
rect 18510 17378 18562 17390
rect 19518 17442 19570 17454
rect 21422 17442 21474 17454
rect 20738 17390 20750 17442
rect 20802 17390 20814 17442
rect 19518 17378 19570 17390
rect 21422 17378 21474 17390
rect 21758 17442 21810 17454
rect 21758 17378 21810 17390
rect 25454 17442 25506 17454
rect 25454 17378 25506 17390
rect 26574 17442 26626 17454
rect 26574 17378 26626 17390
rect 27022 17442 27074 17454
rect 27022 17378 27074 17390
rect 1344 17274 40656 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 40656 17274
rect 1344 17188 40656 17222
rect 15262 17106 15314 17118
rect 15262 17042 15314 17054
rect 20078 17106 20130 17118
rect 20078 17042 20130 17054
rect 16046 16994 16098 17006
rect 16046 16930 16098 16942
rect 17726 16994 17778 17006
rect 17726 16930 17778 16942
rect 19966 16994 20018 17006
rect 19966 16930 20018 16942
rect 21758 16994 21810 17006
rect 21758 16930 21810 16942
rect 21870 16994 21922 17006
rect 27346 16942 27358 16994
rect 27410 16942 27422 16994
rect 21870 16930 21922 16942
rect 17278 16882 17330 16894
rect 4274 16830 4286 16882
rect 4338 16830 4350 16882
rect 15362 16830 15374 16882
rect 15426 16830 15438 16882
rect 15810 16830 15822 16882
rect 15874 16830 15886 16882
rect 17278 16818 17330 16830
rect 17502 16882 17554 16894
rect 17502 16818 17554 16830
rect 17838 16882 17890 16894
rect 28590 16882 28642 16894
rect 28018 16830 28030 16882
rect 28082 16830 28094 16882
rect 37650 16830 37662 16882
rect 37714 16830 37726 16882
rect 17838 16818 17890 16830
rect 28590 16818 28642 16830
rect 15598 16770 15650 16782
rect 25218 16718 25230 16770
rect 25282 16718 25294 16770
rect 15598 16706 15650 16718
rect 1934 16658 1986 16670
rect 1934 16594 1986 16606
rect 21870 16658 21922 16670
rect 21870 16594 21922 16606
rect 40014 16658 40066 16670
rect 40014 16594 40066 16606
rect 1344 16490 40656 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 40656 16490
rect 1344 16404 40656 16438
rect 20302 16322 20354 16334
rect 20302 16258 20354 16270
rect 20526 16322 20578 16334
rect 20526 16258 20578 16270
rect 22206 16322 22258 16334
rect 22206 16258 22258 16270
rect 13458 16158 13470 16210
rect 13522 16158 13534 16210
rect 15586 16158 15598 16210
rect 15650 16158 15662 16210
rect 25330 16158 25342 16210
rect 25394 16158 25406 16210
rect 27458 16158 27470 16210
rect 27522 16158 27534 16210
rect 21310 16098 21362 16110
rect 16258 16046 16270 16098
rect 16322 16046 16334 16098
rect 20738 16046 20750 16098
rect 20802 16046 20814 16098
rect 21310 16034 21362 16046
rect 21646 16098 21698 16110
rect 21646 16034 21698 16046
rect 21870 16098 21922 16110
rect 21870 16034 21922 16046
rect 22318 16098 22370 16110
rect 27918 16098 27970 16110
rect 22530 16046 22542 16098
rect 22594 16046 22606 16098
rect 24546 16046 24558 16098
rect 24610 16046 24622 16098
rect 22318 16034 22370 16046
rect 27918 16034 27970 16046
rect 16830 15874 16882 15886
rect 16830 15810 16882 15822
rect 20638 15874 20690 15886
rect 20638 15810 20690 15822
rect 21646 15874 21698 15886
rect 21646 15810 21698 15822
rect 1344 15706 40656 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 40656 15706
rect 1344 15620 40656 15654
rect 15374 15538 15426 15550
rect 15374 15474 15426 15486
rect 15262 15426 15314 15438
rect 14130 15374 14142 15426
rect 14194 15374 14206 15426
rect 20962 15374 20974 15426
rect 21026 15374 21038 15426
rect 15262 15362 15314 15374
rect 23550 15314 23602 15326
rect 14914 15262 14926 15314
rect 14978 15262 14990 15314
rect 20178 15262 20190 15314
rect 20242 15262 20254 15314
rect 23550 15250 23602 15262
rect 15822 15202 15874 15214
rect 12002 15150 12014 15202
rect 12066 15150 12078 15202
rect 23090 15150 23102 15202
rect 23154 15150 23166 15202
rect 15822 15138 15874 15150
rect 1344 14922 40656 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 40656 14922
rect 1344 14836 40656 14870
rect 19182 14642 19234 14654
rect 16594 14590 16606 14642
rect 16658 14590 16670 14642
rect 18722 14590 18734 14642
rect 18786 14590 18798 14642
rect 19182 14578 19234 14590
rect 15922 14478 15934 14530
rect 15986 14478 15998 14530
rect 1344 14138 40656 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 40656 14138
rect 1344 14052 40656 14086
rect 22990 13970 23042 13982
rect 22990 13906 23042 13918
rect 20402 13806 20414 13858
rect 20466 13806 20478 13858
rect 19730 13694 19742 13746
rect 19794 13694 19806 13746
rect 22530 13582 22542 13634
rect 22594 13582 22606 13634
rect 1344 13354 40656 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 40656 13354
rect 1344 13268 40656 13302
rect 1344 12570 40656 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 40656 12570
rect 1344 12484 40656 12518
rect 1344 11786 40656 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 40656 11786
rect 1344 11700 40656 11734
rect 1344 11002 40656 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 40656 11002
rect 1344 10916 40656 10950
rect 40238 10722 40290 10734
rect 40238 10658 40290 10670
rect 1344 10218 40656 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 40656 10218
rect 1344 10132 40656 10166
rect 1344 9434 40656 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 40656 9434
rect 1344 9348 40656 9382
rect 1344 8650 40656 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 40656 8650
rect 1344 8564 40656 8598
rect 1344 7866 40656 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 40656 7866
rect 1344 7780 40656 7814
rect 1344 7082 40656 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 40656 7082
rect 1344 6996 40656 7030
rect 1344 6298 40656 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 40656 6298
rect 1344 6212 40656 6246
rect 1344 5514 40656 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 40656 5514
rect 1344 5428 40656 5462
rect 1344 4730 40656 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 40656 4730
rect 1344 4644 40656 4678
rect 1344 3946 40656 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 40656 3946
rect 1344 3860 40656 3894
rect 25566 3666 25618 3678
rect 25566 3602 25618 3614
rect 23538 3502 23550 3554
rect 23602 3502 23614 3554
rect 24546 3502 24558 3554
rect 24610 3502 24622 3554
rect 22194 3390 22206 3442
rect 22258 3390 22270 3442
rect 1344 3162 40656 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 40656 3162
rect 1344 3076 40656 3110
<< via1 >>
rect 18734 38558 18786 38610
rect 19742 38558 19794 38610
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 21758 38222 21810 38274
rect 25566 38222 25618 38274
rect 18174 38110 18226 38162
rect 19742 37998 19794 38050
rect 20750 37998 20802 38050
rect 24558 37998 24610 38050
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 20078 37438 20130 37490
rect 26238 37438 26290 37490
rect 19518 37214 19570 37266
rect 25230 37214 25282 37266
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 19742 36318 19794 36370
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 4286 27806 4338 27858
rect 1934 27582 1986 27634
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 2046 27134 2098 27186
rect 17278 27134 17330 27186
rect 4286 27022 4338 27074
rect 14366 27022 14418 27074
rect 20190 27022 20242 27074
rect 14142 26910 14194 26962
rect 19406 26910 19458 26962
rect 20638 26910 20690 26962
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 15038 26462 15090 26514
rect 19518 26462 19570 26514
rect 19854 26462 19906 26514
rect 18846 26350 18898 26402
rect 4286 26238 4338 26290
rect 14590 26238 14642 26290
rect 15262 26238 15314 26290
rect 37886 26238 37938 26290
rect 11790 26126 11842 26178
rect 13918 26126 13970 26178
rect 15934 26126 15986 26178
rect 18958 26126 19010 26178
rect 25342 26126 25394 26178
rect 39902 26126 39954 26178
rect 1934 26014 1986 26066
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 13582 25678 13634 25730
rect 2046 25566 2098 25618
rect 13470 25566 13522 25618
rect 14702 25566 14754 25618
rect 18734 25566 18786 25618
rect 19182 25566 19234 25618
rect 24782 25566 24834 25618
rect 28030 25566 28082 25618
rect 40014 25566 40066 25618
rect 4286 25454 4338 25506
rect 14366 25454 14418 25506
rect 15038 25454 15090 25506
rect 15822 25454 15874 25506
rect 19294 25454 19346 25506
rect 19518 25454 19570 25506
rect 19630 25454 19682 25506
rect 21870 25454 21922 25506
rect 25230 25454 25282 25506
rect 37662 25454 37714 25506
rect 16606 25342 16658 25394
rect 19070 25342 19122 25394
rect 19966 25342 20018 25394
rect 22654 25342 22706 25394
rect 25902 25342 25954 25394
rect 14590 25230 14642 25282
rect 14814 25230 14866 25282
rect 28478 25230 28530 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 17278 24894 17330 24946
rect 18510 24894 18562 24946
rect 23774 24894 23826 24946
rect 25790 24894 25842 24946
rect 26350 24894 26402 24946
rect 17502 24782 17554 24834
rect 18734 24782 18786 24834
rect 25566 24782 25618 24834
rect 27582 24782 27634 24834
rect 28030 24782 28082 24834
rect 13918 24670 13970 24722
rect 14254 24670 14306 24722
rect 14478 24670 14530 24722
rect 14702 24670 14754 24722
rect 14926 24670 14978 24722
rect 17614 24670 17666 24722
rect 18398 24670 18450 24722
rect 20526 24670 20578 24722
rect 25454 24670 25506 24722
rect 26126 24670 26178 24722
rect 26462 24670 26514 24722
rect 27358 24670 27410 24722
rect 27918 24670 27970 24722
rect 37662 24670 37714 24722
rect 11006 24558 11058 24610
rect 13134 24558 13186 24610
rect 14590 24558 14642 24610
rect 19070 24558 19122 24610
rect 21198 24558 21250 24610
rect 23326 24558 23378 24610
rect 28030 24446 28082 24498
rect 40014 24446 40066 24498
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 12910 24110 12962 24162
rect 12798 23998 12850 24050
rect 20414 23998 20466 24050
rect 21646 23998 21698 24050
rect 22654 23998 22706 24050
rect 28590 23998 28642 24050
rect 29262 23998 29314 24050
rect 18622 23886 18674 23938
rect 20190 23886 20242 23938
rect 20638 23886 20690 23938
rect 20750 23886 20802 23938
rect 21422 23886 21474 23938
rect 22542 23886 22594 23938
rect 23886 23886 23938 23938
rect 25678 23886 25730 23938
rect 21982 23774 22034 23826
rect 22206 23774 22258 23826
rect 22878 23774 22930 23826
rect 23438 23774 23490 23826
rect 23774 23774 23826 23826
rect 26462 23774 26514 23826
rect 14142 23662 14194 23714
rect 15598 23662 15650 23714
rect 15934 23662 15986 23714
rect 18846 23662 18898 23714
rect 21310 23662 21362 23714
rect 23662 23662 23714 23714
rect 23998 23662 24050 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 17502 23326 17554 23378
rect 17950 23326 18002 23378
rect 18062 23326 18114 23378
rect 22318 23326 22370 23378
rect 22430 23326 22482 23378
rect 22542 23326 22594 23378
rect 26462 23326 26514 23378
rect 19294 23214 19346 23266
rect 26126 23214 26178 23266
rect 26238 23214 26290 23266
rect 4286 23102 4338 23154
rect 16830 23102 16882 23154
rect 18174 23102 18226 23154
rect 18622 23102 18674 23154
rect 19070 23102 19122 23154
rect 22206 23102 22258 23154
rect 22766 23102 22818 23154
rect 13918 22990 13970 23042
rect 16046 22990 16098 23042
rect 18398 22990 18450 23042
rect 1934 22878 1986 22930
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 13582 22542 13634 22594
rect 18734 22542 18786 22594
rect 26574 22542 26626 22594
rect 1934 22430 1986 22482
rect 9998 22430 10050 22482
rect 16158 22430 16210 22482
rect 24782 22430 24834 22482
rect 25230 22430 25282 22482
rect 40014 22430 40066 22482
rect 4286 22318 4338 22370
rect 12910 22318 12962 22370
rect 13694 22318 13746 22370
rect 16942 22318 16994 22370
rect 17166 22318 17218 22370
rect 17390 22318 17442 22370
rect 17614 22318 17666 22370
rect 18734 22318 18786 22370
rect 21870 22306 21922 22358
rect 26462 22318 26514 22370
rect 37662 22318 37714 22370
rect 12126 22206 12178 22258
rect 13582 22206 13634 22258
rect 16046 22206 16098 22258
rect 16382 22206 16434 22258
rect 16606 22206 16658 22258
rect 17278 22206 17330 22258
rect 18062 22206 18114 22258
rect 19070 22206 19122 22258
rect 22654 22206 22706 22258
rect 27358 22206 27410 22258
rect 14142 22094 14194 22146
rect 18398 22094 18450 22146
rect 26574 22094 26626 22146
rect 27470 22094 27522 22146
rect 27694 22094 27746 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 13134 21758 13186 21810
rect 18398 21758 18450 21810
rect 21982 21758 22034 21810
rect 23886 21758 23938 21810
rect 24334 21758 24386 21810
rect 24558 21758 24610 21810
rect 26350 21758 26402 21810
rect 14030 21646 14082 21698
rect 20750 21646 20802 21698
rect 23438 21646 23490 21698
rect 13918 21534 13970 21586
rect 18174 21534 18226 21586
rect 20638 21534 20690 21586
rect 20974 21534 21026 21586
rect 21870 21534 21922 21586
rect 22094 21534 22146 21586
rect 22542 21534 22594 21586
rect 23662 21534 23714 21586
rect 24222 21534 24274 21586
rect 25902 21534 25954 21586
rect 29486 21534 29538 21586
rect 37886 21534 37938 21586
rect 23550 21422 23602 21474
rect 26686 21422 26738 21474
rect 28814 21422 28866 21474
rect 40014 21422 40066 21474
rect 13246 21310 13298 21362
rect 13470 21310 13522 21362
rect 25566 21310 25618 21362
rect 25902 21310 25954 21362
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 28590 20974 28642 21026
rect 16830 20862 16882 20914
rect 25230 20862 25282 20914
rect 40014 20862 40066 20914
rect 13694 20750 13746 20802
rect 20750 20750 20802 20802
rect 22654 20750 22706 20802
rect 28590 20750 28642 20802
rect 29374 20750 29426 20802
rect 29934 20750 29986 20802
rect 37662 20750 37714 20802
rect 14366 20638 14418 20690
rect 21310 20638 21362 20690
rect 28254 20638 28306 20690
rect 13470 20526 13522 20578
rect 14702 20526 14754 20578
rect 21646 20526 21698 20578
rect 29598 20526 29650 20578
rect 30270 20526 30322 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 14366 20190 14418 20242
rect 11454 20078 11506 20130
rect 14702 20078 14754 20130
rect 16382 20078 16434 20130
rect 17726 20078 17778 20130
rect 18958 20078 19010 20130
rect 21870 20078 21922 20130
rect 10782 19966 10834 20018
rect 15150 19966 15202 20018
rect 15374 19966 15426 20018
rect 16046 19966 16098 20018
rect 19294 19966 19346 20018
rect 25678 19966 25730 20018
rect 37886 19966 37938 20018
rect 13582 19854 13634 19906
rect 14030 19854 14082 19906
rect 15038 19854 15090 19906
rect 17614 19854 17666 19906
rect 26462 19854 26514 19906
rect 28590 19854 28642 19906
rect 29038 19854 29090 19906
rect 40014 19854 40066 19906
rect 17950 19742 18002 19794
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 14702 19406 14754 19458
rect 15262 19406 15314 19458
rect 19294 19406 19346 19458
rect 19630 19406 19682 19458
rect 22654 19406 22706 19458
rect 22990 19406 23042 19458
rect 40014 19406 40066 19458
rect 12910 19294 12962 19346
rect 16158 19294 16210 19346
rect 21534 19294 21586 19346
rect 21870 19294 21922 19346
rect 22430 19294 22482 19346
rect 24110 19294 24162 19346
rect 25790 19294 25842 19346
rect 26238 19294 26290 19346
rect 26462 19294 26514 19346
rect 10110 19182 10162 19234
rect 13806 19182 13858 19234
rect 15038 19182 15090 19234
rect 16494 19182 16546 19234
rect 17054 19182 17106 19234
rect 17390 19182 17442 19234
rect 19294 19182 19346 19234
rect 20190 19182 20242 19234
rect 21310 19182 21362 19234
rect 21982 19182 22034 19234
rect 24670 19182 24722 19234
rect 24894 19182 24946 19234
rect 26350 19182 26402 19234
rect 26798 19182 26850 19234
rect 27022 19182 27074 19234
rect 27358 19182 27410 19234
rect 37662 19182 37714 19234
rect 10782 19070 10834 19122
rect 14030 19070 14082 19122
rect 14478 19070 14530 19122
rect 16046 19070 16098 19122
rect 18958 19070 19010 19122
rect 20078 19070 20130 19122
rect 20302 19070 20354 19122
rect 23326 19070 23378 19122
rect 24334 19070 24386 19122
rect 25902 19070 25954 19122
rect 14590 18958 14642 19010
rect 15598 18958 15650 19010
rect 17726 18958 17778 19010
rect 21758 18958 21810 19010
rect 23438 18958 23490 19010
rect 23774 18958 23826 19010
rect 25230 18958 25282 19010
rect 25678 18958 25730 19010
rect 27246 18958 27298 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 15486 18622 15538 18674
rect 20638 18622 20690 18674
rect 15038 18510 15090 18562
rect 16270 18510 16322 18562
rect 19742 18510 19794 18562
rect 22766 18510 22818 18562
rect 23998 18510 24050 18562
rect 24110 18510 24162 18562
rect 15710 18398 15762 18450
rect 16046 18398 16098 18450
rect 16382 18398 16434 18450
rect 17390 18398 17442 18450
rect 17614 18398 17666 18450
rect 18622 18398 18674 18450
rect 18846 18398 18898 18450
rect 19966 18398 20018 18450
rect 20414 18398 20466 18450
rect 21534 18398 21586 18450
rect 21758 18398 21810 18450
rect 22430 18398 22482 18450
rect 25230 18398 25282 18450
rect 13134 18286 13186 18338
rect 14926 18286 14978 18338
rect 21310 18286 21362 18338
rect 15374 18174 15426 18226
rect 16830 18174 16882 18226
rect 17838 18174 17890 18226
rect 17950 18174 18002 18226
rect 19182 18174 19234 18226
rect 20750 18174 20802 18226
rect 22206 18174 22258 18226
rect 24110 18174 24162 18226
rect 25454 18174 25506 18226
rect 25790 18174 25842 18226
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 17166 17838 17218 17890
rect 18846 17838 18898 17890
rect 19182 17838 19234 17890
rect 1934 17726 1986 17778
rect 17390 17726 17442 17778
rect 4286 17614 4338 17666
rect 16606 17614 16658 17666
rect 17054 17614 17106 17666
rect 17614 17614 17666 17666
rect 18846 17614 18898 17666
rect 20526 17614 20578 17666
rect 21646 17614 21698 17666
rect 21870 17614 21922 17666
rect 22542 17614 22594 17666
rect 24782 17614 24834 17666
rect 25230 17614 25282 17666
rect 25902 17614 25954 17666
rect 26238 17614 26290 17666
rect 26910 17614 26962 17666
rect 18174 17502 18226 17554
rect 19854 17502 19906 17554
rect 22206 17502 22258 17554
rect 25006 17502 25058 17554
rect 25678 17502 25730 17554
rect 27246 17502 27298 17554
rect 17726 17390 17778 17442
rect 18510 17390 18562 17442
rect 19518 17390 19570 17442
rect 20750 17390 20802 17442
rect 21422 17390 21474 17442
rect 21758 17390 21810 17442
rect 25454 17390 25506 17442
rect 26574 17390 26626 17442
rect 27022 17390 27074 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 15262 17054 15314 17106
rect 20078 17054 20130 17106
rect 16046 16942 16098 16994
rect 17726 16942 17778 16994
rect 19966 16942 20018 16994
rect 21758 16942 21810 16994
rect 21870 16942 21922 16994
rect 27358 16942 27410 16994
rect 4286 16830 4338 16882
rect 15374 16830 15426 16882
rect 15822 16830 15874 16882
rect 17278 16830 17330 16882
rect 17502 16830 17554 16882
rect 17838 16830 17890 16882
rect 28030 16830 28082 16882
rect 28590 16830 28642 16882
rect 37662 16830 37714 16882
rect 15598 16718 15650 16770
rect 25230 16718 25282 16770
rect 1934 16606 1986 16658
rect 21870 16606 21922 16658
rect 40014 16606 40066 16658
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 20302 16270 20354 16322
rect 20526 16270 20578 16322
rect 22206 16270 22258 16322
rect 13470 16158 13522 16210
rect 15598 16158 15650 16210
rect 25342 16158 25394 16210
rect 27470 16158 27522 16210
rect 16270 16046 16322 16098
rect 20750 16046 20802 16098
rect 21310 16046 21362 16098
rect 21646 16046 21698 16098
rect 21870 16046 21922 16098
rect 22318 16046 22370 16098
rect 22542 16046 22594 16098
rect 24558 16046 24610 16098
rect 27918 16046 27970 16098
rect 16830 15822 16882 15874
rect 20638 15822 20690 15874
rect 21646 15822 21698 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 15374 15486 15426 15538
rect 14142 15374 14194 15426
rect 15262 15374 15314 15426
rect 20974 15374 21026 15426
rect 14926 15262 14978 15314
rect 20190 15262 20242 15314
rect 23550 15262 23602 15314
rect 12014 15150 12066 15202
rect 15822 15150 15874 15202
rect 23102 15150 23154 15202
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 16606 14590 16658 14642
rect 18734 14590 18786 14642
rect 19182 14590 19234 14642
rect 15934 14478 15986 14530
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 22990 13918 23042 13970
rect 20414 13806 20466 13858
rect 19742 13694 19794 13746
rect 22542 13582 22594 13634
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 40238 10670 40290 10722
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 25566 3614 25618 3666
rect 23550 3502 23602 3554
rect 24558 3502 24610 3554
rect 22206 3390 22258 3442
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
<< metal2 >>
rect 18144 41200 18256 42000
rect 18816 41200 18928 42000
rect 19488 41200 19600 42000
rect 20160 41200 20272 42000
rect 22848 41200 22960 42000
rect 24192 41200 24304 42000
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 18172 38162 18228 41200
rect 18172 38110 18174 38162
rect 18226 38110 18228 38162
rect 18172 38098 18228 38110
rect 18732 38610 18788 38622
rect 18732 38558 18734 38610
rect 18786 38558 18788 38610
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 4284 27860 4340 27870
rect 4284 27766 4340 27804
rect 14140 27860 14196 27870
rect 1932 27634 1988 27646
rect 1932 27582 1934 27634
rect 1986 27582 1988 27634
rect 1932 26964 1988 27582
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 1932 26898 1988 26908
rect 2044 27186 2100 27198
rect 2044 27134 2046 27186
rect 2098 27134 2100 27186
rect 2044 26292 2100 27134
rect 4284 27076 4340 27086
rect 4284 26982 4340 27020
rect 14140 26962 14196 27804
rect 17276 27186 17332 27198
rect 17276 27134 17278 27186
rect 17330 27134 17332 27186
rect 14140 26910 14142 26962
rect 14194 26910 14196 26962
rect 14140 26898 14196 26910
rect 14364 27074 14420 27086
rect 14364 27022 14366 27074
rect 14418 27022 14420 27074
rect 2044 26226 2100 26236
rect 4284 26292 4340 26302
rect 4284 26198 4340 26236
rect 11788 26292 11844 26302
rect 11788 26178 11844 26236
rect 14364 26292 14420 27022
rect 15036 27076 15092 27086
rect 15036 26514 15092 27020
rect 17276 26964 17332 27134
rect 17276 26898 17332 26908
rect 15036 26462 15038 26514
rect 15090 26462 15092 26514
rect 15036 26450 15092 26462
rect 13916 26180 13972 26190
rect 11788 26126 11790 26178
rect 11842 26126 11844 26178
rect 11788 26114 11844 26126
rect 13580 26178 13972 26180
rect 13580 26126 13918 26178
rect 13970 26126 13972 26178
rect 13580 26124 13972 26126
rect 1932 26066 1988 26078
rect 1932 26014 1934 26066
rect 1986 26014 1988 26066
rect 1932 25620 1988 26014
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 13580 25730 13636 26124
rect 13916 26114 13972 26124
rect 13580 25678 13582 25730
rect 13634 25678 13636 25730
rect 13580 25666 13636 25678
rect 1932 25554 1988 25564
rect 2044 25618 2100 25630
rect 2044 25566 2046 25618
rect 2098 25566 2100 25618
rect 2044 24948 2100 25566
rect 13468 25620 13524 25630
rect 13468 25526 13524 25564
rect 2044 24882 2100 24892
rect 4284 25506 4340 25518
rect 4284 25454 4286 25506
rect 4338 25454 4340 25506
rect 4284 24612 4340 25454
rect 13916 25508 13972 25518
rect 4284 24546 4340 24556
rect 11004 24724 11060 24734
rect 11004 24610 11060 24668
rect 13916 24722 13972 25452
rect 14364 25506 14420 26236
rect 14364 25454 14366 25506
rect 14418 25454 14420 25506
rect 14364 25442 14420 25454
rect 14588 26290 14644 26302
rect 14588 26238 14590 26290
rect 14642 26238 14644 26290
rect 14588 25508 14644 26238
rect 15260 26292 15316 26302
rect 15260 26198 15316 26236
rect 15932 26178 15988 26190
rect 15932 26126 15934 26178
rect 15986 26126 15988 26178
rect 14700 25620 14756 25630
rect 14700 25526 14756 25564
rect 14588 25442 14644 25452
rect 15036 25506 15092 25518
rect 15036 25454 15038 25506
rect 15090 25454 15092 25506
rect 14588 25284 14644 25294
rect 14476 25282 14644 25284
rect 14476 25230 14590 25282
rect 14642 25230 14644 25282
rect 14476 25228 14644 25230
rect 13916 24670 13918 24722
rect 13970 24670 13972 24722
rect 11004 24558 11006 24610
rect 11058 24558 11060 24610
rect 11004 24546 11060 24558
rect 12796 24612 12852 24622
rect 13132 24612 13188 24622
rect 4476 24332 4740 24342
rect 4172 24276 4228 24286
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 1932 22932 1988 22942
rect 1932 22838 1988 22876
rect 1932 22484 1988 22494
rect 1932 22390 1988 22428
rect 4172 20132 4228 24220
rect 12796 24050 12852 24556
rect 12908 24610 13188 24612
rect 12908 24558 13134 24610
rect 13186 24558 13188 24610
rect 12908 24556 13188 24558
rect 12908 24162 12964 24556
rect 13132 24546 13188 24556
rect 12908 24110 12910 24162
rect 12962 24110 12964 24162
rect 12908 24098 12964 24110
rect 12796 23998 12798 24050
rect 12850 23998 12852 24050
rect 12796 23986 12852 23998
rect 13916 23716 13972 24670
rect 14252 24724 14308 24734
rect 14252 24630 14308 24668
rect 14476 24722 14532 25228
rect 14588 25218 14644 25228
rect 14812 25282 14868 25294
rect 14812 25230 14814 25282
rect 14866 25230 14868 25282
rect 14476 24670 14478 24722
rect 14530 24670 14532 24722
rect 14140 23716 14196 23726
rect 13916 23714 14196 23716
rect 13916 23662 14142 23714
rect 14194 23662 14196 23714
rect 13916 23660 14196 23662
rect 4284 23156 4340 23166
rect 4284 23062 4340 23100
rect 13916 23156 13972 23166
rect 13916 23042 13972 23100
rect 13916 22990 13918 23042
rect 13970 22990 13972 23042
rect 13916 22978 13972 22990
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 13580 22596 13636 22606
rect 13580 22594 14084 22596
rect 13580 22542 13582 22594
rect 13634 22542 14084 22594
rect 13580 22540 14084 22542
rect 13580 22530 13636 22540
rect 9996 22482 10052 22494
rect 9996 22430 9998 22482
rect 10050 22430 10052 22482
rect 4284 22372 4340 22382
rect 4284 22278 4340 22316
rect 9996 22260 10052 22430
rect 12908 22370 12964 22382
rect 12908 22318 12910 22370
rect 12962 22318 12964 22370
rect 9996 22194 10052 22204
rect 12124 22258 12180 22270
rect 12124 22206 12126 22258
rect 12178 22206 12180 22258
rect 12124 21812 12180 22206
rect 12908 22148 12964 22318
rect 13692 22372 13748 22382
rect 13692 22278 13748 22316
rect 13580 22260 13636 22270
rect 13580 22166 13636 22204
rect 12908 22082 12964 22092
rect 12124 21746 12180 21756
rect 13132 21812 13188 21822
rect 13132 21718 13188 21756
rect 14028 21698 14084 22540
rect 14028 21646 14030 21698
rect 14082 21646 14084 21698
rect 14028 21634 14084 21646
rect 14140 22148 14196 23660
rect 14476 23492 14532 24670
rect 14700 24724 14756 24734
rect 14812 24724 14868 25230
rect 14700 24722 14868 24724
rect 14700 24670 14702 24722
rect 14754 24670 14868 24722
rect 14700 24668 14868 24670
rect 14700 24658 14756 24668
rect 14588 24612 14644 24622
rect 14588 24518 14644 24556
rect 14812 23716 14868 24668
rect 14812 23650 14868 23660
rect 14924 24722 14980 24734
rect 14924 24670 14926 24722
rect 14978 24670 14980 24722
rect 14924 23604 14980 24670
rect 14924 23538 14980 23548
rect 14476 23426 14532 23436
rect 15036 22260 15092 25454
rect 15820 25508 15876 25518
rect 15932 25508 15988 26126
rect 18732 25620 18788 38558
rect 18844 37492 18900 41200
rect 19516 38668 19572 41200
rect 19516 38612 19684 38668
rect 18844 37426 18900 37436
rect 19516 37266 19572 37278
rect 19516 37214 19518 37266
rect 19570 37214 19572 37266
rect 18844 26964 18900 26974
rect 19404 26962 19460 26974
rect 19404 26910 19406 26962
rect 19458 26910 19460 26962
rect 19404 26908 19460 26910
rect 18844 26402 18900 26908
rect 18844 26350 18846 26402
rect 18898 26350 18900 26402
rect 18844 26338 18900 26350
rect 19180 26852 19460 26908
rect 19516 26964 19572 37214
rect 19628 36372 19684 38612
rect 19740 38610 19796 38622
rect 19740 38558 19742 38610
rect 19794 38558 19796 38610
rect 19740 38050 19796 38558
rect 20188 38276 20244 41200
rect 20188 38210 20244 38220
rect 21756 38276 21812 38286
rect 21756 38182 21812 38220
rect 22876 38276 22932 41200
rect 22876 38210 22932 38220
rect 19740 37998 19742 38050
rect 19794 37998 19796 38050
rect 19740 37986 19796 37998
rect 20748 38050 20804 38062
rect 20748 37998 20750 38050
rect 20802 37998 20804 38050
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 20076 37492 20132 37502
rect 20076 37398 20132 37436
rect 19740 36372 19796 36382
rect 19628 36370 19796 36372
rect 19628 36318 19742 36370
rect 19794 36318 19796 36370
rect 19628 36316 19796 36318
rect 19740 36306 19796 36316
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 15876 25452 15988 25508
rect 18508 25618 18788 25620
rect 18508 25566 18734 25618
rect 18786 25566 18788 25618
rect 18508 25564 18788 25566
rect 15820 25414 15876 25452
rect 16604 25394 16660 25406
rect 16604 25342 16606 25394
rect 16658 25342 16660 25394
rect 16604 24948 16660 25342
rect 16604 24882 16660 24892
rect 17276 24948 17332 24958
rect 17276 24854 17332 24892
rect 18508 24946 18564 25564
rect 18732 25554 18788 25564
rect 18956 26178 19012 26190
rect 18956 26126 18958 26178
rect 19010 26126 19012 26178
rect 18956 25508 19012 26126
rect 19180 25618 19236 26852
rect 19516 26514 19572 26908
rect 20188 27074 20244 27086
rect 20188 27022 20190 27074
rect 20242 27022 20244 27074
rect 20188 26908 20244 27022
rect 20636 26962 20692 26974
rect 20636 26910 20638 26962
rect 20690 26910 20692 26962
rect 20636 26908 20692 26910
rect 20188 26852 20692 26908
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 19516 26462 19518 26514
rect 19570 26462 19572 26514
rect 19516 26450 19572 26462
rect 19852 26516 19908 26526
rect 19852 26422 19908 26460
rect 19180 25566 19182 25618
rect 19234 25566 19236 25618
rect 19180 25554 19236 25566
rect 18956 25442 19012 25452
rect 19292 25506 19348 25518
rect 19292 25454 19294 25506
rect 19346 25454 19348 25506
rect 18508 24894 18510 24946
rect 18562 24894 18564 24946
rect 18508 24882 18564 24894
rect 19068 25394 19124 25406
rect 19068 25342 19070 25394
rect 19122 25342 19124 25394
rect 17500 24836 17556 24846
rect 17500 24742 17556 24780
rect 18732 24836 18788 24846
rect 19068 24836 19124 25342
rect 18732 24742 18788 24780
rect 18956 24780 19124 24836
rect 17612 24724 17668 24734
rect 17612 24722 18116 24724
rect 17612 24670 17614 24722
rect 17666 24670 18116 24722
rect 17612 24668 18116 24670
rect 17612 24658 17668 24668
rect 17500 24500 17556 24510
rect 17164 24444 17500 24500
rect 15596 23716 15652 23726
rect 15596 23622 15652 23660
rect 15932 23714 15988 23726
rect 15932 23662 15934 23714
rect 15986 23662 15988 23714
rect 15036 22194 15092 22204
rect 13916 21586 13972 21598
rect 13916 21534 13918 21586
rect 13970 21534 13972 21586
rect 13244 21362 13300 21374
rect 13244 21310 13246 21362
rect 13298 21310 13300 21362
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 4172 20066 4228 20076
rect 11452 20580 11508 20590
rect 11452 20130 11508 20524
rect 11452 20078 11454 20130
rect 11506 20078 11508 20130
rect 11452 20066 11508 20078
rect 10780 20018 10836 20030
rect 10780 19966 10782 20018
rect 10834 19966 10836 20018
rect 10108 19908 10164 19918
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 10108 19234 10164 19852
rect 10780 19908 10836 19966
rect 10780 19842 10836 19852
rect 13244 19796 13300 21310
rect 13468 21362 13524 21374
rect 13468 21310 13470 21362
rect 13522 21310 13524 21362
rect 13468 20580 13524 21310
rect 13692 20804 13748 20814
rect 13468 20486 13524 20524
rect 13580 20802 13748 20804
rect 13580 20750 13694 20802
rect 13746 20750 13748 20802
rect 13580 20748 13748 20750
rect 13580 20356 13636 20748
rect 13692 20738 13748 20748
rect 13916 20692 13972 21534
rect 13916 20626 13972 20636
rect 13468 20300 13636 20356
rect 13468 20020 13524 20300
rect 13692 20244 13748 20254
rect 14140 20188 14196 22092
rect 14364 20690 14420 20702
rect 14364 20638 14366 20690
rect 14418 20638 14420 20690
rect 13468 19954 13524 19964
rect 13580 20132 13748 20188
rect 14028 20132 14196 20188
rect 14252 20244 14308 20254
rect 14364 20244 14420 20638
rect 14700 20580 14756 20590
rect 14700 20578 14868 20580
rect 14700 20526 14702 20578
rect 14754 20526 14868 20578
rect 14700 20524 14868 20526
rect 14700 20514 14756 20524
rect 14308 20242 14420 20244
rect 14308 20190 14366 20242
rect 14418 20190 14420 20242
rect 14308 20188 14420 20190
rect 14252 20178 14308 20188
rect 14364 20178 14420 20188
rect 13580 19906 13636 20132
rect 13580 19854 13582 19906
rect 13634 19854 13636 19906
rect 13580 19842 13636 19854
rect 13916 19908 13972 19918
rect 14028 19908 14084 20132
rect 14700 20130 14756 20142
rect 14700 20078 14702 20130
rect 14754 20078 14756 20130
rect 13972 19906 14084 19908
rect 13972 19854 14030 19906
rect 14082 19854 14084 19906
rect 13972 19852 14084 19854
rect 13244 19730 13300 19740
rect 12908 19348 12964 19358
rect 12908 19254 12964 19292
rect 13804 19348 13860 19358
rect 10108 19182 10110 19234
rect 10162 19182 10164 19234
rect 10108 19170 10164 19182
rect 13804 19234 13860 19292
rect 13804 19182 13806 19234
rect 13858 19182 13860 19234
rect 13804 19170 13860 19182
rect 10780 19122 10836 19134
rect 10780 19070 10782 19122
rect 10834 19070 10836 19122
rect 10780 18340 10836 19070
rect 10780 18274 10836 18284
rect 13132 18564 13188 18574
rect 13132 18338 13188 18508
rect 13916 18564 13972 19852
rect 14028 19842 14084 19852
rect 14588 19908 14644 19918
rect 14476 19348 14532 19358
rect 14028 19124 14084 19134
rect 14028 19030 14084 19068
rect 14476 19122 14532 19292
rect 14476 19070 14478 19122
rect 14530 19070 14532 19122
rect 14476 19058 14532 19070
rect 14588 19010 14644 19852
rect 14700 19684 14756 20078
rect 14700 19618 14756 19628
rect 14700 19460 14756 19470
rect 14812 19460 14868 20524
rect 15148 20020 15204 20030
rect 15148 19926 15204 19964
rect 15372 20018 15428 20030
rect 15372 19966 15374 20018
rect 15426 19966 15428 20018
rect 15036 19908 15092 19918
rect 15036 19814 15092 19852
rect 15260 19460 15316 19470
rect 14700 19458 15260 19460
rect 14700 19406 14702 19458
rect 14754 19406 15260 19458
rect 14700 19404 15260 19406
rect 14700 19394 14756 19404
rect 15260 19366 15316 19404
rect 14588 18958 14590 19010
rect 14642 18958 14644 19010
rect 14588 18788 14644 18958
rect 14588 18722 14644 18732
rect 15036 19234 15092 19246
rect 15036 19182 15038 19234
rect 15090 19182 15092 19234
rect 15036 19124 15092 19182
rect 13916 18498 13972 18508
rect 15036 18562 15092 19068
rect 15372 19012 15428 19966
rect 15932 19908 15988 23662
rect 16828 23380 16884 23390
rect 16828 23154 16884 23324
rect 16828 23102 16830 23154
rect 16882 23102 16884 23154
rect 16044 23042 16100 23054
rect 16044 22990 16046 23042
rect 16098 22990 16100 23042
rect 16044 22484 16100 22990
rect 16156 22484 16212 22494
rect 16044 22482 16212 22484
rect 16044 22430 16158 22482
rect 16210 22430 16212 22482
rect 16044 22428 16212 22430
rect 16156 22418 16212 22428
rect 16044 22260 16100 22270
rect 16044 22166 16100 22204
rect 16380 22260 16436 22270
rect 16604 22260 16660 22270
rect 16380 22258 16548 22260
rect 16380 22206 16382 22258
rect 16434 22206 16548 22258
rect 16380 22204 16548 22206
rect 16380 22194 16436 22204
rect 16492 20188 16548 22204
rect 16604 22166 16660 22204
rect 16828 20914 16884 23102
rect 16940 23156 16996 23166
rect 16940 22370 16996 23100
rect 16940 22318 16942 22370
rect 16994 22318 16996 22370
rect 16940 22306 16996 22318
rect 17164 22370 17220 24444
rect 17500 24434 17556 24444
rect 17948 23604 18004 23614
rect 17500 23380 17556 23390
rect 17500 23286 17556 23324
rect 17948 23378 18004 23548
rect 17948 23326 17950 23378
rect 18002 23326 18004 23378
rect 17948 23314 18004 23326
rect 18060 23378 18116 24668
rect 18396 24722 18452 24734
rect 18396 24670 18398 24722
rect 18450 24670 18452 24722
rect 18396 24500 18452 24670
rect 18396 24434 18452 24444
rect 18284 24052 18340 24062
rect 18172 23604 18228 23614
rect 18284 23604 18340 23996
rect 18620 23940 18676 23950
rect 18620 23938 18788 23940
rect 18620 23886 18622 23938
rect 18674 23886 18788 23938
rect 18620 23884 18788 23886
rect 18620 23874 18676 23884
rect 18228 23548 18340 23604
rect 18172 23538 18228 23548
rect 18060 23326 18062 23378
rect 18114 23326 18116 23378
rect 18060 23314 18116 23326
rect 18172 23154 18228 23166
rect 18172 23102 18174 23154
rect 18226 23102 18228 23154
rect 18172 22820 18228 23102
rect 17164 22318 17166 22370
rect 17218 22318 17220 22370
rect 16828 20862 16830 20914
rect 16882 20862 16884 20914
rect 16828 20188 16884 20862
rect 16380 20130 16436 20142
rect 16492 20132 16660 20188
rect 16828 20132 16996 20188
rect 16380 20078 16382 20130
rect 16434 20078 16436 20130
rect 15932 19842 15988 19852
rect 16044 20018 16100 20030
rect 16044 19966 16046 20018
rect 16098 19966 16100 20018
rect 16044 19348 16100 19966
rect 16380 20020 16436 20078
rect 16380 19954 16436 19964
rect 16492 19684 16548 19694
rect 16268 19460 16324 19470
rect 16044 19282 16100 19292
rect 16156 19346 16212 19358
rect 16156 19294 16158 19346
rect 16210 19294 16212 19346
rect 16044 19124 16100 19134
rect 15596 19012 15652 19022
rect 15372 19010 15652 19012
rect 15372 18958 15598 19010
rect 15650 18958 15652 19010
rect 15372 18956 15652 18958
rect 15596 18900 15652 18956
rect 15596 18834 15652 18844
rect 15484 18676 15540 18686
rect 15484 18582 15540 18620
rect 15036 18510 15038 18562
rect 15090 18510 15092 18562
rect 15036 18498 15092 18510
rect 15708 18450 15764 18462
rect 15708 18398 15710 18450
rect 15762 18398 15764 18450
rect 13132 18286 13134 18338
rect 13186 18286 13188 18338
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 1932 17780 1988 17790
rect 1932 17686 1988 17724
rect 4284 17668 4340 17678
rect 4284 17574 4340 17612
rect 4284 16884 4340 16894
rect 4284 16790 4340 16828
rect 12012 16884 12068 16894
rect 1932 16658 1988 16670
rect 1932 16606 1934 16658
rect 1986 16606 1988 16658
rect 1932 16212 1988 16606
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 1932 16146 1988 16156
rect 12012 15428 12068 16828
rect 12012 15202 12068 15372
rect 12012 15150 12014 15202
rect 12066 15150 12068 15202
rect 12012 15138 12068 15150
rect 13132 15204 13188 18286
rect 14924 18340 14980 18350
rect 14924 18246 14980 18284
rect 15372 18228 15428 18238
rect 13468 17668 13524 17678
rect 13468 16210 13524 17612
rect 13468 16158 13470 16210
rect 13522 16158 13524 16210
rect 13468 16146 13524 16158
rect 14140 17108 14196 17118
rect 14140 15426 14196 17052
rect 15260 17108 15316 17118
rect 15260 17014 15316 17052
rect 15372 16882 15428 18172
rect 15708 18004 15764 18398
rect 16044 18450 16100 19068
rect 16044 18398 16046 18450
rect 16098 18398 16100 18450
rect 16044 18386 16100 18398
rect 16156 18228 16212 19294
rect 16268 18562 16324 19404
rect 16492 19234 16548 19628
rect 16492 19182 16494 19234
rect 16546 19182 16548 19234
rect 16492 19170 16548 19182
rect 16604 19012 16660 20132
rect 16604 18946 16660 18956
rect 16268 18510 16270 18562
rect 16322 18510 16324 18562
rect 16268 18498 16324 18510
rect 16380 18452 16436 18462
rect 16380 18358 16436 18396
rect 16156 18162 16212 18172
rect 16828 18228 16884 18238
rect 16828 18134 16884 18172
rect 16940 18004 16996 20132
rect 17052 19796 17108 19806
rect 17052 19234 17108 19740
rect 17052 19182 17054 19234
rect 17106 19182 17108 19234
rect 17052 18452 17108 19182
rect 17164 18676 17220 22318
rect 17388 22764 18228 22820
rect 17388 22370 17444 22764
rect 18284 22596 18340 23548
rect 18620 23604 18676 23614
rect 18620 23154 18676 23548
rect 18620 23102 18622 23154
rect 18674 23102 18676 23154
rect 18620 23090 18676 23102
rect 18396 23044 18452 23054
rect 18396 23042 18564 23044
rect 18396 22990 18398 23042
rect 18450 22990 18564 23042
rect 18396 22988 18564 22990
rect 18396 22978 18452 22988
rect 18508 22708 18564 22988
rect 18732 22932 18788 23884
rect 18844 23716 18900 23726
rect 18844 23622 18900 23660
rect 18956 23604 19012 24780
rect 18956 23538 19012 23548
rect 19068 24610 19124 24622
rect 19068 24558 19070 24610
rect 19122 24558 19124 24610
rect 19068 23380 19124 24558
rect 19292 23492 19348 25454
rect 19516 25506 19572 25518
rect 19516 25454 19518 25506
rect 19570 25454 19572 25506
rect 19068 23314 19124 23324
rect 19180 23436 19348 23492
rect 19404 23940 19460 23950
rect 19404 23492 19460 23884
rect 19068 23154 19124 23166
rect 19068 23102 19070 23154
rect 19122 23102 19124 23154
rect 19068 22932 19124 23102
rect 18732 22876 19124 22932
rect 18732 22708 18788 22718
rect 18508 22652 18732 22708
rect 18060 22540 18340 22596
rect 18732 22594 18788 22652
rect 18732 22542 18734 22594
rect 18786 22542 18788 22594
rect 17388 22318 17390 22370
rect 17442 22318 17444 22370
rect 17276 22260 17332 22270
rect 17276 22166 17332 22204
rect 17388 20020 17444 22318
rect 17612 22370 17668 22382
rect 17612 22318 17614 22370
rect 17666 22318 17668 22370
rect 17612 21588 17668 22318
rect 18060 22258 18116 22540
rect 18732 22530 18788 22542
rect 18060 22206 18062 22258
rect 18114 22206 18116 22258
rect 18060 22194 18116 22206
rect 18732 22370 18788 22382
rect 18732 22318 18734 22370
rect 18786 22318 18788 22370
rect 18284 22148 18340 22158
rect 18284 21812 18340 22092
rect 18396 22148 18452 22158
rect 18732 22148 18788 22318
rect 18396 22146 18788 22148
rect 18396 22094 18398 22146
rect 18450 22094 18788 22146
rect 18396 22092 18788 22094
rect 18396 22082 18452 22092
rect 18396 21812 18452 21822
rect 18284 21810 18452 21812
rect 18284 21758 18398 21810
rect 18450 21758 18452 21810
rect 18284 21756 18452 21758
rect 17612 21522 17668 21532
rect 18172 21588 18228 21598
rect 18172 21494 18228 21532
rect 18284 20188 18340 21756
rect 18396 21746 18452 21756
rect 17388 19954 17444 19964
rect 17724 20130 17780 20142
rect 17724 20078 17726 20130
rect 17778 20078 17780 20130
rect 17612 19908 17668 19918
rect 17612 19814 17668 19852
rect 17724 19684 17780 20078
rect 17724 19618 17780 19628
rect 17836 20132 18340 20188
rect 17388 19460 17444 19470
rect 17388 19234 17444 19404
rect 17836 19236 17892 20132
rect 17948 19796 18004 19806
rect 17948 19702 18004 19740
rect 17388 19182 17390 19234
rect 17442 19182 17444 19234
rect 17388 19170 17444 19182
rect 17612 19180 17892 19236
rect 17164 18610 17220 18620
rect 17500 18788 17556 18798
rect 17388 18452 17444 18462
rect 17052 18386 17108 18396
rect 17276 18450 17444 18452
rect 17276 18398 17390 18450
rect 17442 18398 17444 18450
rect 17276 18396 17444 18398
rect 15708 17938 15764 17948
rect 16828 17948 16996 18004
rect 17276 18116 17332 18396
rect 17388 18386 17444 18396
rect 16604 17668 16660 17678
rect 16604 17574 16660 17612
rect 16044 17556 16100 17566
rect 15372 16830 15374 16882
rect 15426 16830 15428 16882
rect 15372 16818 15428 16830
rect 15596 16996 15652 17006
rect 15596 16770 15652 16940
rect 16044 16994 16100 17500
rect 16044 16942 16046 16994
rect 16098 16942 16100 16994
rect 16044 16930 16100 16942
rect 15596 16718 15598 16770
rect 15650 16718 15652 16770
rect 15596 16706 15652 16718
rect 15708 16884 15764 16894
rect 15596 16212 15652 16222
rect 15708 16212 15764 16828
rect 15596 16210 15764 16212
rect 15596 16158 15598 16210
rect 15650 16158 15764 16210
rect 15596 16156 15764 16158
rect 15820 16882 15876 16894
rect 15820 16830 15822 16882
rect 15874 16830 15876 16882
rect 15596 16146 15652 16156
rect 15820 15988 15876 16830
rect 16604 16324 16660 16334
rect 15372 15932 15876 15988
rect 16268 16098 16324 16110
rect 16268 16046 16270 16098
rect 16322 16046 16324 16098
rect 15372 15538 15428 15932
rect 15372 15486 15374 15538
rect 15426 15486 15428 15538
rect 15372 15474 15428 15486
rect 14140 15374 14142 15426
rect 14194 15374 14196 15426
rect 14140 15362 14196 15374
rect 15260 15428 15316 15438
rect 15260 15334 15316 15372
rect 13132 15138 13188 15148
rect 14924 15314 14980 15326
rect 14924 15262 14926 15314
rect 14978 15262 14980 15314
rect 14924 15204 14980 15262
rect 14924 15138 14980 15148
rect 15820 15204 15876 15214
rect 15932 15204 15988 15214
rect 15820 15202 15932 15204
rect 15820 15150 15822 15202
rect 15874 15150 15932 15202
rect 15820 15148 15932 15150
rect 15820 15138 15876 15148
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 15932 14530 15988 15148
rect 16268 15204 16324 16046
rect 16268 15138 16324 15148
rect 16604 14642 16660 16268
rect 16828 15874 16884 17948
rect 17164 17892 17220 17902
rect 17164 17798 17220 17836
rect 17052 17780 17108 17790
rect 17052 17666 17108 17724
rect 17052 17614 17054 17666
rect 17106 17614 17108 17666
rect 17052 17602 17108 17614
rect 17276 16882 17332 18060
rect 17388 17780 17444 17790
rect 17500 17780 17556 18732
rect 17612 18450 17668 19180
rect 17724 19012 17780 19022
rect 17724 18918 17780 18956
rect 17612 18398 17614 18450
rect 17666 18398 17668 18450
rect 17612 18386 17668 18398
rect 18172 18452 18228 18462
rect 17836 18228 17892 18238
rect 17388 17778 17556 17780
rect 17388 17726 17390 17778
rect 17442 17726 17556 17778
rect 17388 17724 17556 17726
rect 17612 18004 17668 18014
rect 17388 17714 17444 17724
rect 17612 17666 17668 17948
rect 17836 18004 17892 18172
rect 17836 17938 17892 17948
rect 17948 18226 18004 18238
rect 17948 18174 17950 18226
rect 18002 18174 18004 18226
rect 17612 17614 17614 17666
rect 17666 17614 17668 17666
rect 17612 17602 17668 17614
rect 17724 17444 17780 17454
rect 17724 17442 17892 17444
rect 17724 17390 17726 17442
rect 17778 17390 17892 17442
rect 17724 17388 17892 17390
rect 17724 17378 17780 17388
rect 17724 16996 17780 17006
rect 17724 16902 17780 16940
rect 17276 16830 17278 16882
rect 17330 16830 17332 16882
rect 17276 16818 17332 16830
rect 17500 16884 17556 16894
rect 17500 16790 17556 16828
rect 17836 16882 17892 17388
rect 17836 16830 17838 16882
rect 17890 16830 17892 16882
rect 17836 16818 17892 16830
rect 17948 16324 18004 18174
rect 18172 17554 18228 18396
rect 18620 18452 18676 18462
rect 18620 18358 18676 18396
rect 18732 17892 18788 22092
rect 19068 22258 19124 22876
rect 19068 22206 19070 22258
rect 19122 22206 19124 22258
rect 18956 20132 19012 20142
rect 18956 20038 19012 20076
rect 18956 19124 19012 19134
rect 18956 19030 19012 19068
rect 18844 18452 18900 18462
rect 18844 18358 18900 18396
rect 19068 18228 19124 22206
rect 19180 22148 19236 23436
rect 19404 23426 19460 23436
rect 19292 23268 19348 23278
rect 19292 22372 19348 23212
rect 19292 22306 19348 22316
rect 19180 22082 19236 22092
rect 19516 20188 19572 25454
rect 19628 25506 19684 25518
rect 19628 25454 19630 25506
rect 19682 25454 19684 25506
rect 19628 23716 19684 25454
rect 19852 25508 19908 25518
rect 20524 25508 20580 26852
rect 20748 26516 20804 37998
rect 24220 37492 24276 41200
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 25564 38276 25620 38286
rect 25564 38182 25620 38220
rect 24220 37426 24276 37436
rect 24556 38050 24612 38062
rect 24556 37998 24558 38050
rect 24610 37998 24612 38050
rect 20748 26450 20804 26460
rect 23884 25620 23940 25630
rect 19908 25452 20020 25508
rect 19852 25442 19908 25452
rect 19964 25394 20020 25452
rect 19964 25342 19966 25394
rect 20018 25342 20020 25394
rect 19964 25330 20020 25342
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 20524 24722 20580 25452
rect 21868 25508 21924 25518
rect 21868 25414 21924 25452
rect 23436 25508 23492 25518
rect 20524 24670 20526 24722
rect 20578 24670 20580 24722
rect 20524 24658 20580 24670
rect 22652 25394 22708 25406
rect 22652 25342 22654 25394
rect 22706 25342 22708 25394
rect 21196 24612 21252 24622
rect 21196 24610 21364 24612
rect 21196 24558 21198 24610
rect 21250 24558 21364 24610
rect 21196 24556 21364 24558
rect 21196 24546 21252 24556
rect 20412 24052 20468 24062
rect 20412 23958 20468 23996
rect 19628 23650 19684 23660
rect 20188 23940 20244 23950
rect 20636 23940 20692 23950
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 20188 23268 20244 23884
rect 20188 23202 20244 23212
rect 20524 23938 20692 23940
rect 20524 23886 20638 23938
rect 20690 23886 20692 23938
rect 20524 23884 20692 23886
rect 20524 23828 20580 23884
rect 20636 23874 20692 23884
rect 20748 23940 20804 23950
rect 20748 23846 20804 23884
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 20412 21588 20468 21598
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 19292 20132 19348 20142
rect 19516 20132 19684 20188
rect 19292 20018 19348 20076
rect 19292 19966 19294 20018
rect 19346 19966 19348 20018
rect 19292 19954 19348 19966
rect 19292 19460 19348 19470
rect 19292 19366 19348 19404
rect 19628 19458 19684 20132
rect 19628 19406 19630 19458
rect 19682 19406 19684 19458
rect 19628 19348 19684 19406
rect 19628 19282 19684 19292
rect 20188 19908 20244 19918
rect 19292 19234 19348 19246
rect 19292 19182 19294 19234
rect 19346 19182 19348 19234
rect 19292 18452 19348 19182
rect 20188 19236 20244 19852
rect 20412 19236 20468 21532
rect 20524 19460 20580 23772
rect 21308 23714 21364 24556
rect 21644 24052 21700 24062
rect 21644 23958 21700 23996
rect 22652 24050 22708 25342
rect 23436 25060 23492 25452
rect 23772 25060 23828 25070
rect 23436 25004 23772 25060
rect 23772 24946 23828 25004
rect 23772 24894 23774 24946
rect 23826 24894 23828 24946
rect 23772 24882 23828 24894
rect 22876 24612 22932 24622
rect 22652 23998 22654 24050
rect 22706 23998 22708 24050
rect 22652 23986 22708 23998
rect 22764 24556 22876 24612
rect 21308 23662 21310 23714
rect 21362 23662 21364 23714
rect 21308 23650 21364 23662
rect 21420 23938 21476 23950
rect 21420 23886 21422 23938
rect 21474 23886 21476 23938
rect 21420 23716 21476 23886
rect 22540 23940 22596 23950
rect 22540 23846 22596 23884
rect 21980 23828 22036 23838
rect 21980 23734 22036 23772
rect 22204 23828 22260 23838
rect 22204 23826 22484 23828
rect 22204 23774 22206 23826
rect 22258 23774 22484 23826
rect 22204 23772 22484 23774
rect 22204 23762 22260 23772
rect 21420 23650 21476 23660
rect 22316 23380 22372 23390
rect 21980 23378 22372 23380
rect 21980 23326 22318 23378
rect 22370 23326 22372 23378
rect 21980 23324 22372 23326
rect 20860 22708 20916 22718
rect 20748 21698 20804 21710
rect 20748 21646 20750 21698
rect 20802 21646 20804 21698
rect 20636 21588 20692 21598
rect 20636 21494 20692 21532
rect 20748 21028 20804 21646
rect 20636 20972 20804 21028
rect 20636 19908 20692 20972
rect 20748 20804 20804 20814
rect 20748 20710 20804 20748
rect 20636 19842 20692 19852
rect 20748 19460 20804 19470
rect 20524 19404 20748 19460
rect 20412 19180 20692 19236
rect 20188 19142 20244 19180
rect 20076 19122 20132 19134
rect 20076 19070 20078 19122
rect 20130 19070 20132 19122
rect 20076 19012 20132 19070
rect 20300 19122 20356 19134
rect 20300 19070 20302 19122
rect 20354 19070 20356 19122
rect 20076 18956 20244 19012
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 19292 18386 19348 18396
rect 19740 18562 19796 18574
rect 19740 18510 19742 18562
rect 19794 18510 19796 18562
rect 19740 18452 19796 18510
rect 19740 18386 19796 18396
rect 19964 18450 20020 18462
rect 19964 18398 19966 18450
rect 20018 18398 20020 18450
rect 19180 18228 19236 18238
rect 19068 18226 19236 18228
rect 19068 18174 19182 18226
rect 19234 18174 19236 18226
rect 19068 18172 19236 18174
rect 18844 17892 18900 17902
rect 18788 17890 18900 17892
rect 18788 17838 18846 17890
rect 18898 17838 18900 17890
rect 18788 17836 18900 17838
rect 18732 17798 18788 17836
rect 18844 17826 18900 17836
rect 18956 17780 19012 17790
rect 19068 17780 19124 18172
rect 19180 18162 19236 18172
rect 19852 18228 19908 18238
rect 19180 17892 19236 17902
rect 19180 17798 19236 17836
rect 19012 17724 19124 17780
rect 18956 17714 19012 17724
rect 18172 17502 18174 17554
rect 18226 17502 18228 17554
rect 18172 17490 18228 17502
rect 18844 17666 18900 17678
rect 18844 17614 18846 17666
rect 18898 17614 18900 17666
rect 17948 16258 18004 16268
rect 18508 17444 18564 17454
rect 18844 17444 18900 17614
rect 19852 17554 19908 18172
rect 19852 17502 19854 17554
rect 19906 17502 19908 17554
rect 19852 17490 19908 17502
rect 19964 17892 20020 18398
rect 19964 17556 20020 17836
rect 19964 17490 20020 17500
rect 20188 17892 20244 18956
rect 20300 18340 20356 19070
rect 20636 18674 20692 19180
rect 20636 18622 20638 18674
rect 20690 18622 20692 18674
rect 20636 18610 20692 18622
rect 20412 18564 20468 18574
rect 20412 18450 20468 18508
rect 20748 18452 20804 19404
rect 20412 18398 20414 18450
rect 20466 18398 20468 18450
rect 20412 18386 20468 18398
rect 20636 18396 20804 18452
rect 20300 18274 20356 18284
rect 20636 18116 20692 18396
rect 18508 17442 18844 17444
rect 18508 17390 18510 17442
rect 18562 17390 18844 17442
rect 18508 17388 18844 17390
rect 16828 15822 16830 15874
rect 16882 15822 16884 15874
rect 16828 15204 16884 15822
rect 16828 15138 16884 15148
rect 16604 14590 16606 14642
rect 16658 14590 16660 14642
rect 16604 14578 16660 14590
rect 18508 14644 18564 17388
rect 18844 17350 18900 17388
rect 19516 17444 19572 17454
rect 19516 17350 19572 17388
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 19964 17108 20020 17118
rect 19964 16994 20020 17052
rect 20076 17108 20132 17118
rect 20188 17108 20244 17836
rect 20076 17106 20244 17108
rect 20076 17054 20078 17106
rect 20130 17054 20244 17106
rect 20076 17052 20244 17054
rect 20300 18060 20692 18116
rect 20748 18228 20804 18238
rect 20076 17042 20132 17052
rect 19964 16942 19966 16994
rect 20018 16942 20020 16994
rect 19964 16930 20020 16942
rect 20300 16322 20356 18060
rect 20748 18004 20804 18172
rect 20524 17948 20804 18004
rect 20524 17892 20580 17948
rect 20524 17666 20580 17836
rect 20524 17614 20526 17666
rect 20578 17614 20580 17666
rect 20524 17602 20580 17614
rect 20748 17780 20804 17790
rect 20748 17442 20804 17724
rect 20748 17390 20750 17442
rect 20802 17390 20804 17442
rect 20748 17220 20804 17390
rect 20748 17154 20804 17164
rect 20300 16270 20302 16322
rect 20354 16270 20356 16322
rect 20300 16258 20356 16270
rect 20524 16324 20580 16334
rect 20860 16324 20916 22652
rect 21980 22596 22036 23324
rect 22316 23314 22372 23324
rect 22428 23378 22484 23772
rect 22764 23716 22820 24556
rect 22876 24546 22932 24556
rect 23324 24612 23380 24622
rect 23324 24518 23380 24556
rect 23884 23938 23940 25564
rect 24556 24612 24612 37998
rect 26236 37492 26292 37502
rect 26236 37398 26292 37436
rect 25228 37266 25284 37278
rect 25228 37214 25230 37266
rect 25282 37214 25284 37266
rect 25228 26852 25284 37214
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 24780 26796 25284 26852
rect 24780 25620 24836 26796
rect 37884 26290 37940 26302
rect 37884 26238 37886 26290
rect 37938 26238 37940 26290
rect 25340 26180 25396 26190
rect 24780 25526 24836 25564
rect 25228 26178 25396 26180
rect 25228 26126 25342 26178
rect 25394 26126 25396 26178
rect 25228 26124 25396 26126
rect 25228 25506 25284 26124
rect 25340 26114 25396 26124
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 25228 25454 25230 25506
rect 25282 25454 25284 25506
rect 25228 25284 25284 25454
rect 28028 25618 28084 25630
rect 28028 25566 28030 25618
rect 28082 25566 28084 25618
rect 25900 25396 25956 25406
rect 25116 25060 25172 25070
rect 25228 25060 25284 25228
rect 25788 25394 25956 25396
rect 25788 25342 25902 25394
rect 25954 25342 25956 25394
rect 25788 25340 25956 25342
rect 25172 25004 25396 25060
rect 25116 24994 25172 25004
rect 24556 24546 24612 24556
rect 25340 23940 25396 25004
rect 25788 24946 25844 25340
rect 25900 25330 25956 25340
rect 27356 25396 27412 25406
rect 25788 24894 25790 24946
rect 25842 24894 25844 24946
rect 25788 24882 25844 24894
rect 26348 24948 26404 24958
rect 26348 24854 26404 24892
rect 27356 24948 27412 25340
rect 28028 25396 28084 25566
rect 37660 25508 37716 25518
rect 37660 25414 37716 25452
rect 28028 25330 28084 25340
rect 28476 25284 28532 25294
rect 28476 25190 28532 25228
rect 25564 24836 25620 24846
rect 25564 24834 25732 24836
rect 25564 24782 25566 24834
rect 25618 24782 25732 24834
rect 25564 24780 25732 24782
rect 25564 24770 25620 24780
rect 25452 24722 25508 24734
rect 25452 24670 25454 24722
rect 25506 24670 25508 24722
rect 25452 24164 25508 24670
rect 25676 24724 25732 24780
rect 26124 24724 26180 24734
rect 26460 24724 26516 24734
rect 25676 24722 26180 24724
rect 25676 24670 26126 24722
rect 26178 24670 26180 24722
rect 25676 24668 26180 24670
rect 26124 24658 26180 24668
rect 26348 24668 26460 24724
rect 26124 24500 26180 24510
rect 25452 24108 25844 24164
rect 25676 23940 25732 23950
rect 23884 23886 23886 23938
rect 23938 23886 23940 23938
rect 23884 23874 23940 23886
rect 25228 23938 25732 23940
rect 25228 23886 25678 23938
rect 25730 23886 25732 23938
rect 25228 23884 25732 23886
rect 22876 23828 22932 23838
rect 23436 23828 23492 23838
rect 22876 23734 22932 23772
rect 23212 23826 23492 23828
rect 23212 23774 23438 23826
rect 23490 23774 23492 23826
rect 23212 23772 23492 23774
rect 22428 23326 22430 23378
rect 22482 23326 22484 23378
rect 22428 23314 22484 23326
rect 22540 23660 22820 23716
rect 22540 23378 22596 23660
rect 22540 23326 22542 23378
rect 22594 23326 22596 23378
rect 22540 23314 22596 23326
rect 22204 23156 22260 23166
rect 22764 23156 22820 23166
rect 22204 23154 22708 23156
rect 22204 23102 22206 23154
rect 22258 23102 22708 23154
rect 22204 23100 22708 23102
rect 22204 23090 22260 23100
rect 21756 22540 22036 22596
rect 21308 21700 21364 21710
rect 20972 21588 21028 21598
rect 20972 21494 21028 21532
rect 21308 20692 21364 21644
rect 21308 20598 21364 20636
rect 21644 20578 21700 20590
rect 21644 20526 21646 20578
rect 21698 20526 21700 20578
rect 21532 19796 21588 19806
rect 21420 19684 21476 19694
rect 21196 19236 21252 19246
rect 21196 17668 21252 19180
rect 21308 19234 21364 19246
rect 21308 19182 21310 19234
rect 21362 19182 21364 19234
rect 21308 18340 21364 19182
rect 21420 18452 21476 19628
rect 21532 19346 21588 19740
rect 21532 19294 21534 19346
rect 21586 19294 21588 19346
rect 21532 19282 21588 19294
rect 21532 18452 21588 18462
rect 21420 18450 21588 18452
rect 21420 18398 21534 18450
rect 21586 18398 21588 18450
rect 21420 18396 21588 18398
rect 21644 18452 21700 20526
rect 21756 19348 21812 22540
rect 22652 22484 22708 23100
rect 22764 23062 22820 23100
rect 22652 22428 22820 22484
rect 21868 22358 21924 22370
rect 21868 22306 21870 22358
rect 21922 22306 21924 22358
rect 21868 22036 21924 22306
rect 22652 22260 22708 22270
rect 21868 21970 21924 21980
rect 21980 22258 22708 22260
rect 21980 22206 22654 22258
rect 22706 22206 22708 22258
rect 21980 22204 22708 22206
rect 21980 21810 22036 22204
rect 22652 22194 22708 22204
rect 21980 21758 21982 21810
rect 22034 21758 22036 21810
rect 21980 21746 22036 21758
rect 22764 21812 22820 22428
rect 21868 21588 21924 21598
rect 21868 21494 21924 21532
rect 22092 21586 22148 21598
rect 22092 21534 22094 21586
rect 22146 21534 22148 21586
rect 21868 20804 21924 20814
rect 21868 20130 21924 20748
rect 21868 20078 21870 20130
rect 21922 20078 21924 20130
rect 21868 20066 21924 20078
rect 21980 20244 22036 20254
rect 21868 19348 21924 19358
rect 21756 19346 21924 19348
rect 21756 19294 21870 19346
rect 21922 19294 21924 19346
rect 21756 19292 21924 19294
rect 21868 19282 21924 19292
rect 21980 19234 22036 20188
rect 22092 20132 22148 21534
rect 22540 21586 22596 21598
rect 22540 21534 22542 21586
rect 22594 21534 22596 21586
rect 22540 21476 22596 21534
rect 22540 21410 22596 21420
rect 22652 20804 22708 20814
rect 22652 20710 22708 20748
rect 22148 20076 22484 20132
rect 22092 20066 22148 20076
rect 22428 19346 22484 20076
rect 22652 19684 22708 19694
rect 22652 19458 22708 19628
rect 22652 19406 22654 19458
rect 22706 19406 22708 19458
rect 22652 19394 22708 19406
rect 22428 19294 22430 19346
rect 22482 19294 22484 19346
rect 22428 19282 22484 19294
rect 21980 19182 21982 19234
rect 22034 19182 22036 19234
rect 21980 19170 22036 19182
rect 21756 19012 21812 19022
rect 21756 19010 21924 19012
rect 21756 18958 21758 19010
rect 21810 18958 21924 19010
rect 21756 18956 21924 18958
rect 21756 18946 21812 18956
rect 21756 18452 21812 18462
rect 21644 18396 21756 18452
rect 21532 18386 21588 18396
rect 21756 18358 21812 18396
rect 21868 18452 21924 18956
rect 22764 18562 22820 21756
rect 22988 21364 23044 21374
rect 22988 20244 23044 21308
rect 22988 19458 23044 20188
rect 23212 20188 23268 23772
rect 23436 23762 23492 23772
rect 23772 23828 23828 23838
rect 23772 23734 23828 23772
rect 23660 23714 23716 23726
rect 23660 23662 23662 23714
rect 23714 23662 23716 23714
rect 23660 22372 23716 23662
rect 23660 22306 23716 22316
rect 23996 23714 24052 23726
rect 23996 23662 23998 23714
rect 24050 23662 24052 23714
rect 23996 23156 24052 23662
rect 23884 21924 23940 21934
rect 23884 21810 23940 21868
rect 23884 21758 23886 21810
rect 23938 21758 23940 21810
rect 23884 21746 23940 21758
rect 23436 21700 23492 21710
rect 23436 21606 23492 21644
rect 23660 21586 23716 21598
rect 23660 21534 23662 21586
rect 23714 21534 23716 21586
rect 23548 21476 23604 21486
rect 23548 21382 23604 21420
rect 23660 20188 23716 21534
rect 23996 20188 24052 23100
rect 24556 23044 24612 23054
rect 24332 21812 24388 21822
rect 24332 21718 24388 21756
rect 24556 21810 24612 22988
rect 24780 22482 24836 22494
rect 24780 22430 24782 22482
rect 24834 22430 24836 22482
rect 24780 21924 24836 22430
rect 24780 21858 24836 21868
rect 25228 22482 25284 23884
rect 25676 23874 25732 23884
rect 25788 23044 25844 24108
rect 26124 23266 26180 24444
rect 26236 23716 26292 23726
rect 26348 23716 26404 24668
rect 26460 24630 26516 24668
rect 27356 24722 27412 24892
rect 29260 25172 29316 25182
rect 27580 24836 27636 24846
rect 27580 24742 27636 24780
rect 28028 24836 28084 24846
rect 28028 24834 28196 24836
rect 28028 24782 28030 24834
rect 28082 24782 28196 24834
rect 28028 24780 28196 24782
rect 28028 24770 28084 24780
rect 27356 24670 27358 24722
rect 27410 24670 27412 24722
rect 27356 24658 27412 24670
rect 27916 24724 27972 24734
rect 27916 24630 27972 24668
rect 28140 24612 28196 24780
rect 28140 24546 28196 24556
rect 28588 24612 28644 24622
rect 28028 24500 28084 24510
rect 28028 24406 28084 24444
rect 28588 24050 28644 24556
rect 28588 23998 28590 24050
rect 28642 23998 28644 24050
rect 28588 23986 28644 23998
rect 29260 24050 29316 25116
rect 37884 24836 37940 26238
rect 39900 26178 39956 26190
rect 39900 26126 39902 26178
rect 39954 26126 39956 26178
rect 39900 25620 39956 26126
rect 39900 25554 39956 25564
rect 40012 25618 40068 25630
rect 40012 25566 40014 25618
rect 40066 25566 40068 25618
rect 40012 24948 40068 25566
rect 40012 24882 40068 24892
rect 37884 24770 37940 24780
rect 37660 24724 37716 24734
rect 37660 24630 37716 24668
rect 40012 24498 40068 24510
rect 40012 24446 40014 24498
rect 40066 24446 40068 24498
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 40012 24276 40068 24446
rect 40012 24210 40068 24220
rect 29260 23998 29262 24050
rect 29314 23998 29316 24050
rect 29260 23986 29316 23998
rect 26292 23660 26404 23716
rect 26460 23826 26516 23838
rect 26460 23774 26462 23826
rect 26514 23774 26516 23826
rect 26236 23650 26292 23660
rect 26460 23378 26516 23774
rect 26460 23326 26462 23378
rect 26514 23326 26516 23378
rect 26460 23314 26516 23326
rect 26124 23214 26126 23266
rect 26178 23214 26180 23266
rect 26124 23202 26180 23214
rect 26236 23268 26292 23278
rect 26236 23266 26404 23268
rect 26236 23214 26238 23266
rect 26290 23214 26404 23266
rect 26236 23212 26404 23214
rect 26236 23202 26292 23212
rect 25788 22978 25844 22988
rect 26348 22708 26404 23212
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 26348 22652 26628 22708
rect 35196 22698 35460 22708
rect 26572 22594 26628 22652
rect 26572 22542 26574 22594
rect 26626 22542 26628 22594
rect 26572 22530 26628 22542
rect 25228 22430 25230 22482
rect 25282 22430 25284 22482
rect 25228 22036 25284 22430
rect 40012 22482 40068 22494
rect 40012 22430 40014 22482
rect 40066 22430 40068 22482
rect 24556 21758 24558 21810
rect 24610 21758 24612 21810
rect 24556 21746 24612 21758
rect 24220 21586 24276 21598
rect 24220 21534 24222 21586
rect 24274 21534 24276 21586
rect 24220 20188 24276 21534
rect 24444 21588 24500 21598
rect 24444 20188 24500 21532
rect 25228 20916 25284 21980
rect 25228 20822 25284 20860
rect 25452 22372 25508 22382
rect 23212 20132 23716 20188
rect 23772 20132 24052 20188
rect 24108 20132 24276 20188
rect 24332 20132 24500 20188
rect 22988 19406 22990 19458
rect 23042 19406 23044 19458
rect 22988 19394 23044 19406
rect 22764 18510 22766 18562
rect 22818 18510 22820 18562
rect 21980 18452 22036 18462
rect 21868 18396 21980 18452
rect 21308 18246 21364 18284
rect 21868 18116 21924 18396
rect 21980 18386 22036 18396
rect 22428 18450 22484 18462
rect 22428 18398 22430 18450
rect 22482 18398 22484 18450
rect 22204 18228 22260 18238
rect 21868 18050 21924 18060
rect 22092 18226 22260 18228
rect 22092 18174 22206 18226
rect 22258 18174 22260 18226
rect 22092 18172 22260 18174
rect 21644 17668 21700 17678
rect 21196 17666 21700 17668
rect 21196 17614 21646 17666
rect 21698 17614 21700 17666
rect 21196 17612 21700 17614
rect 21644 17602 21700 17612
rect 21868 17668 21924 17678
rect 21868 17574 21924 17612
rect 21420 17442 21476 17454
rect 21420 17390 21422 17442
rect 21474 17390 21476 17442
rect 21420 17220 21476 17390
rect 21420 17154 21476 17164
rect 21644 17444 21700 17454
rect 20524 16322 21364 16324
rect 20524 16270 20526 16322
rect 20578 16270 21364 16322
rect 20524 16268 21364 16270
rect 20524 16258 20580 16268
rect 20748 16100 20804 16110
rect 20748 16006 20804 16044
rect 21308 16098 21364 16268
rect 21308 16046 21310 16098
rect 21362 16046 21364 16098
rect 21308 16034 21364 16046
rect 21644 16098 21700 17388
rect 21756 17442 21812 17454
rect 21756 17390 21758 17442
rect 21810 17390 21812 17442
rect 21756 16994 21812 17390
rect 22092 17444 22148 18172
rect 22204 18162 22260 18172
rect 22428 18228 22484 18398
rect 22428 18162 22484 18172
rect 22540 18452 22596 18462
rect 22540 17666 22596 18396
rect 22540 17614 22542 17666
rect 22594 17614 22596 17666
rect 22540 17602 22596 17614
rect 22204 17556 22260 17566
rect 22204 17462 22260 17500
rect 22092 17378 22148 17388
rect 22204 17220 22260 17230
rect 21756 16942 21758 16994
rect 21810 16942 21812 16994
rect 21756 16930 21812 16942
rect 21868 16996 21924 17006
rect 21868 16994 22036 16996
rect 21868 16942 21870 16994
rect 21922 16942 22036 16994
rect 21868 16940 22036 16942
rect 21868 16930 21924 16940
rect 21644 16046 21646 16098
rect 21698 16046 21700 16098
rect 21644 16034 21700 16046
rect 21868 16658 21924 16670
rect 21868 16606 21870 16658
rect 21922 16606 21924 16658
rect 21868 16098 21924 16606
rect 21868 16046 21870 16098
rect 21922 16046 21924 16098
rect 21868 16034 21924 16046
rect 20636 15876 20692 15886
rect 20412 15874 20692 15876
rect 20412 15822 20638 15874
rect 20690 15822 20692 15874
rect 20412 15820 20692 15822
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 19628 15316 19684 15326
rect 19180 15204 19236 15214
rect 18732 14644 18788 14654
rect 18508 14642 18788 14644
rect 18508 14590 18734 14642
rect 18786 14590 18788 14642
rect 18508 14588 18788 14590
rect 18732 14578 18788 14588
rect 19180 14642 19236 15148
rect 19180 14590 19182 14642
rect 19234 14590 19236 14642
rect 19180 14578 19236 14590
rect 15932 14478 15934 14530
rect 15986 14478 15988 14530
rect 15932 14466 15988 14478
rect 19628 13748 19684 15260
rect 20188 15316 20244 15326
rect 20188 15222 20244 15260
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 20412 13858 20468 15820
rect 20636 15810 20692 15820
rect 21644 15874 21700 15886
rect 21644 15822 21646 15874
rect 21698 15822 21700 15874
rect 21644 15652 21700 15822
rect 20972 15596 21700 15652
rect 20972 15426 21028 15596
rect 20972 15374 20974 15426
rect 21026 15374 21028 15426
rect 20972 15362 21028 15374
rect 21980 15204 22036 16940
rect 22204 16322 22260 17164
rect 22764 16996 22820 18510
rect 23324 19122 23380 19134
rect 23324 19070 23326 19122
rect 23378 19070 23380 19122
rect 23324 18452 23380 19070
rect 23324 18386 23380 18396
rect 23436 19010 23492 19022
rect 23436 18958 23438 19010
rect 23490 18958 23492 19010
rect 23436 18116 23492 18958
rect 23436 17668 23492 18060
rect 23436 17602 23492 17612
rect 23548 18340 23604 20132
rect 23772 19010 23828 20132
rect 24108 19348 24164 20132
rect 23772 18958 23774 19010
rect 23826 18958 23828 19010
rect 23772 18452 23828 18958
rect 23772 18386 23828 18396
rect 23884 19346 24164 19348
rect 23884 19294 24110 19346
rect 24162 19294 24164 19346
rect 23884 19292 24164 19294
rect 23548 17556 23604 18284
rect 23772 18004 23828 18014
rect 23884 18004 23940 19292
rect 24108 19282 24164 19292
rect 23996 19124 24052 19134
rect 23996 18562 24052 19068
rect 24332 19122 24388 20132
rect 25452 19348 25508 22316
rect 26460 22372 26516 22382
rect 26460 22278 26516 22316
rect 37660 22370 37716 22382
rect 37660 22318 37662 22370
rect 37714 22318 37716 22370
rect 27356 22258 27412 22270
rect 27356 22206 27358 22258
rect 27410 22206 27412 22258
rect 26572 22146 26628 22158
rect 26572 22094 26574 22146
rect 26626 22094 26628 22146
rect 26348 22036 26404 22046
rect 26348 21810 26404 21980
rect 26348 21758 26350 21810
rect 26402 21758 26404 21810
rect 26348 21746 26404 21758
rect 25900 21588 25956 21626
rect 25900 21522 25956 21532
rect 25564 21364 25620 21374
rect 25564 21270 25620 21308
rect 25900 21362 25956 21374
rect 25900 21310 25902 21362
rect 25954 21310 25956 21362
rect 25900 21028 25956 21310
rect 25900 20962 25956 20972
rect 25676 20916 25732 20926
rect 25676 20132 25732 20860
rect 26572 20804 26628 22094
rect 27356 21700 27412 22206
rect 26684 21476 26740 21486
rect 26684 21474 26964 21476
rect 26684 21422 26686 21474
rect 26738 21422 26964 21474
rect 26684 21420 26964 21422
rect 26684 21410 26740 21420
rect 26684 21028 26740 21038
rect 26740 20972 26852 21028
rect 26684 20962 26740 20972
rect 25452 19282 25508 19292
rect 25564 20076 25732 20132
rect 24332 19070 24334 19122
rect 24386 19070 24388 19122
rect 23996 18510 23998 18562
rect 24050 18510 24052 18562
rect 23996 18498 24052 18510
rect 24108 18564 24164 18574
rect 24332 18564 24388 19070
rect 24108 18562 24388 18564
rect 24108 18510 24110 18562
rect 24162 18510 24388 18562
rect 24108 18508 24388 18510
rect 24668 19234 24724 19246
rect 24668 19182 24670 19234
rect 24722 19182 24724 19234
rect 24108 18498 24164 18508
rect 24108 18228 24164 18238
rect 24108 18134 24164 18172
rect 23828 17948 23940 18004
rect 23772 17938 23828 17948
rect 24220 17668 24276 18508
rect 24668 18340 24724 19182
rect 24892 19236 24948 19246
rect 24892 19234 25172 19236
rect 24892 19182 24894 19234
rect 24946 19182 25172 19234
rect 24892 19180 25172 19182
rect 24892 19170 24948 19180
rect 24668 18274 24724 18284
rect 24220 17602 24276 17612
rect 24780 17666 24836 17678
rect 24780 17614 24782 17666
rect 24834 17614 24836 17666
rect 23548 17490 23604 17500
rect 24780 17220 24836 17614
rect 25004 17668 25060 17678
rect 25116 17668 25172 19180
rect 25564 19124 25620 20076
rect 25676 20018 25732 20076
rect 25676 19966 25678 20018
rect 25730 19966 25732 20018
rect 25676 19954 25732 19966
rect 26348 20692 26404 20702
rect 25788 19348 25844 19358
rect 26236 19348 26292 19358
rect 25788 19346 26292 19348
rect 25788 19294 25790 19346
rect 25842 19294 26238 19346
rect 26290 19294 26292 19346
rect 25788 19292 26292 19294
rect 25788 19282 25844 19292
rect 26236 19282 26292 19292
rect 26348 19234 26404 20636
rect 26460 19906 26516 19918
rect 26460 19854 26462 19906
rect 26514 19854 26516 19906
rect 26460 19346 26516 19854
rect 26460 19294 26462 19346
rect 26514 19294 26516 19346
rect 26460 19282 26516 19294
rect 26348 19182 26350 19234
rect 26402 19182 26404 19234
rect 26348 19170 26404 19182
rect 25340 19068 25620 19124
rect 25900 19124 25956 19134
rect 25228 19012 25284 19022
rect 25228 18918 25284 18956
rect 25228 18452 25284 18462
rect 25228 18358 25284 18396
rect 25228 17668 25284 17678
rect 25116 17666 25284 17668
rect 25116 17614 25230 17666
rect 25282 17614 25284 17666
rect 25116 17612 25284 17614
rect 25004 17554 25060 17612
rect 25004 17502 25006 17554
rect 25058 17502 25060 17554
rect 25004 17490 25060 17502
rect 25228 17444 25284 17612
rect 25228 17378 25284 17388
rect 24836 17164 25284 17220
rect 24780 17126 24836 17164
rect 22764 16930 22820 16940
rect 25228 16770 25284 17164
rect 25228 16718 25230 16770
rect 25282 16718 25284 16770
rect 25228 16706 25284 16718
rect 25340 16548 25396 19068
rect 25900 19030 25956 19068
rect 25676 19012 25732 19022
rect 25676 18918 25732 18956
rect 25452 18228 25508 18238
rect 25452 18134 25508 18172
rect 25788 18228 25844 18238
rect 25788 18226 26292 18228
rect 25788 18174 25790 18226
rect 25842 18174 26292 18226
rect 25788 18172 26292 18174
rect 25788 18162 25844 18172
rect 25900 18004 25956 18014
rect 25900 17666 25956 17948
rect 25900 17614 25902 17666
rect 25954 17614 25956 17666
rect 25900 17602 25956 17614
rect 26236 17666 26292 18172
rect 26572 18004 26628 20748
rect 26796 19234 26852 20972
rect 26908 20132 26964 21420
rect 26964 20076 27076 20132
rect 26908 20066 26964 20076
rect 26796 19182 26798 19234
rect 26850 19182 26852 19234
rect 26796 19170 26852 19182
rect 27020 19234 27076 20076
rect 27020 19182 27022 19234
rect 27074 19182 27076 19234
rect 27020 19170 27076 19182
rect 27356 19234 27412 21644
rect 27468 22146 27524 22158
rect 27468 22094 27470 22146
rect 27522 22094 27524 22146
rect 27468 19908 27524 22094
rect 27692 22146 27748 22158
rect 27692 22094 27694 22146
rect 27746 22094 27748 22146
rect 27692 20692 27748 22094
rect 37660 21924 37716 22318
rect 40012 22260 40068 22430
rect 40012 22194 40068 22204
rect 37660 21858 37716 21868
rect 29484 21586 29540 21598
rect 29484 21534 29486 21586
rect 29538 21534 29540 21586
rect 28812 21476 28868 21486
rect 28588 21474 28868 21476
rect 28588 21422 28814 21474
rect 28866 21422 28868 21474
rect 28588 21420 28868 21422
rect 28588 21026 28644 21420
rect 28812 21410 28868 21420
rect 28588 20974 28590 21026
rect 28642 20974 28644 21026
rect 28588 20962 28644 20974
rect 28588 20804 28644 20814
rect 28588 20710 28644 20748
rect 29372 20804 29428 20814
rect 29372 20710 29428 20748
rect 27692 20626 27748 20636
rect 28252 20690 28308 20702
rect 28252 20638 28254 20690
rect 28306 20638 28308 20690
rect 27468 19842 27524 19852
rect 27356 19182 27358 19234
rect 27410 19182 27412 19234
rect 27356 19170 27412 19182
rect 27244 19012 27300 19022
rect 28252 19012 28308 20638
rect 29484 20188 29540 21534
rect 37884 21586 37940 21598
rect 37884 21534 37886 21586
rect 37938 21534 37940 21586
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 29932 20804 29988 20814
rect 29596 20580 29652 20590
rect 29596 20486 29652 20524
rect 29036 20132 29540 20188
rect 29932 20132 29988 20748
rect 37660 20804 37716 20814
rect 37660 20710 37716 20748
rect 30268 20580 30324 20590
rect 30268 20486 30324 20524
rect 37884 20468 37940 21534
rect 40012 21588 40068 21598
rect 40012 21474 40068 21532
rect 40012 21422 40014 21474
rect 40066 21422 40068 21474
rect 40012 21410 40068 21422
rect 40012 20916 40068 20926
rect 40012 20822 40068 20860
rect 37884 20402 37940 20412
rect 28588 19908 28644 19918
rect 28588 19814 28644 19852
rect 29036 19906 29092 20132
rect 29036 19854 29038 19906
rect 29090 19854 29092 19906
rect 27244 19010 28308 19012
rect 27244 18958 27246 19010
rect 27298 18958 28308 19010
rect 27244 18956 28308 18958
rect 27244 18946 27300 18956
rect 26572 17938 26628 17948
rect 26236 17614 26238 17666
rect 26290 17614 26292 17666
rect 26236 17602 26292 17614
rect 26908 17668 26964 17678
rect 26908 17574 26964 17612
rect 25676 17556 25732 17566
rect 25676 17462 25732 17500
rect 27244 17556 27300 17566
rect 27244 17462 27300 17500
rect 22204 16270 22206 16322
rect 22258 16270 22260 16322
rect 22204 16258 22260 16270
rect 25228 16492 25396 16548
rect 25452 17442 25508 17454
rect 25452 17390 25454 17442
rect 25506 17390 25508 17442
rect 22316 16100 22372 16110
rect 22316 16006 22372 16044
rect 22540 16098 22596 16110
rect 22540 16046 22542 16098
rect 22594 16046 22596 16098
rect 21980 15138 22036 15148
rect 20412 13806 20414 13858
rect 20466 13806 20468 13858
rect 20412 13794 20468 13806
rect 19740 13748 19796 13758
rect 19628 13746 19796 13748
rect 19628 13694 19742 13746
rect 19794 13694 19796 13746
rect 19628 13692 19796 13694
rect 19740 13682 19796 13692
rect 22540 13634 22596 16046
rect 24556 16100 24612 16110
rect 22988 15316 23044 15326
rect 22988 13970 23044 15260
rect 23548 15316 23604 15326
rect 23548 15222 23604 15260
rect 24556 15316 24612 16044
rect 25228 16100 25284 16492
rect 25340 16212 25396 16222
rect 25452 16212 25508 17390
rect 26572 17444 26628 17454
rect 26572 17350 26628 17388
rect 27020 17442 27076 17454
rect 27020 17390 27022 17442
rect 27074 17390 27076 17442
rect 27020 17332 27076 17390
rect 27020 17266 27076 17276
rect 27356 17444 27412 17454
rect 27356 16994 27412 17388
rect 27356 16942 27358 16994
rect 27410 16942 27412 16994
rect 27356 16930 27412 16942
rect 27468 17332 27524 17342
rect 25340 16210 25508 16212
rect 25340 16158 25342 16210
rect 25394 16158 25508 16210
rect 25340 16156 25508 16158
rect 27468 16210 27524 17276
rect 28028 16884 28084 16894
rect 28588 16884 28644 16894
rect 29036 16884 29092 19854
rect 29932 19124 29988 20076
rect 40012 20132 40068 20142
rect 37884 20018 37940 20030
rect 37884 19966 37886 20018
rect 37938 19966 37940 20018
rect 37660 19796 37716 19806
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 37660 19234 37716 19740
rect 37660 19182 37662 19234
rect 37714 19182 37716 19234
rect 37660 19170 37716 19182
rect 29932 19058 29988 19068
rect 37884 19124 37940 19966
rect 40012 19906 40068 20076
rect 40012 19854 40014 19906
rect 40066 19854 40068 19906
rect 40012 19842 40068 19854
rect 40012 19572 40068 19582
rect 40012 19458 40068 19516
rect 40012 19406 40014 19458
rect 40066 19406 40068 19458
rect 40012 19394 40068 19406
rect 37884 19058 37940 19068
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 27468 16158 27470 16210
rect 27522 16158 27524 16210
rect 25340 16146 25396 16156
rect 27468 16146 27524 16158
rect 27916 16882 29092 16884
rect 27916 16830 28030 16882
rect 28082 16830 28590 16882
rect 28642 16830 29092 16882
rect 27916 16828 29092 16830
rect 37660 17332 37716 17342
rect 37660 16882 37716 17276
rect 37660 16830 37662 16882
rect 37714 16830 37716 16882
rect 25228 16034 25284 16044
rect 27916 16100 27972 16828
rect 28028 16818 28084 16828
rect 28588 16818 28644 16828
rect 37660 16818 37716 16830
rect 40012 16658 40068 16670
rect 40012 16606 40014 16658
rect 40066 16606 40068 16658
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 40012 16212 40068 16606
rect 40012 16146 40068 16156
rect 27916 16006 27972 16044
rect 24556 15250 24612 15260
rect 23100 15204 23156 15214
rect 23100 15110 23156 15148
rect 24444 15204 24500 15214
rect 22988 13918 22990 13970
rect 23042 13918 23044 13970
rect 22988 13906 23044 13918
rect 22540 13582 22542 13634
rect 22594 13582 22596 13634
rect 22540 13524 22596 13582
rect 22540 13458 22596 13468
rect 23548 13524 23604 13534
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 22876 3668 22932 3678
rect 22204 3442 22260 3454
rect 22204 3390 22206 3442
rect 22258 3390 22260 3442
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 22204 800 22260 3390
rect 22876 800 22932 3612
rect 23548 3554 23604 13468
rect 24444 8428 24500 15148
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 40236 10722 40292 10734
rect 40236 10670 40238 10722
rect 40290 10670 40292 10722
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 40236 10164 40292 10670
rect 40236 10098 40292 10108
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 24444 8372 24612 8428
rect 23548 3502 23550 3554
rect 23602 3502 23604 3554
rect 23548 3490 23604 3502
rect 24556 3554 24612 8372
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 25564 3668 25620 3678
rect 25564 3574 25620 3612
rect 24556 3502 24558 3554
rect 24610 3502 24612 3554
rect 24556 3490 24612 3502
rect 22176 0 22288 800
rect 22848 0 22960 800
<< via2 >>
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 4284 27858 4340 27860
rect 4284 27806 4286 27858
rect 4286 27806 4338 27858
rect 4338 27806 4340 27858
rect 4284 27804 4340 27806
rect 14140 27804 14196 27860
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 1932 26908 1988 26964
rect 4284 27074 4340 27076
rect 4284 27022 4286 27074
rect 4286 27022 4338 27074
rect 4338 27022 4340 27074
rect 4284 27020 4340 27022
rect 2044 26236 2100 26292
rect 4284 26290 4340 26292
rect 4284 26238 4286 26290
rect 4286 26238 4338 26290
rect 4338 26238 4340 26290
rect 4284 26236 4340 26238
rect 11788 26236 11844 26292
rect 15036 27020 15092 27076
rect 17276 26908 17332 26964
rect 14364 26236 14420 26292
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 1932 25564 1988 25620
rect 13468 25618 13524 25620
rect 13468 25566 13470 25618
rect 13470 25566 13522 25618
rect 13522 25566 13524 25618
rect 13468 25564 13524 25566
rect 2044 24892 2100 24948
rect 13916 25452 13972 25508
rect 4284 24556 4340 24612
rect 11004 24668 11060 24724
rect 15260 26290 15316 26292
rect 15260 26238 15262 26290
rect 15262 26238 15314 26290
rect 15314 26238 15316 26290
rect 15260 26236 15316 26238
rect 14700 25618 14756 25620
rect 14700 25566 14702 25618
rect 14702 25566 14754 25618
rect 14754 25566 14756 25618
rect 14700 25564 14756 25566
rect 14588 25452 14644 25508
rect 12796 24556 12852 24612
rect 4476 24330 4532 24332
rect 4172 24220 4228 24276
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 1932 22930 1988 22932
rect 1932 22878 1934 22930
rect 1934 22878 1986 22930
rect 1986 22878 1988 22930
rect 1932 22876 1988 22878
rect 1932 22482 1988 22484
rect 1932 22430 1934 22482
rect 1934 22430 1986 22482
rect 1986 22430 1988 22482
rect 1932 22428 1988 22430
rect 14252 24722 14308 24724
rect 14252 24670 14254 24722
rect 14254 24670 14306 24722
rect 14306 24670 14308 24722
rect 14252 24668 14308 24670
rect 4284 23154 4340 23156
rect 4284 23102 4286 23154
rect 4286 23102 4338 23154
rect 4338 23102 4340 23154
rect 4284 23100 4340 23102
rect 13916 23100 13972 23156
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 4284 22370 4340 22372
rect 4284 22318 4286 22370
rect 4286 22318 4338 22370
rect 4338 22318 4340 22370
rect 4284 22316 4340 22318
rect 9996 22204 10052 22260
rect 13692 22370 13748 22372
rect 13692 22318 13694 22370
rect 13694 22318 13746 22370
rect 13746 22318 13748 22370
rect 13692 22316 13748 22318
rect 13580 22258 13636 22260
rect 13580 22206 13582 22258
rect 13582 22206 13634 22258
rect 13634 22206 13636 22258
rect 13580 22204 13636 22206
rect 12908 22092 12964 22148
rect 12124 21756 12180 21812
rect 13132 21810 13188 21812
rect 13132 21758 13134 21810
rect 13134 21758 13186 21810
rect 13186 21758 13188 21810
rect 13132 21756 13188 21758
rect 14588 24610 14644 24612
rect 14588 24558 14590 24610
rect 14590 24558 14642 24610
rect 14642 24558 14644 24610
rect 14588 24556 14644 24558
rect 14812 23660 14868 23716
rect 14924 23548 14980 23604
rect 14476 23436 14532 23492
rect 18844 37436 18900 37492
rect 18844 26908 18900 26964
rect 20188 38220 20244 38276
rect 21756 38274 21812 38276
rect 21756 38222 21758 38274
rect 21758 38222 21810 38274
rect 21810 38222 21812 38274
rect 21756 38220 21812 38222
rect 22876 38220 22932 38276
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 20076 37490 20132 37492
rect 20076 37438 20078 37490
rect 20078 37438 20130 37490
rect 20130 37438 20132 37490
rect 20076 37436 20132 37438
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 19516 26908 19572 26964
rect 15820 25506 15876 25508
rect 15820 25454 15822 25506
rect 15822 25454 15874 25506
rect 15874 25454 15876 25506
rect 15820 25452 15876 25454
rect 16604 24892 16660 24948
rect 17276 24946 17332 24948
rect 17276 24894 17278 24946
rect 17278 24894 17330 24946
rect 17330 24894 17332 24946
rect 17276 24892 17332 24894
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 19852 26514 19908 26516
rect 19852 26462 19854 26514
rect 19854 26462 19906 26514
rect 19906 26462 19908 26514
rect 19852 26460 19908 26462
rect 18956 25452 19012 25508
rect 17500 24834 17556 24836
rect 17500 24782 17502 24834
rect 17502 24782 17554 24834
rect 17554 24782 17556 24834
rect 17500 24780 17556 24782
rect 18732 24834 18788 24836
rect 18732 24782 18734 24834
rect 18734 24782 18786 24834
rect 18786 24782 18788 24834
rect 18732 24780 18788 24782
rect 17500 24444 17556 24500
rect 15596 23714 15652 23716
rect 15596 23662 15598 23714
rect 15598 23662 15650 23714
rect 15650 23662 15652 23714
rect 15596 23660 15652 23662
rect 15036 22204 15092 22260
rect 14140 22146 14196 22148
rect 14140 22094 14142 22146
rect 14142 22094 14194 22146
rect 14194 22094 14196 22146
rect 14140 22092 14196 22094
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 4172 20076 4228 20132
rect 11452 20524 11508 20580
rect 10108 19852 10164 19908
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 10780 19852 10836 19908
rect 13468 20578 13524 20580
rect 13468 20526 13470 20578
rect 13470 20526 13522 20578
rect 13522 20526 13524 20578
rect 13468 20524 13524 20526
rect 13916 20636 13972 20692
rect 13692 20188 13748 20244
rect 13468 19964 13524 20020
rect 14252 20188 14308 20244
rect 13916 19852 13972 19908
rect 13244 19740 13300 19796
rect 12908 19346 12964 19348
rect 12908 19294 12910 19346
rect 12910 19294 12962 19346
rect 12962 19294 12964 19346
rect 12908 19292 12964 19294
rect 13804 19292 13860 19348
rect 10780 18284 10836 18340
rect 13132 18508 13188 18564
rect 14588 19852 14644 19908
rect 14476 19292 14532 19348
rect 14028 19122 14084 19124
rect 14028 19070 14030 19122
rect 14030 19070 14082 19122
rect 14082 19070 14084 19122
rect 14028 19068 14084 19070
rect 14700 19628 14756 19684
rect 15148 20018 15204 20020
rect 15148 19966 15150 20018
rect 15150 19966 15202 20018
rect 15202 19966 15204 20018
rect 15148 19964 15204 19966
rect 15036 19906 15092 19908
rect 15036 19854 15038 19906
rect 15038 19854 15090 19906
rect 15090 19854 15092 19906
rect 15036 19852 15092 19854
rect 15260 19458 15316 19460
rect 15260 19406 15262 19458
rect 15262 19406 15314 19458
rect 15314 19406 15316 19458
rect 15260 19404 15316 19406
rect 14588 18732 14644 18788
rect 15036 19068 15092 19124
rect 13916 18508 13972 18564
rect 16828 23324 16884 23380
rect 16044 22258 16100 22260
rect 16044 22206 16046 22258
rect 16046 22206 16098 22258
rect 16098 22206 16100 22258
rect 16044 22204 16100 22206
rect 16604 22258 16660 22260
rect 16604 22206 16606 22258
rect 16606 22206 16658 22258
rect 16658 22206 16660 22258
rect 16604 22204 16660 22206
rect 16940 23100 16996 23156
rect 17948 23548 18004 23604
rect 17500 23378 17556 23380
rect 17500 23326 17502 23378
rect 17502 23326 17554 23378
rect 17554 23326 17556 23378
rect 17500 23324 17556 23326
rect 18396 24444 18452 24500
rect 18284 23996 18340 24052
rect 18172 23548 18228 23604
rect 15932 19852 15988 19908
rect 16380 19964 16436 20020
rect 16492 19628 16548 19684
rect 16268 19404 16324 19460
rect 16044 19292 16100 19348
rect 16044 19122 16100 19124
rect 16044 19070 16046 19122
rect 16046 19070 16098 19122
rect 16098 19070 16100 19122
rect 16044 19068 16100 19070
rect 15596 18844 15652 18900
rect 15484 18674 15540 18676
rect 15484 18622 15486 18674
rect 15486 18622 15538 18674
rect 15538 18622 15540 18674
rect 15484 18620 15540 18622
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 1932 17778 1988 17780
rect 1932 17726 1934 17778
rect 1934 17726 1986 17778
rect 1986 17726 1988 17778
rect 1932 17724 1988 17726
rect 4284 17666 4340 17668
rect 4284 17614 4286 17666
rect 4286 17614 4338 17666
rect 4338 17614 4340 17666
rect 4284 17612 4340 17614
rect 4284 16882 4340 16884
rect 4284 16830 4286 16882
rect 4286 16830 4338 16882
rect 4338 16830 4340 16882
rect 4284 16828 4340 16830
rect 12012 16828 12068 16884
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 1932 16156 1988 16212
rect 12012 15372 12068 15428
rect 14924 18338 14980 18340
rect 14924 18286 14926 18338
rect 14926 18286 14978 18338
rect 14978 18286 14980 18338
rect 14924 18284 14980 18286
rect 15372 18226 15428 18228
rect 15372 18174 15374 18226
rect 15374 18174 15426 18226
rect 15426 18174 15428 18226
rect 15372 18172 15428 18174
rect 13468 17612 13524 17668
rect 14140 17052 14196 17108
rect 15260 17106 15316 17108
rect 15260 17054 15262 17106
rect 15262 17054 15314 17106
rect 15314 17054 15316 17106
rect 15260 17052 15316 17054
rect 16604 18956 16660 19012
rect 16380 18450 16436 18452
rect 16380 18398 16382 18450
rect 16382 18398 16434 18450
rect 16434 18398 16436 18450
rect 16380 18396 16436 18398
rect 16156 18172 16212 18228
rect 16828 18226 16884 18228
rect 16828 18174 16830 18226
rect 16830 18174 16882 18226
rect 16882 18174 16884 18226
rect 16828 18172 16884 18174
rect 17052 19740 17108 19796
rect 18620 23548 18676 23604
rect 18844 23714 18900 23716
rect 18844 23662 18846 23714
rect 18846 23662 18898 23714
rect 18898 23662 18900 23714
rect 18844 23660 18900 23662
rect 18956 23548 19012 23604
rect 19068 23324 19124 23380
rect 19404 23884 19460 23940
rect 19404 23436 19460 23492
rect 18732 22652 18788 22708
rect 17276 22258 17332 22260
rect 17276 22206 17278 22258
rect 17278 22206 17330 22258
rect 17330 22206 17332 22258
rect 17276 22204 17332 22206
rect 18284 22092 18340 22148
rect 17612 21532 17668 21588
rect 18172 21586 18228 21588
rect 18172 21534 18174 21586
rect 18174 21534 18226 21586
rect 18226 21534 18228 21586
rect 18172 21532 18228 21534
rect 17388 19964 17444 20020
rect 17612 19906 17668 19908
rect 17612 19854 17614 19906
rect 17614 19854 17666 19906
rect 17666 19854 17668 19906
rect 17612 19852 17668 19854
rect 17724 19628 17780 19684
rect 17388 19404 17444 19460
rect 17948 19794 18004 19796
rect 17948 19742 17950 19794
rect 17950 19742 18002 19794
rect 18002 19742 18004 19794
rect 17948 19740 18004 19742
rect 17164 18620 17220 18676
rect 17500 18732 17556 18788
rect 17052 18396 17108 18452
rect 15708 17948 15764 18004
rect 17276 18060 17332 18116
rect 16604 17666 16660 17668
rect 16604 17614 16606 17666
rect 16606 17614 16658 17666
rect 16658 17614 16660 17666
rect 16604 17612 16660 17614
rect 16044 17500 16100 17556
rect 15596 16940 15652 16996
rect 15708 16828 15764 16884
rect 16604 16268 16660 16324
rect 15260 15426 15316 15428
rect 15260 15374 15262 15426
rect 15262 15374 15314 15426
rect 15314 15374 15316 15426
rect 15260 15372 15316 15374
rect 13132 15148 13188 15204
rect 14924 15148 14980 15204
rect 15932 15148 15988 15204
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 16268 15148 16324 15204
rect 17164 17890 17220 17892
rect 17164 17838 17166 17890
rect 17166 17838 17218 17890
rect 17218 17838 17220 17890
rect 17164 17836 17220 17838
rect 17052 17724 17108 17780
rect 17724 19010 17780 19012
rect 17724 18958 17726 19010
rect 17726 18958 17778 19010
rect 17778 18958 17780 19010
rect 17724 18956 17780 18958
rect 18172 18396 18228 18452
rect 17836 18226 17892 18228
rect 17836 18174 17838 18226
rect 17838 18174 17890 18226
rect 17890 18174 17892 18226
rect 17836 18172 17892 18174
rect 17612 17948 17668 18004
rect 17836 17948 17892 18004
rect 17724 16994 17780 16996
rect 17724 16942 17726 16994
rect 17726 16942 17778 16994
rect 17778 16942 17780 16994
rect 17724 16940 17780 16942
rect 17500 16882 17556 16884
rect 17500 16830 17502 16882
rect 17502 16830 17554 16882
rect 17554 16830 17556 16882
rect 17500 16828 17556 16830
rect 18620 18450 18676 18452
rect 18620 18398 18622 18450
rect 18622 18398 18674 18450
rect 18674 18398 18676 18450
rect 18620 18396 18676 18398
rect 18956 20130 19012 20132
rect 18956 20078 18958 20130
rect 18958 20078 19010 20130
rect 19010 20078 19012 20130
rect 18956 20076 19012 20078
rect 18956 19122 19012 19124
rect 18956 19070 18958 19122
rect 18958 19070 19010 19122
rect 19010 19070 19012 19122
rect 18956 19068 19012 19070
rect 18844 18450 18900 18452
rect 18844 18398 18846 18450
rect 18846 18398 18898 18450
rect 18898 18398 18900 18450
rect 18844 18396 18900 18398
rect 19292 23266 19348 23268
rect 19292 23214 19294 23266
rect 19294 23214 19346 23266
rect 19346 23214 19348 23266
rect 19292 23212 19348 23214
rect 19292 22316 19348 22372
rect 19180 22092 19236 22148
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 25564 38274 25620 38276
rect 25564 38222 25566 38274
rect 25566 38222 25618 38274
rect 25618 38222 25620 38274
rect 25564 38220 25620 38222
rect 24220 37436 24276 37492
rect 20748 26460 20804 26516
rect 23884 25564 23940 25620
rect 19852 25452 19908 25508
rect 20524 25452 20580 25508
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 21868 25506 21924 25508
rect 21868 25454 21870 25506
rect 21870 25454 21922 25506
rect 21922 25454 21924 25506
rect 21868 25452 21924 25454
rect 23436 25452 23492 25508
rect 20412 24050 20468 24052
rect 20412 23998 20414 24050
rect 20414 23998 20466 24050
rect 20466 23998 20468 24050
rect 20412 23996 20468 23998
rect 19628 23660 19684 23716
rect 20188 23938 20244 23940
rect 20188 23886 20190 23938
rect 20190 23886 20242 23938
rect 20242 23886 20244 23938
rect 20188 23884 20244 23886
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 20188 23212 20244 23268
rect 20748 23938 20804 23940
rect 20748 23886 20750 23938
rect 20750 23886 20802 23938
rect 20802 23886 20804 23938
rect 20748 23884 20804 23886
rect 20524 23772 20580 23828
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 20412 21532 20468 21588
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 19292 20076 19348 20132
rect 19292 19458 19348 19460
rect 19292 19406 19294 19458
rect 19294 19406 19346 19458
rect 19346 19406 19348 19458
rect 19292 19404 19348 19406
rect 19628 19292 19684 19348
rect 20188 19852 20244 19908
rect 20188 19234 20244 19236
rect 20188 19182 20190 19234
rect 20190 19182 20242 19234
rect 20242 19182 20244 19234
rect 20188 19180 20244 19182
rect 21644 24050 21700 24052
rect 21644 23998 21646 24050
rect 21646 23998 21698 24050
rect 21698 23998 21700 24050
rect 21644 23996 21700 23998
rect 23772 25004 23828 25060
rect 22876 24556 22932 24612
rect 22540 23938 22596 23940
rect 22540 23886 22542 23938
rect 22542 23886 22594 23938
rect 22594 23886 22596 23938
rect 22540 23884 22596 23886
rect 21980 23826 22036 23828
rect 21980 23774 21982 23826
rect 21982 23774 22034 23826
rect 22034 23774 22036 23826
rect 21980 23772 22036 23774
rect 21420 23660 21476 23716
rect 20860 22652 20916 22708
rect 20636 21586 20692 21588
rect 20636 21534 20638 21586
rect 20638 21534 20690 21586
rect 20690 21534 20692 21586
rect 20636 21532 20692 21534
rect 20748 20802 20804 20804
rect 20748 20750 20750 20802
rect 20750 20750 20802 20802
rect 20802 20750 20804 20802
rect 20748 20748 20804 20750
rect 20636 19852 20692 19908
rect 20748 19404 20804 19460
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 19292 18396 19348 18452
rect 19740 18396 19796 18452
rect 18732 17836 18788 17892
rect 19852 18172 19908 18228
rect 19180 17890 19236 17892
rect 19180 17838 19182 17890
rect 19182 17838 19234 17890
rect 19234 17838 19236 17890
rect 19180 17836 19236 17838
rect 18956 17724 19012 17780
rect 17948 16268 18004 16324
rect 19964 17836 20020 17892
rect 19964 17500 20020 17556
rect 20412 18508 20468 18564
rect 20300 18284 20356 18340
rect 20188 17836 20244 17892
rect 18844 17388 18900 17444
rect 16828 15148 16884 15204
rect 19516 17442 19572 17444
rect 19516 17390 19518 17442
rect 19518 17390 19570 17442
rect 19570 17390 19572 17442
rect 19516 17388 19572 17390
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 19964 17052 20020 17108
rect 20748 18226 20804 18228
rect 20748 18174 20750 18226
rect 20750 18174 20802 18226
rect 20802 18174 20804 18226
rect 20748 18172 20804 18174
rect 20524 17836 20580 17892
rect 20748 17724 20804 17780
rect 20748 17164 20804 17220
rect 23324 24610 23380 24612
rect 23324 24558 23326 24610
rect 23326 24558 23378 24610
rect 23378 24558 23380 24610
rect 23324 24556 23380 24558
rect 26236 37490 26292 37492
rect 26236 37438 26238 37490
rect 26238 37438 26290 37490
rect 26290 37438 26292 37490
rect 26236 37436 26292 37438
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 24780 25618 24836 25620
rect 24780 25566 24782 25618
rect 24782 25566 24834 25618
rect 24834 25566 24836 25618
rect 24780 25564 24836 25566
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 25228 25228 25284 25284
rect 25116 25004 25172 25060
rect 24556 24556 24612 24612
rect 27356 25340 27412 25396
rect 26348 24946 26404 24948
rect 26348 24894 26350 24946
rect 26350 24894 26402 24946
rect 26402 24894 26404 24946
rect 26348 24892 26404 24894
rect 37660 25506 37716 25508
rect 37660 25454 37662 25506
rect 37662 25454 37714 25506
rect 37714 25454 37716 25506
rect 37660 25452 37716 25454
rect 28028 25340 28084 25396
rect 28476 25282 28532 25284
rect 28476 25230 28478 25282
rect 28478 25230 28530 25282
rect 28530 25230 28532 25282
rect 28476 25228 28532 25230
rect 27356 24892 27412 24948
rect 26460 24722 26516 24724
rect 26460 24670 26462 24722
rect 26462 24670 26514 24722
rect 26514 24670 26516 24722
rect 26460 24668 26516 24670
rect 26124 24444 26180 24500
rect 22876 23826 22932 23828
rect 22876 23774 22878 23826
rect 22878 23774 22930 23826
rect 22930 23774 22932 23826
rect 22876 23772 22932 23774
rect 21308 21644 21364 21700
rect 20972 21586 21028 21588
rect 20972 21534 20974 21586
rect 20974 21534 21026 21586
rect 21026 21534 21028 21586
rect 20972 21532 21028 21534
rect 21308 20690 21364 20692
rect 21308 20638 21310 20690
rect 21310 20638 21362 20690
rect 21362 20638 21364 20690
rect 21308 20636 21364 20638
rect 21532 19740 21588 19796
rect 21420 19628 21476 19684
rect 21196 19180 21252 19236
rect 22764 23154 22820 23156
rect 22764 23102 22766 23154
rect 22766 23102 22818 23154
rect 22818 23102 22820 23154
rect 22764 23100 22820 23102
rect 21868 21980 21924 22036
rect 22764 21756 22820 21812
rect 21868 21586 21924 21588
rect 21868 21534 21870 21586
rect 21870 21534 21922 21586
rect 21922 21534 21924 21586
rect 21868 21532 21924 21534
rect 21868 20748 21924 20804
rect 21980 20188 22036 20244
rect 22540 21420 22596 21476
rect 22652 20802 22708 20804
rect 22652 20750 22654 20802
rect 22654 20750 22706 20802
rect 22706 20750 22708 20802
rect 22652 20748 22708 20750
rect 22092 20076 22148 20132
rect 22652 19628 22708 19684
rect 21756 18450 21812 18452
rect 21756 18398 21758 18450
rect 21758 18398 21810 18450
rect 21810 18398 21812 18450
rect 21756 18396 21812 18398
rect 22988 21308 23044 21364
rect 22988 20188 23044 20244
rect 23772 23826 23828 23828
rect 23772 23774 23774 23826
rect 23774 23774 23826 23826
rect 23826 23774 23828 23826
rect 23772 23772 23828 23774
rect 23660 22316 23716 22372
rect 23996 23100 24052 23156
rect 23884 21868 23940 21924
rect 23436 21698 23492 21700
rect 23436 21646 23438 21698
rect 23438 21646 23490 21698
rect 23490 21646 23492 21698
rect 23436 21644 23492 21646
rect 23548 21474 23604 21476
rect 23548 21422 23550 21474
rect 23550 21422 23602 21474
rect 23602 21422 23604 21474
rect 23548 21420 23604 21422
rect 24556 22988 24612 23044
rect 24332 21810 24388 21812
rect 24332 21758 24334 21810
rect 24334 21758 24386 21810
rect 24386 21758 24388 21810
rect 24332 21756 24388 21758
rect 24780 21868 24836 21924
rect 29260 25116 29316 25172
rect 27580 24834 27636 24836
rect 27580 24782 27582 24834
rect 27582 24782 27634 24834
rect 27634 24782 27636 24834
rect 27580 24780 27636 24782
rect 27916 24722 27972 24724
rect 27916 24670 27918 24722
rect 27918 24670 27970 24722
rect 27970 24670 27972 24722
rect 27916 24668 27972 24670
rect 28140 24556 28196 24612
rect 28588 24556 28644 24612
rect 28028 24498 28084 24500
rect 28028 24446 28030 24498
rect 28030 24446 28082 24498
rect 28082 24446 28084 24498
rect 28028 24444 28084 24446
rect 39900 25564 39956 25620
rect 40012 24892 40068 24948
rect 37884 24780 37940 24836
rect 37660 24722 37716 24724
rect 37660 24670 37662 24722
rect 37662 24670 37714 24722
rect 37714 24670 37716 24722
rect 37660 24668 37716 24670
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 40012 24220 40068 24276
rect 26236 23660 26292 23716
rect 25788 22988 25844 23044
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 25228 21980 25284 22036
rect 24444 21532 24500 21588
rect 25228 20914 25284 20916
rect 25228 20862 25230 20914
rect 25230 20862 25282 20914
rect 25282 20862 25284 20914
rect 25228 20860 25284 20862
rect 25452 22316 25508 22372
rect 21980 18396 22036 18452
rect 21308 18338 21364 18340
rect 21308 18286 21310 18338
rect 21310 18286 21362 18338
rect 21362 18286 21364 18338
rect 21308 18284 21364 18286
rect 21868 18060 21924 18116
rect 21868 17666 21924 17668
rect 21868 17614 21870 17666
rect 21870 17614 21922 17666
rect 21922 17614 21924 17666
rect 21868 17612 21924 17614
rect 21420 17164 21476 17220
rect 21644 17388 21700 17444
rect 20748 16098 20804 16100
rect 20748 16046 20750 16098
rect 20750 16046 20802 16098
rect 20802 16046 20804 16098
rect 20748 16044 20804 16046
rect 22428 18172 22484 18228
rect 22540 18396 22596 18452
rect 22204 17554 22260 17556
rect 22204 17502 22206 17554
rect 22206 17502 22258 17554
rect 22258 17502 22260 17554
rect 22204 17500 22260 17502
rect 22092 17388 22148 17444
rect 22204 17164 22260 17220
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 19628 15260 19684 15316
rect 19180 15148 19236 15204
rect 20188 15314 20244 15316
rect 20188 15262 20190 15314
rect 20190 15262 20242 15314
rect 20242 15262 20244 15314
rect 20188 15260 20244 15262
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 23324 18396 23380 18452
rect 23436 18060 23492 18116
rect 23436 17612 23492 17668
rect 23772 18396 23828 18452
rect 23548 18284 23604 18340
rect 23996 19068 24052 19124
rect 26460 22370 26516 22372
rect 26460 22318 26462 22370
rect 26462 22318 26514 22370
rect 26514 22318 26516 22370
rect 26460 22316 26516 22318
rect 26348 21980 26404 22036
rect 25900 21586 25956 21588
rect 25900 21534 25902 21586
rect 25902 21534 25954 21586
rect 25954 21534 25956 21586
rect 25900 21532 25956 21534
rect 25564 21362 25620 21364
rect 25564 21310 25566 21362
rect 25566 21310 25618 21362
rect 25618 21310 25620 21362
rect 25564 21308 25620 21310
rect 25900 20972 25956 21028
rect 25676 20860 25732 20916
rect 27356 21644 27412 21700
rect 26684 20972 26740 21028
rect 26572 20748 26628 20804
rect 25452 19292 25508 19348
rect 24108 18226 24164 18228
rect 24108 18174 24110 18226
rect 24110 18174 24162 18226
rect 24162 18174 24164 18226
rect 24108 18172 24164 18174
rect 23772 17948 23828 18004
rect 24668 18284 24724 18340
rect 24220 17612 24276 17668
rect 23548 17500 23604 17556
rect 25004 17612 25060 17668
rect 26348 20636 26404 20692
rect 25900 19122 25956 19124
rect 25900 19070 25902 19122
rect 25902 19070 25954 19122
rect 25954 19070 25956 19122
rect 25900 19068 25956 19070
rect 25228 19010 25284 19012
rect 25228 18958 25230 19010
rect 25230 18958 25282 19010
rect 25282 18958 25284 19010
rect 25228 18956 25284 18958
rect 25228 18450 25284 18452
rect 25228 18398 25230 18450
rect 25230 18398 25282 18450
rect 25282 18398 25284 18450
rect 25228 18396 25284 18398
rect 25228 17388 25284 17444
rect 24780 17164 24836 17220
rect 22764 16940 22820 16996
rect 25676 19010 25732 19012
rect 25676 18958 25678 19010
rect 25678 18958 25730 19010
rect 25730 18958 25732 19010
rect 25676 18956 25732 18958
rect 25452 18226 25508 18228
rect 25452 18174 25454 18226
rect 25454 18174 25506 18226
rect 25506 18174 25508 18226
rect 25452 18172 25508 18174
rect 25900 17948 25956 18004
rect 26908 20076 26964 20132
rect 40012 22204 40068 22260
rect 37660 21868 37716 21924
rect 28588 20802 28644 20804
rect 28588 20750 28590 20802
rect 28590 20750 28642 20802
rect 28642 20750 28644 20802
rect 28588 20748 28644 20750
rect 29372 20802 29428 20804
rect 29372 20750 29374 20802
rect 29374 20750 29426 20802
rect 29426 20750 29428 20802
rect 29372 20748 29428 20750
rect 27692 20636 27748 20692
rect 27468 19852 27524 19908
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 29932 20802 29988 20804
rect 29932 20750 29934 20802
rect 29934 20750 29986 20802
rect 29986 20750 29988 20802
rect 29932 20748 29988 20750
rect 29596 20578 29652 20580
rect 29596 20526 29598 20578
rect 29598 20526 29650 20578
rect 29650 20526 29652 20578
rect 29596 20524 29652 20526
rect 37660 20802 37716 20804
rect 37660 20750 37662 20802
rect 37662 20750 37714 20802
rect 37714 20750 37716 20802
rect 37660 20748 37716 20750
rect 30268 20578 30324 20580
rect 30268 20526 30270 20578
rect 30270 20526 30322 20578
rect 30322 20526 30324 20578
rect 30268 20524 30324 20526
rect 40012 21532 40068 21588
rect 40012 20914 40068 20916
rect 40012 20862 40014 20914
rect 40014 20862 40066 20914
rect 40066 20862 40068 20914
rect 40012 20860 40068 20862
rect 37884 20412 37940 20468
rect 28588 19906 28644 19908
rect 28588 19854 28590 19906
rect 28590 19854 28642 19906
rect 28642 19854 28644 19906
rect 28588 19852 28644 19854
rect 26572 17948 26628 18004
rect 26908 17666 26964 17668
rect 26908 17614 26910 17666
rect 26910 17614 26962 17666
rect 26962 17614 26964 17666
rect 26908 17612 26964 17614
rect 25676 17554 25732 17556
rect 25676 17502 25678 17554
rect 25678 17502 25730 17554
rect 25730 17502 25732 17554
rect 25676 17500 25732 17502
rect 27244 17554 27300 17556
rect 27244 17502 27246 17554
rect 27246 17502 27298 17554
rect 27298 17502 27300 17554
rect 27244 17500 27300 17502
rect 22316 16098 22372 16100
rect 22316 16046 22318 16098
rect 22318 16046 22370 16098
rect 22370 16046 22372 16098
rect 22316 16044 22372 16046
rect 21980 15148 22036 15204
rect 24556 16098 24612 16100
rect 24556 16046 24558 16098
rect 24558 16046 24610 16098
rect 24610 16046 24612 16098
rect 24556 16044 24612 16046
rect 22988 15260 23044 15316
rect 23548 15314 23604 15316
rect 23548 15262 23550 15314
rect 23550 15262 23602 15314
rect 23602 15262 23604 15314
rect 23548 15260 23604 15262
rect 26572 17442 26628 17444
rect 26572 17390 26574 17442
rect 26574 17390 26626 17442
rect 26626 17390 26628 17442
rect 26572 17388 26628 17390
rect 27020 17276 27076 17332
rect 27356 17388 27412 17444
rect 27468 17276 27524 17332
rect 29932 20076 29988 20132
rect 40012 20076 40068 20132
rect 37660 19740 37716 19796
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 29932 19068 29988 19124
rect 40012 19516 40068 19572
rect 37884 19068 37940 19124
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 37660 17276 37716 17332
rect 25228 16044 25284 16100
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 40012 16156 40068 16212
rect 27916 16098 27972 16100
rect 27916 16046 27918 16098
rect 27918 16046 27970 16098
rect 27970 16046 27972 16098
rect 27916 16044 27972 16046
rect 24556 15260 24612 15316
rect 23100 15202 23156 15204
rect 23100 15150 23102 15202
rect 23102 15150 23154 15202
rect 23154 15150 23156 15202
rect 23100 15148 23156 15150
rect 24444 15148 24500 15204
rect 22540 13468 22596 13524
rect 23548 13468 23604 13524
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 22876 3612 22932 3668
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 40236 10108 40292 10164
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 25564 3666 25620 3668
rect 25564 3614 25566 3666
rect 25566 3614 25618 3666
rect 25618 3614 25620 3666
rect 25564 3612 25620 3614
<< metal3 >>
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 20178 38220 20188 38276
rect 20244 38220 21756 38276
rect 21812 38220 21822 38276
rect 22866 38220 22876 38276
rect 22932 38220 25564 38276
rect 25620 38220 25630 38276
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 18834 37436 18844 37492
rect 18900 37436 20076 37492
rect 20132 37436 20142 37492
rect 24210 37436 24220 37492
rect 24276 37436 26236 37492
rect 26292 37436 26302 37492
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 4274 27804 4284 27860
rect 4340 27804 14140 27860
rect 14196 27804 14206 27860
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 4274 27020 4284 27076
rect 4340 27020 15036 27076
rect 15092 27020 15102 27076
rect 0 26964 800 26992
rect 0 26908 1932 26964
rect 1988 26908 1998 26964
rect 17266 26908 17276 26964
rect 17332 26908 18844 26964
rect 18900 26908 19516 26964
rect 19572 26908 19582 26964
rect 0 26880 800 26908
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 19842 26460 19852 26516
rect 19908 26460 20748 26516
rect 20804 26460 20814 26516
rect 0 26292 800 26320
rect 0 26236 2044 26292
rect 2100 26236 2110 26292
rect 4274 26236 4284 26292
rect 4340 26236 11788 26292
rect 11844 26236 14364 26292
rect 14420 26236 15260 26292
rect 15316 26236 15326 26292
rect 0 26208 800 26236
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 0 25620 800 25648
rect 41200 25620 42000 25648
rect 0 25564 1932 25620
rect 1988 25564 1998 25620
rect 13458 25564 13468 25620
rect 13524 25564 14700 25620
rect 14756 25564 14766 25620
rect 23874 25564 23884 25620
rect 23940 25564 24780 25620
rect 24836 25564 24846 25620
rect 39890 25564 39900 25620
rect 39956 25564 42000 25620
rect 0 25536 800 25564
rect 41200 25536 42000 25564
rect 13906 25452 13916 25508
rect 13972 25452 14588 25508
rect 14644 25452 15820 25508
rect 15876 25452 15886 25508
rect 18946 25452 18956 25508
rect 19012 25452 19852 25508
rect 19908 25452 19918 25508
rect 20514 25452 20524 25508
rect 20580 25452 21868 25508
rect 21924 25452 23436 25508
rect 23492 25452 23502 25508
rect 31892 25452 37660 25508
rect 37716 25452 37726 25508
rect 31892 25396 31948 25452
rect 27346 25340 27356 25396
rect 27412 25340 28028 25396
rect 28084 25340 31948 25396
rect 25218 25228 25228 25284
rect 25284 25228 28476 25284
rect 28532 25228 28542 25284
rect 28476 25172 28532 25228
rect 28476 25116 29260 25172
rect 29316 25116 29326 25172
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 23762 25004 23772 25060
rect 23828 25004 25116 25060
rect 25172 25004 25182 25060
rect 0 24948 800 24976
rect 41200 24948 42000 24976
rect 0 24892 2044 24948
rect 2100 24892 2110 24948
rect 16594 24892 16604 24948
rect 16660 24892 17276 24948
rect 17332 24892 17342 24948
rect 26338 24892 26348 24948
rect 26404 24892 27356 24948
rect 27412 24892 27422 24948
rect 40002 24892 40012 24948
rect 40068 24892 42000 24948
rect 0 24864 800 24892
rect 41200 24864 42000 24892
rect 17490 24780 17500 24836
rect 17556 24780 18732 24836
rect 18788 24780 18798 24836
rect 27570 24780 27580 24836
rect 27636 24780 37884 24836
rect 37940 24780 37950 24836
rect 8372 24668 11004 24724
rect 11060 24668 14252 24724
rect 14308 24668 14318 24724
rect 26450 24668 26460 24724
rect 26516 24668 27916 24724
rect 27972 24668 27982 24724
rect 31892 24668 37660 24724
rect 37716 24668 37726 24724
rect 8372 24612 8428 24668
rect 31892 24612 31948 24668
rect 4274 24556 4284 24612
rect 4340 24556 8428 24612
rect 12786 24556 12796 24612
rect 12852 24556 14588 24612
rect 14644 24556 14654 24612
rect 22866 24556 22876 24612
rect 22932 24556 23324 24612
rect 23380 24556 24556 24612
rect 24612 24556 24622 24612
rect 28130 24556 28140 24612
rect 28196 24556 28588 24612
rect 28644 24556 31948 24612
rect 17490 24444 17500 24500
rect 17556 24444 18396 24500
rect 18452 24444 18462 24500
rect 26114 24444 26124 24500
rect 26180 24444 28028 24500
rect 28084 24444 28094 24500
rect 0 24276 800 24304
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 41200 24276 42000 24304
rect 0 24220 4172 24276
rect 4228 24220 4238 24276
rect 40002 24220 40012 24276
rect 40068 24220 42000 24276
rect 0 24192 800 24220
rect 41200 24192 42000 24220
rect 18274 23996 18284 24052
rect 18340 23996 20412 24052
rect 20468 23996 21644 24052
rect 21700 23996 21710 24052
rect 19394 23884 19404 23940
rect 19460 23884 20188 23940
rect 20244 23884 20254 23940
rect 20738 23884 20748 23940
rect 20804 23884 22540 23940
rect 22596 23884 22606 23940
rect 20514 23772 20524 23828
rect 20580 23772 21980 23828
rect 22036 23772 22046 23828
rect 22866 23772 22876 23828
rect 22932 23772 23772 23828
rect 23828 23772 23838 23828
rect 14802 23660 14812 23716
rect 14868 23660 15596 23716
rect 15652 23660 18676 23716
rect 18834 23660 18844 23716
rect 18900 23660 19628 23716
rect 19684 23660 21420 23716
rect 21476 23660 26236 23716
rect 26292 23660 26302 23716
rect 18620 23604 18676 23660
rect 14914 23548 14924 23604
rect 14980 23548 17948 23604
rect 18004 23548 18172 23604
rect 18228 23548 18238 23604
rect 18610 23548 18620 23604
rect 18676 23548 18956 23604
rect 19012 23548 19022 23604
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 14466 23436 14476 23492
rect 14532 23436 19404 23492
rect 19460 23436 19470 23492
rect 16818 23324 16828 23380
rect 16884 23324 17500 23380
rect 17556 23324 19068 23380
rect 19124 23324 19134 23380
rect 19282 23212 19292 23268
rect 19348 23212 20188 23268
rect 20244 23212 20254 23268
rect 4274 23100 4284 23156
rect 4340 23100 13916 23156
rect 13972 23100 16940 23156
rect 16996 23100 17006 23156
rect 22754 23100 22764 23156
rect 22820 23100 23996 23156
rect 24052 23100 24062 23156
rect 24546 22988 24556 23044
rect 24612 22988 25788 23044
rect 25844 22988 25854 23044
rect 0 22932 800 22960
rect 0 22876 1932 22932
rect 1988 22876 1998 22932
rect 0 22848 800 22876
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 18722 22652 18732 22708
rect 18788 22652 20860 22708
rect 20916 22652 20926 22708
rect 1922 22428 1932 22484
rect 1988 22428 1998 22484
rect 0 22260 800 22288
rect 1932 22260 1988 22428
rect 4274 22316 4284 22372
rect 4340 22316 8428 22372
rect 13682 22316 13692 22372
rect 13748 22316 19292 22372
rect 19348 22316 19358 22372
rect 23650 22316 23660 22372
rect 23716 22316 25452 22372
rect 25508 22316 26460 22372
rect 26516 22316 26526 22372
rect 0 22204 1988 22260
rect 8372 22260 8428 22316
rect 41200 22260 42000 22288
rect 8372 22204 9996 22260
rect 10052 22204 13580 22260
rect 13636 22204 13646 22260
rect 15026 22204 15036 22260
rect 15092 22204 16044 22260
rect 16100 22204 16110 22260
rect 16594 22204 16604 22260
rect 16660 22204 17276 22260
rect 17332 22204 17342 22260
rect 40002 22204 40012 22260
rect 40068 22204 42000 22260
rect 0 22176 800 22204
rect 16044 22148 16100 22204
rect 41200 22176 42000 22204
rect 12898 22092 12908 22148
rect 12964 22092 14140 22148
rect 14196 22092 14206 22148
rect 16044 22092 18284 22148
rect 18340 22092 19180 22148
rect 19236 22092 19246 22148
rect 21858 21980 21868 22036
rect 21924 21980 25228 22036
rect 25284 21980 26348 22036
rect 26404 21980 26414 22036
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 23874 21868 23884 21924
rect 23940 21868 24780 21924
rect 24836 21868 37660 21924
rect 37716 21868 37726 21924
rect 12114 21756 12124 21812
rect 12180 21756 13132 21812
rect 13188 21756 13198 21812
rect 22754 21756 22764 21812
rect 22820 21756 24332 21812
rect 24388 21756 24398 21812
rect 21298 21644 21308 21700
rect 21364 21644 23436 21700
rect 23492 21644 27356 21700
rect 27412 21644 27422 21700
rect 41200 21588 42000 21616
rect 17602 21532 17612 21588
rect 17668 21532 18172 21588
rect 18228 21532 20412 21588
rect 20468 21532 20636 21588
rect 20692 21532 20702 21588
rect 20962 21532 20972 21588
rect 21028 21532 21868 21588
rect 21924 21532 21934 21588
rect 24434 21532 24444 21588
rect 24500 21532 25900 21588
rect 25956 21532 25966 21588
rect 40002 21532 40012 21588
rect 40068 21532 42000 21588
rect 41200 21504 42000 21532
rect 22530 21420 22540 21476
rect 22596 21420 23548 21476
rect 23604 21420 23614 21476
rect 22978 21308 22988 21364
rect 23044 21308 25564 21364
rect 25620 21308 25630 21364
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 25890 20972 25900 21028
rect 25956 20972 26684 21028
rect 26740 20972 26750 21028
rect 41200 20916 42000 20944
rect 25218 20860 25228 20916
rect 25284 20860 25676 20916
rect 25732 20860 25742 20916
rect 40002 20860 40012 20916
rect 40068 20860 42000 20916
rect 41200 20832 42000 20860
rect 20738 20748 20748 20804
rect 20804 20748 21868 20804
rect 21924 20748 22652 20804
rect 22708 20748 22718 20804
rect 26562 20748 26572 20804
rect 26628 20748 28588 20804
rect 28644 20748 28654 20804
rect 29362 20748 29372 20804
rect 29428 20748 29932 20804
rect 29988 20748 29998 20804
rect 31892 20748 37660 20804
rect 37716 20748 37726 20804
rect 13906 20636 13916 20692
rect 13972 20636 21308 20692
rect 21364 20636 21374 20692
rect 26338 20636 26348 20692
rect 26404 20636 27692 20692
rect 27748 20636 27758 20692
rect 31892 20580 31948 20748
rect 11442 20524 11452 20580
rect 11508 20524 13468 20580
rect 13524 20524 13534 20580
rect 29586 20524 29596 20580
rect 29652 20524 29662 20580
rect 30258 20524 30268 20580
rect 30324 20524 31948 20580
rect 29596 20468 29652 20524
rect 29596 20412 37884 20468
rect 37940 20412 37950 20468
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 41200 20244 42000 20272
rect 13682 20188 13692 20244
rect 13748 20188 14252 20244
rect 14308 20188 14318 20244
rect 21970 20188 21980 20244
rect 22036 20188 22988 20244
rect 23044 20188 23054 20244
rect 40012 20188 42000 20244
rect 40012 20132 40068 20188
rect 41200 20160 42000 20188
rect 4162 20076 4172 20132
rect 4228 20076 18956 20132
rect 19012 20076 19292 20132
rect 19348 20076 19358 20132
rect 20132 20076 22092 20132
rect 22148 20076 22158 20132
rect 26898 20076 26908 20132
rect 26964 20076 29932 20132
rect 29988 20076 29998 20132
rect 40002 20076 40012 20132
rect 40068 20076 40078 20132
rect 20132 20020 20188 20076
rect 13458 19964 13468 20020
rect 13524 19964 15148 20020
rect 15204 19964 15214 20020
rect 16370 19964 16380 20020
rect 16436 19964 17388 20020
rect 17444 19964 20188 20020
rect 10098 19852 10108 19908
rect 10164 19852 10780 19908
rect 10836 19852 13916 19908
rect 13972 19852 13982 19908
rect 14578 19852 14588 19908
rect 14644 19852 15036 19908
rect 15092 19852 15932 19908
rect 15988 19852 15998 19908
rect 16828 19852 17612 19908
rect 17668 19852 18228 19908
rect 20178 19852 20188 19908
rect 20244 19852 20636 19908
rect 20692 19852 20702 19908
rect 27458 19852 27468 19908
rect 27524 19852 28588 19908
rect 28644 19852 31948 19908
rect 16828 19796 16884 19852
rect 18172 19796 18228 19852
rect 31892 19796 31948 19852
rect 13234 19740 13244 19796
rect 13300 19740 16884 19796
rect 17042 19740 17052 19796
rect 17108 19740 17948 19796
rect 18004 19740 18014 19796
rect 18172 19740 21532 19796
rect 21588 19740 21598 19796
rect 31892 19740 37660 19796
rect 37716 19740 37726 19796
rect 14690 19628 14700 19684
rect 14756 19628 16492 19684
rect 16548 19628 17724 19684
rect 17780 19628 21420 19684
rect 21476 19628 22652 19684
rect 22708 19628 22718 19684
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 41200 19572 42000 19600
rect 40002 19516 40012 19572
rect 40068 19516 42000 19572
rect 41200 19488 42000 19516
rect 15250 19404 15260 19460
rect 15316 19404 16268 19460
rect 16324 19404 17388 19460
rect 17444 19404 17454 19460
rect 19282 19404 19292 19460
rect 19348 19404 20748 19460
rect 20804 19404 20814 19460
rect 12898 19292 12908 19348
rect 12964 19292 13804 19348
rect 13860 19292 14476 19348
rect 14532 19292 16044 19348
rect 16100 19292 16110 19348
rect 19618 19292 19628 19348
rect 19684 19292 25452 19348
rect 25508 19292 25518 19348
rect 18060 19180 20188 19236
rect 20244 19180 21196 19236
rect 21252 19180 21262 19236
rect 14018 19068 14028 19124
rect 14084 19068 15036 19124
rect 15092 19068 16044 19124
rect 16100 19068 16110 19124
rect 18060 19012 18116 19180
rect 25452 19124 25508 19292
rect 18946 19068 18956 19124
rect 19012 19068 23996 19124
rect 24052 19068 24062 19124
rect 25452 19068 25900 19124
rect 25956 19068 25966 19124
rect 29922 19068 29932 19124
rect 29988 19068 37884 19124
rect 37940 19068 37950 19124
rect 16594 18956 16604 19012
rect 16660 18956 17724 19012
rect 17780 18956 18116 19012
rect 18956 18900 19012 19068
rect 25218 18956 25228 19012
rect 25284 18956 25676 19012
rect 25732 18956 25742 19012
rect 15586 18844 15596 18900
rect 15652 18844 19012 18900
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 14578 18732 14588 18788
rect 14644 18732 17500 18788
rect 17556 18732 17566 18788
rect 15474 18620 15484 18676
rect 15540 18620 17164 18676
rect 17220 18620 17230 18676
rect 13122 18508 13132 18564
rect 13188 18508 13916 18564
rect 13972 18508 13982 18564
rect 20374 18508 20412 18564
rect 20468 18508 20478 18564
rect 16370 18396 16380 18452
rect 16436 18396 17052 18452
rect 17108 18396 18172 18452
rect 18228 18396 18620 18452
rect 18676 18396 18686 18452
rect 18834 18396 18844 18452
rect 18900 18396 19292 18452
rect 19348 18396 19740 18452
rect 19796 18396 21756 18452
rect 21812 18396 21822 18452
rect 21970 18396 21980 18452
rect 22036 18396 22540 18452
rect 22596 18396 23324 18452
rect 23380 18396 23390 18452
rect 23762 18396 23772 18452
rect 23828 18396 25228 18452
rect 25284 18396 25294 18452
rect 10770 18284 10780 18340
rect 10836 18284 14924 18340
rect 14980 18284 20300 18340
rect 20356 18284 21308 18340
rect 21364 18284 21374 18340
rect 23538 18284 23548 18340
rect 23604 18284 24668 18340
rect 24724 18284 24734 18340
rect 15362 18172 15372 18228
rect 15428 18172 16156 18228
rect 16212 18172 16222 18228
rect 16818 18172 16828 18228
rect 16884 18172 17836 18228
rect 17892 18172 17902 18228
rect 19842 18172 19852 18228
rect 19908 18172 20412 18228
rect 20468 18172 20478 18228
rect 20738 18172 20748 18228
rect 20804 18172 22428 18228
rect 22484 18172 22494 18228
rect 24098 18172 24108 18228
rect 24164 18172 25452 18228
rect 25508 18172 25518 18228
rect 16156 18116 16212 18172
rect 20300 18116 20356 18172
rect 16156 18060 17276 18116
rect 17332 18060 17342 18116
rect 17612 18060 19180 18116
rect 19236 18060 19246 18116
rect 20300 18060 21868 18116
rect 21924 18060 21934 18116
rect 23426 18060 23436 18116
rect 23492 18060 25956 18116
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 17612 18004 17668 18060
rect 25900 18004 25956 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 15698 17948 15708 18004
rect 15764 17948 17612 18004
rect 17668 17948 17678 18004
rect 17826 17948 17836 18004
rect 17892 17948 23772 18004
rect 23828 17948 23838 18004
rect 25890 17948 25900 18004
rect 25956 17948 26572 18004
rect 26628 17948 26638 18004
rect 17154 17836 17164 17892
rect 17220 17836 18732 17892
rect 18788 17836 18798 17892
rect 19170 17836 19180 17892
rect 19236 17836 19964 17892
rect 20020 17836 20030 17892
rect 20178 17836 20188 17892
rect 20244 17836 20524 17892
rect 20580 17836 20590 17892
rect 1922 17724 1932 17780
rect 1988 17724 1998 17780
rect 17042 17724 17052 17780
rect 17108 17724 18956 17780
rect 19012 17724 19022 17780
rect 19170 17724 19180 17780
rect 19236 17724 20748 17780
rect 20804 17724 20814 17780
rect 0 17556 800 17584
rect 1932 17556 1988 17724
rect 4274 17612 4284 17668
rect 4340 17612 13468 17668
rect 13524 17612 16604 17668
rect 16660 17612 16670 17668
rect 16828 17612 21700 17668
rect 21858 17612 21868 17668
rect 21924 17612 23436 17668
rect 23492 17612 23502 17668
rect 24210 17612 24220 17668
rect 24276 17612 25004 17668
rect 25060 17612 26908 17668
rect 26964 17612 26974 17668
rect 16828 17556 16884 17612
rect 21644 17556 21700 17612
rect 0 17500 1988 17556
rect 16034 17500 16044 17556
rect 16100 17500 16884 17556
rect 19954 17500 19964 17556
rect 20020 17500 20244 17556
rect 21644 17500 22204 17556
rect 22260 17500 23548 17556
rect 23604 17500 23614 17556
rect 25666 17500 25676 17556
rect 25732 17500 27244 17556
rect 27300 17500 27310 17556
rect 0 17472 800 17500
rect 18834 17388 18844 17444
rect 18900 17388 19516 17444
rect 19572 17388 19582 17444
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 20188 17108 20244 17500
rect 21634 17388 21644 17444
rect 21700 17388 22092 17444
rect 22148 17388 25228 17444
rect 25284 17388 25294 17444
rect 26562 17388 26572 17444
rect 26628 17388 27356 17444
rect 27412 17388 27422 17444
rect 27010 17276 27020 17332
rect 27076 17276 27468 17332
rect 27524 17276 37660 17332
rect 37716 17276 37726 17332
rect 20738 17164 20748 17220
rect 20804 17164 21420 17220
rect 21476 17164 22204 17220
rect 22260 17164 22270 17220
rect 24770 17164 24780 17220
rect 24836 17164 24846 17220
rect 24780 17108 24836 17164
rect 14130 17052 14140 17108
rect 14196 17052 15260 17108
rect 15316 17052 15326 17108
rect 19954 17052 19964 17108
rect 20020 17052 24836 17108
rect 15586 16940 15596 16996
rect 15652 16940 17724 16996
rect 17780 16940 22764 16996
rect 22820 16940 22830 16996
rect 4274 16828 4284 16884
rect 4340 16828 12012 16884
rect 12068 16828 12078 16884
rect 15698 16828 15708 16884
rect 15764 16828 17500 16884
rect 17556 16828 17566 16884
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 16594 16268 16604 16324
rect 16660 16268 17948 16324
rect 18004 16268 18014 16324
rect 0 16212 800 16240
rect 41200 16212 42000 16240
rect 0 16156 1932 16212
rect 1988 16156 1998 16212
rect 40002 16156 40012 16212
rect 40068 16156 42000 16212
rect 0 16128 800 16156
rect 41200 16128 42000 16156
rect 20738 16044 20748 16100
rect 20804 16044 22316 16100
rect 22372 16044 22382 16100
rect 24546 16044 24556 16100
rect 24612 16044 25228 16100
rect 25284 16044 27916 16100
rect 27972 16044 27982 16100
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 12002 15372 12012 15428
rect 12068 15372 15260 15428
rect 15316 15372 15326 15428
rect 19618 15260 19628 15316
rect 19684 15260 20188 15316
rect 20244 15260 22988 15316
rect 23044 15260 23548 15316
rect 23604 15260 24556 15316
rect 24612 15260 24622 15316
rect 13122 15148 13132 15204
rect 13188 15148 14924 15204
rect 14980 15148 15932 15204
rect 15988 15148 16268 15204
rect 16324 15148 16828 15204
rect 16884 15148 19180 15204
rect 19236 15148 19246 15204
rect 21970 15148 21980 15204
rect 22036 15148 23100 15204
rect 23156 15148 24444 15204
rect 24500 15148 24510 15204
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 22530 13468 22540 13524
rect 22596 13468 23548 13524
rect 23604 13468 23614 13524
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 41200 10164 42000 10192
rect 40226 10108 40236 10164
rect 40292 10108 42000 10164
rect 41200 10080 42000 10108
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 22866 3612 22876 3668
rect 22932 3612 25564 3668
rect 25620 3612 25630 3668
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
<< via3 >>
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 20412 18508 20468 18564
rect 20412 18172 20468 18228
rect 19180 18060 19236 18116
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 19180 17724 19236 17780
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
<< metal4 >>
rect 4448 38444 4768 38476
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 19808 37660 20128 38476
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19808 34524 20128 36036
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 19808 23548 20128 25060
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 19808 21980 20128 23492
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 19180 18116 19236 18126
rect 19180 17780 19236 18060
rect 19180 17714 19236 17724
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 17276 20128 18788
rect 35168 38444 35488 38476
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 20412 18564 20468 18574
rect 20412 18228 20468 18508
rect 20412 18162 20468 18172
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _087_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 24528 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _088_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 26768 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _089_
timestamp 1698175906
transform 1 0 13552 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _090_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 15232 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _091_
timestamp 1698175906
transform 1 0 14224 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _092_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 20272 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _093_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21168 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _094_
timestamp 1698175906
transform 1 0 19376 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _095_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 23184 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _096_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 25200 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _097_
timestamp 1698175906
transform 1 0 14224 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _098_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 14896 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _099_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 14896 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _100_
timestamp 1698175906
transform 1 0 14896 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _101_
timestamp 1698175906
transform -1 0 14000 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _102_
timestamp 1698175906
transform -1 0 18704 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _103_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 15904 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _104_
timestamp 1698175906
transform 1 0 19824 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _105_
timestamp 1698175906
transform -1 0 20944 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _106_
timestamp 1698175906
transform 1 0 17920 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _107_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 17248 0 1 18816
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _108_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17248 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _109_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 24528 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _110_
timestamp 1698175906
transform 1 0 23856 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _111_
timestamp 1698175906
transform 1 0 25088 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _112_
timestamp 1698175906
transform 1 0 26096 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _113_
timestamp 1698175906
transform 1 0 18816 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _114_
timestamp 1698175906
transform -1 0 19376 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _115_
timestamp 1698175906
transform 1 0 18480 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _116_
timestamp 1698175906
transform -1 0 19264 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _117_
timestamp 1698175906
transform 1 0 20272 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _118_
timestamp 1698175906
transform 1 0 22064 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _119_
timestamp 1698175906
transform -1 0 20944 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _120_
timestamp 1698175906
transform 1 0 17248 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _121_
timestamp 1698175906
transform -1 0 20608 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _122_
timestamp 1698175906
transform 1 0 26320 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _123_
timestamp 1698175906
transform 1 0 18368 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _124_
timestamp 1698175906
transform 1 0 27776 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _125_
timestamp 1698175906
transform 1 0 25984 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _126_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 22064 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _127_
timestamp 1698175906
transform 1 0 21616 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _128_
timestamp 1698175906
transform -1 0 22064 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _129_
timestamp 1698175906
transform -1 0 16128 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _130_
timestamp 1698175906
transform -1 0 18592 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _131_
timestamp 1698175906
transform 1 0 18816 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _132_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 14112 0 -1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _133_
timestamp 1698175906
transform 1 0 12656 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _134_
timestamp 1698175906
transform 1 0 14224 0 1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _135_
timestamp 1698175906
transform 1 0 13328 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _136_
timestamp 1698175906
transform 1 0 18704 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _137_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 20160 0 1 25088
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _138_
timestamp 1698175906
transform -1 0 26656 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _139_
timestamp 1698175906
transform 1 0 22288 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _140_
timestamp 1698175906
transform 1 0 24080 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _141_
timestamp 1698175906
transform 1 0 25312 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _142_
timestamp 1698175906
transform -1 0 22736 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _143_
timestamp 1698175906
transform 1 0 24528 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _144_
timestamp 1698175906
transform -1 0 21840 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _145_
timestamp 1698175906
transform 1 0 27216 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _146_
timestamp 1698175906
transform 1 0 25536 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _147_
timestamp 1698175906
transform -1 0 18144 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _148_
timestamp 1698175906
transform -1 0 13888 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _149_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 14224 0 -1 21952
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _150_
timestamp 1698175906
transform 1 0 15904 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _151_
timestamp 1698175906
transform 1 0 22288 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _152_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21168 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _153_
timestamp 1698175906
transform 1 0 21952 0 -1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _154_
timestamp 1698175906
transform -1 0 22400 0 1 23520
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _155_
timestamp 1698175906
transform 1 0 25424 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _156_
timestamp 1698175906
transform -1 0 27552 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _157_
timestamp 1698175906
transform 1 0 28112 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _158_
timestamp 1698175906
transform 1 0 16576 0 1 17248
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _159_
timestamp 1698175906
transform 1 0 17248 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _160_
timestamp 1698175906
transform 1 0 20048 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _161_
timestamp 1698175906
transform 1 0 23296 0 1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _162_
timestamp 1698175906
transform -1 0 23072 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _163_
timestamp 1698175906
transform 1 0 20496 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _164_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 23296 0 -1 21952
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _165_
timestamp 1698175906
transform 1 0 21728 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _166_
timestamp 1698175906
transform 1 0 15120 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _167_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 16240 0 -1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _168_
timestamp 1698175906
transform 1 0 15232 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _169_
timestamp 1698175906
transform 1 0 18256 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _170_
timestamp 1698175906
transform -1 0 18816 0 -1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _171_
timestamp 1698175906
transform -1 0 17808 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _172_
timestamp 1698175906
transform 1 0 16800 0 1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _173_
timestamp 1698175906
transform 1 0 15904 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _174_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 24416 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _175_
timestamp 1698175906
transform 1 0 9856 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _176_
timestamp 1698175906
transform 1 0 10528 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _177_
timestamp 1698175906
transform 1 0 15680 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _178_
timestamp 1698175906
transform -1 0 28336 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _179_
timestamp 1698175906
transform 1 0 19488 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _180_
timestamp 1698175906
transform 1 0 25536 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _181_
timestamp 1698175906
transform 1 0 20048 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _182_
timestamp 1698175906
transform -1 0 14112 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _183_
timestamp 1698175906
transform -1 0 14896 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _184_
timestamp 1698175906
transform -1 0 20384 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _185_
timestamp 1698175906
transform 1 0 24976 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _186_
timestamp 1698175906
transform 1 0 25536 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _187_
timestamp 1698175906
transform -1 0 13104 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _188_
timestamp 1698175906
transform 1 0 20272 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _189_
timestamp 1698175906
transform -1 0 29792 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _190_
timestamp 1698175906
transform -1 0 16576 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _191_
timestamp 1698175906
transform 1 0 21728 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _192_
timestamp 1698175906
transform 1 0 21728 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _193_
timestamp 1698175906
transform -1 0 15120 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _194_
timestamp 1698175906
transform 1 0 15680 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _195_
timestamp 1698175906
transform -1 0 17024 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _198_
timestamp 1698175906
transform -1 0 14672 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _199_
timestamp 1698175906
transform 1 0 29120 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _200_
timestamp 1698175906
transform 1 0 19376 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _201_
timestamp 1698175906
transform 1 0 29792 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _202_
timestamp 1698175906
transform 1 0 27104 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _203_
timestamp 1698175906
transform -1 0 15568 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__174__CLK dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 27888 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__175__CLK
timestamp 1698175906
transform 1 0 13104 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__176__CLK
timestamp 1698175906
transform 1 0 14000 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__177__CLK
timestamp 1698175906
transform 1 0 19152 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__178__CLK
timestamp 1698175906
transform 1 0 28560 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__179__CLK
timestamp 1698175906
transform 1 0 22960 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__180__CLK
timestamp 1698175906
transform 1 0 29232 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__181__CLK
timestamp 1698175906
transform 1 0 23520 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__182__CLK
timestamp 1698175906
transform 1 0 14112 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__183__CLK
timestamp 1698175906
transform -1 0 16016 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__184__CLK
timestamp 1698175906
transform 1 0 20608 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__185__CLK
timestamp 1698175906
transform 1 0 28448 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__186__CLK
timestamp 1698175906
transform 1 0 29008 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__187__CLK
timestamp 1698175906
transform 1 0 14112 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__188__CLK
timestamp 1698175906
transform 1 0 23744 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__189__CLK
timestamp 1698175906
transform 1 0 26320 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__190__CLK
timestamp 1698175906
transform 1 0 16800 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__191__CLK
timestamp 1698175906
transform 1 0 25312 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__192__CLK
timestamp 1698175906
transform 1 0 25200 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__193__CLK
timestamp 1698175906
transform 1 0 15792 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__194__CLK
timestamp 1698175906
transform 1 0 19040 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__195__CLK
timestamp 1698175906
transform 1 0 17472 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1698175906
transform 1 0 18928 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19152 0 -1 20384
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1698175906
transform -1 0 20944 0 1 20384
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1698175906
transform 1 0 22512 0 1 20384
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1568 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698175906
transform 1 0 5376 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698175906
transform 1 0 9184 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698175906
transform 1 0 12992 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_138
timestamp 1698175906
transform 1 0 16800 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_172 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 20608 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_176 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21056 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_232
timestamp 1698175906
transform 1 0 27328 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_236
timestamp 1698175906
transform 1 0 27776 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_240
timestamp 1698175906
transform 1 0 28224 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_274
timestamp 1698175906
transform 1 0 32032 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_308
timestamp 1698175906
transform 1 0 35840 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_342
timestamp 1698175906
transform 1 0 39648 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_346
timestamp 1698175906
transform 1 0 40096 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_348 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 40320 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1568 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698175906
transform 1 0 8736 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698175906
transform 1 0 9408 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698175906
transform 1 0 16576 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_142
timestamp 1698175906
transform 1 0 17248 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_206
timestamp 1698175906
transform 1 0 24416 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_212
timestamp 1698175906
transform 1 0 25088 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_276
timestamp 1698175906
transform 1 0 32256 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_282
timestamp 1698175906
transform 1 0 32928 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_346
timestamp 1698175906
transform 1 0 40096 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_348
timestamp 1698175906
transform 1 0 40320 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698175906
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698175906
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698175906
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698175906
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_107
timestamp 1698175906
transform 1 0 13328 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_171
timestamp 1698175906
transform 1 0 20496 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_177
timestamp 1698175906
transform 1 0 21168 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_241
timestamp 1698175906
transform 1 0 28336 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698175906
transform 1 0 29008 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698175906
transform 1 0 36176 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_317
timestamp 1698175906
transform 1 0 36848 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698175906
transform 1 0 1568 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698175906
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698175906
transform 1 0 9408 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698175906
transform 1 0 16576 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_142
timestamp 1698175906
transform 1 0 17248 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_206
timestamp 1698175906
transform 1 0 24416 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_212
timestamp 1698175906
transform 1 0 25088 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_276
timestamp 1698175906
transform 1 0 32256 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_282
timestamp 1698175906
transform 1 0 32928 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_346
timestamp 1698175906
transform 1 0 40096 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_348
timestamp 1698175906
transform 1 0 40320 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698175906
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698175906
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698175906
transform 1 0 5488 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698175906
transform 1 0 12656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_107
timestamp 1698175906
transform 1 0 13328 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698175906
transform 1 0 20496 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_177
timestamp 1698175906
transform 1 0 21168 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_241
timestamp 1698175906
transform 1 0 28336 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698175906
transform 1 0 29008 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698175906
transform 1 0 36176 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_317
timestamp 1698175906
transform 1 0 36848 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698175906
transform 1 0 1568 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698175906
transform 1 0 8736 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698175906
transform 1 0 9408 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698175906
transform 1 0 16576 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_142
timestamp 1698175906
transform 1 0 17248 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_206
timestamp 1698175906
transform 1 0 24416 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_212
timestamp 1698175906
transform 1 0 25088 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698175906
transform 1 0 32256 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_282
timestamp 1698175906
transform 1 0 32928 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_346
timestamp 1698175906
transform 1 0 40096 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_348
timestamp 1698175906
transform 1 0 40320 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698175906
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698175906
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698175906
transform 1 0 5488 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698175906
transform 1 0 12656 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_107
timestamp 1698175906
transform 1 0 13328 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_171
timestamp 1698175906
transform 1 0 20496 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_177
timestamp 1698175906
transform 1 0 21168 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_241
timestamp 1698175906
transform 1 0 28336 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_247
timestamp 1698175906
transform 1 0 29008 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_311
timestamp 1698175906
transform 1 0 36176 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_317
timestamp 1698175906
transform 1 0 36848 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698175906
transform 1 0 1568 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698175906
transform 1 0 8736 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_72
timestamp 1698175906
transform 1 0 9408 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698175906
transform 1 0 16576 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_142
timestamp 1698175906
transform 1 0 17248 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_206
timestamp 1698175906
transform 1 0 24416 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_212
timestamp 1698175906
transform 1 0 25088 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_276
timestamp 1698175906
transform 1 0 32256 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_282
timestamp 1698175906
transform 1 0 32928 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_346
timestamp 1698175906
transform 1 0 40096 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_348
timestamp 1698175906
transform 1 0 40320 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698175906
transform 1 0 1568 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698175906
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_37
timestamp 1698175906
transform 1 0 5488 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_101
timestamp 1698175906
transform 1 0 12656 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_107
timestamp 1698175906
transform 1 0 13328 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_171
timestamp 1698175906
transform 1 0 20496 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_177
timestamp 1698175906
transform 1 0 21168 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_241
timestamp 1698175906
transform 1 0 28336 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_247
timestamp 1698175906
transform 1 0 29008 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_311
timestamp 1698175906
transform 1 0 36176 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_317
timestamp 1698175906
transform 1 0 36848 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698175906
transform 1 0 1568 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698175906
transform 1 0 8736 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_72
timestamp 1698175906
transform 1 0 9408 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_136
timestamp 1698175906
transform 1 0 16576 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_142
timestamp 1698175906
transform 1 0 17248 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_206
timestamp 1698175906
transform 1 0 24416 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_212
timestamp 1698175906
transform 1 0 25088 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_276
timestamp 1698175906
transform 1 0 32256 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_9_282
timestamp 1698175906
transform 1 0 32928 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_314 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 36512 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_330 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 38304 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_338
timestamp 1698175906
transform 1 0 39200 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_342
timestamp 1698175906
transform 1 0 39648 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_344
timestamp 1698175906
transform 1 0 39872 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698175906
transform 1 0 1568 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698175906
transform 1 0 5152 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_37
timestamp 1698175906
transform 1 0 5488 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698175906
transform 1 0 12656 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_107
timestamp 1698175906
transform 1 0 13328 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_171
timestamp 1698175906
transform 1 0 20496 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_177
timestamp 1698175906
transform 1 0 21168 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_241
timestamp 1698175906
transform 1 0 28336 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_247
timestamp 1698175906
transform 1 0 29008 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_311
timestamp 1698175906
transform 1 0 36176 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_317
timestamp 1698175906
transform 1 0 36848 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2
timestamp 1698175906
transform 1 0 1568 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698175906
transform 1 0 8736 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_72
timestamp 1698175906
transform 1 0 9408 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698175906
transform 1 0 16576 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_142
timestamp 1698175906
transform 1 0 17248 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_206
timestamp 1698175906
transform 1 0 24416 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_212
timestamp 1698175906
transform 1 0 25088 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_276
timestamp 1698175906
transform 1 0 32256 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_282
timestamp 1698175906
transform 1 0 32928 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_346
timestamp 1698175906
transform 1 0 40096 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_348
timestamp 1698175906
transform 1 0 40320 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698175906
transform 1 0 1568 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698175906
transform 1 0 5152 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_37
timestamp 1698175906
transform 1 0 5488 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698175906
transform 1 0 12656 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_107
timestamp 1698175906
transform 1 0 13328 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_171
timestamp 1698175906
transform 1 0 20496 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_177
timestamp 1698175906
transform 1 0 21168 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_241
timestamp 1698175906
transform 1 0 28336 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_247
timestamp 1698175906
transform 1 0 29008 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_311
timestamp 1698175906
transform 1 0 36176 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_317
timestamp 1698175906
transform 1 0 36848 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_2
timestamp 1698175906
transform 1 0 1568 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_66
timestamp 1698175906
transform 1 0 8736 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_72
timestamp 1698175906
transform 1 0 9408 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_136
timestamp 1698175906
transform 1 0 16576 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_142
timestamp 1698175906
transform 1 0 17248 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_158
timestamp 1698175906
transform 1 0 19040 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_191
timestamp 1698175906
transform 1 0 22736 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_195
timestamp 1698175906
transform 1 0 23184 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_203
timestamp 1698175906
transform 1 0 24080 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_207
timestamp 1698175906
transform 1 0 24528 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_209
timestamp 1698175906
transform 1 0 24752 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_212
timestamp 1698175906
transform 1 0 25088 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_276
timestamp 1698175906
transform 1 0 32256 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_282
timestamp 1698175906
transform 1 0 32928 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_346
timestamp 1698175906
transform 1 0 40096 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_348
timestamp 1698175906
transform 1 0 40320 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698175906
transform 1 0 1568 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698175906
transform 1 0 5152 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_37
timestamp 1698175906
transform 1 0 5488 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_101
timestamp 1698175906
transform 1 0 12656 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_107
timestamp 1698175906
transform 1 0 13328 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_123
timestamp 1698175906
transform 1 0 15120 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_127
timestamp 1698175906
transform 1 0 15568 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_157
timestamp 1698175906
transform 1 0 18928 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_161
timestamp 1698175906
transform 1 0 19376 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_169
timestamp 1698175906
transform 1 0 20272 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_173
timestamp 1698175906
transform 1 0 20720 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_177
timestamp 1698175906
transform 1 0 21168 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_241
timestamp 1698175906
transform 1 0 28336 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_247
timestamp 1698175906
transform 1 0 29008 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_311
timestamp 1698175906
transform 1 0 36176 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_317
timestamp 1698175906
transform 1 0 36848 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_2
timestamp 1698175906
transform 1 0 1568 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_66
timestamp 1698175906
transform 1 0 8736 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_72
timestamp 1698175906
transform 1 0 9408 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_88
timestamp 1698175906
transform 1 0 11200 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_92
timestamp 1698175906
transform 1 0 11648 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_127
timestamp 1698175906
transform 1 0 15568 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_131
timestamp 1698175906
transform 1 0 16016 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_139
timestamp 1698175906
transform 1 0 16912 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_142
timestamp 1698175906
transform 1 0 17248 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_158
timestamp 1698175906
transform 1 0 19040 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_166
timestamp 1698175906
transform 1 0 19936 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_196
timestamp 1698175906
transform 1 0 23296 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_200
timestamp 1698175906
transform 1 0 23744 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_208
timestamp 1698175906
transform 1 0 24640 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_212
timestamp 1698175906
transform 1 0 25088 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_276
timestamp 1698175906
transform 1 0 32256 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_282
timestamp 1698175906
transform 1 0 32928 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_346
timestamp 1698175906
transform 1 0 40096 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_348
timestamp 1698175906
transform 1 0 40320 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_2
timestamp 1698175906
transform 1 0 1568 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698175906
transform 1 0 5152 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_37
timestamp 1698175906
transform 1 0 5488 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_101
timestamp 1698175906
transform 1 0 12656 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_136
timestamp 1698175906
transform 1 0 16576 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_140
timestamp 1698175906
transform 1 0 17024 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_156
timestamp 1698175906
transform 1 0 18816 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_164
timestamp 1698175906
transform 1 0 19712 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_166
timestamp 1698175906
transform 1 0 19936 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_191
timestamp 1698175906
transform 1 0 22736 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_199
timestamp 1698175906
transform 1 0 23632 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_203
timestamp 1698175906
transform 1 0 24080 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_205
timestamp 1698175906
transform 1 0 24304 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_235
timestamp 1698175906
transform 1 0 27664 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_239
timestamp 1698175906
transform 1 0 28112 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_243
timestamp 1698175906
transform 1 0 28560 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_247
timestamp 1698175906
transform 1 0 29008 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_311
timestamp 1698175906
transform 1 0 36176 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_317
timestamp 1698175906
transform 1 0 36848 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_28
timestamp 1698175906
transform 1 0 4480 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_60
timestamp 1698175906
transform 1 0 8064 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_68
timestamp 1698175906
transform 1 0 8960 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_72
timestamp 1698175906
transform 1 0 9408 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_104
timestamp 1698175906
transform 1 0 12992 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_120
timestamp 1698175906
transform 1 0 14784 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_122
timestamp 1698175906
transform 1 0 15008 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_133
timestamp 1698175906
transform 1 0 16240 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_137
timestamp 1698175906
transform 1 0 16688 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_139
timestamp 1698175906
transform 1 0 16912 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_150
timestamp 1698175906
transform 1 0 18144 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_158
timestamp 1698175906
transform 1 0 19040 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_162
timestamp 1698175906
transform 1 0 19488 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_164
timestamp 1698175906
transform 1 0 19712 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_169
timestamp 1698175906
transform 1 0 20272 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_177
timestamp 1698175906
transform 1 0 21168 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_186
timestamp 1698175906
transform 1 0 22176 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_202
timestamp 1698175906
transform 1 0 23968 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_241
timestamp 1698175906
transform 1 0 28336 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_245
timestamp 1698175906
transform 1 0 28784 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_277
timestamp 1698175906
transform 1 0 32368 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_279
timestamp 1698175906
transform 1 0 32592 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_282
timestamp 1698175906
transform 1 0 32928 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_314
timestamp 1698175906
transform 1 0 36512 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_322
timestamp 1698175906
transform 1 0 37408 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_28
timestamp 1698175906
transform 1 0 4480 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_32
timestamp 1698175906
transform 1 0 4928 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698175906
transform 1 0 5152 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_37
timestamp 1698175906
transform 1 0 5488 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_101
timestamp 1698175906
transform 1 0 12656 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_107
timestamp 1698175906
transform 1 0 13328 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_123
timestamp 1698175906
transform 1 0 15120 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_131
timestamp 1698175906
transform 1 0 16016 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_135
timestamp 1698175906
transform 1 0 16464 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_147
timestamp 1698175906
transform 1 0 17808 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_167
timestamp 1698175906
transform 1 0 20048 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_191
timestamp 1698175906
transform 1 0 22736 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_232
timestamp 1698175906
transform 1 0 27328 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_240
timestamp 1698175906
transform 1 0 28224 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_244
timestamp 1698175906
transform 1 0 28672 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_247
timestamp 1698175906
transform 1 0 29008 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_311
timestamp 1698175906
transform 1 0 36176 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_317
timestamp 1698175906
transform 1 0 36848 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_2
timestamp 1698175906
transform 1 0 1568 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_66
timestamp 1698175906
transform 1 0 8736 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_72
timestamp 1698175906
transform 1 0 9408 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_104
timestamp 1698175906
transform 1 0 12992 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_107
timestamp 1698175906
transform 1 0 13328 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_115
timestamp 1698175906
transform 1 0 14224 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_119
timestamp 1698175906
transform 1 0 14672 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_150
timestamp 1698175906
transform 1 0 18144 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_152
timestamp 1698175906
transform 1 0 18368 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_161
timestamp 1698175906
transform 1 0 19376 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_175
timestamp 1698175906
transform 1 0 20944 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_193
timestamp 1698175906
transform 1 0 22960 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_206
timestamp 1698175906
transform 1 0 24416 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_220
timestamp 1698175906
transform 1 0 25984 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_252
timestamp 1698175906
transform 1 0 29568 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_268
timestamp 1698175906
transform 1 0 31360 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_276
timestamp 1698175906
transform 1 0 32256 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_282
timestamp 1698175906
transform 1 0 32928 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_346
timestamp 1698175906
transform 1 0 40096 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_348
timestamp 1698175906
transform 1 0 40320 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_2
timestamp 1698175906
transform 1 0 1568 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698175906
transform 1 0 5152 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_37
timestamp 1698175906
transform 1 0 5488 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_69
timestamp 1698175906
transform 1 0 9072 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_73
timestamp 1698175906
transform 1 0 9520 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_75
timestamp 1698175906
transform 1 0 9744 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_107
timestamp 1698175906
transform 1 0 13328 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_148
timestamp 1698175906
transform 1 0 17920 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_172
timestamp 1698175906
transform 1 0 20608 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_174
timestamp 1698175906
transform 1 0 20832 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_215
timestamp 1698175906
transform 1 0 25424 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_224
timestamp 1698175906
transform 1 0 26432 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_234
timestamp 1698175906
transform 1 0 27552 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_242
timestamp 1698175906
transform 1 0 28448 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_244
timestamp 1698175906
transform 1 0 28672 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_247
timestamp 1698175906
transform 1 0 29008 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_311
timestamp 1698175906
transform 1 0 36176 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_317
timestamp 1698175906
transform 1 0 36848 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_321
timestamp 1698175906
transform 1 0 37296 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_2
timestamp 1698175906
transform 1 0 1568 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_66
timestamp 1698175906
transform 1 0 8736 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_72
timestamp 1698175906
transform 1 0 9408 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_80
timestamp 1698175906
transform 1 0 10304 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_111
timestamp 1698175906
transform 1 0 13776 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_127
timestamp 1698175906
transform 1 0 15568 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_129
timestamp 1698175906
transform 1 0 15792 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_136
timestamp 1698175906
transform 1 0 16576 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_142
timestamp 1698175906
transform 1 0 17248 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_150
timestamp 1698175906
transform 1 0 18144 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_154
timestamp 1698175906
transform 1 0 18592 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_156
timestamp 1698175906
transform 1 0 18816 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_209
timestamp 1698175906
transform 1 0 24752 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_212
timestamp 1698175906
transform 1 0 25088 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_245
timestamp 1698175906
transform 1 0 28784 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_249
timestamp 1698175906
transform 1 0 29232 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_265
timestamp 1698175906
transform 1 0 31024 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_273
timestamp 1698175906
transform 1 0 31920 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_277
timestamp 1698175906
transform 1 0 32368 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_279
timestamp 1698175906
transform 1 0 32592 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_282
timestamp 1698175906
transform 1 0 32928 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_314
timestamp 1698175906
transform 1 0 36512 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_322
timestamp 1698175906
transform 1 0 37408 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_2
timestamp 1698175906
transform 1 0 1568 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698175906
transform 1 0 5152 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_37
timestamp 1698175906
transform 1 0 5488 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_101
timestamp 1698175906
transform 1 0 12656 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_113
timestamp 1698175906
transform 1 0 14000 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_121
timestamp 1698175906
transform 1 0 14896 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_183
timestamp 1698175906
transform 1 0 21840 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_187
timestamp 1698175906
transform 1 0 22288 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_247
timestamp 1698175906
transform 1 0 29008 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_260
timestamp 1698175906
transform 1 0 30464 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_292
timestamp 1698175906
transform 1 0 34048 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_308
timestamp 1698175906
transform 1 0 35840 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_312
timestamp 1698175906
transform 1 0 36288 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_314
timestamp 1698175906
transform 1 0 36512 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_317
timestamp 1698175906
transform 1 0 36848 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_321
timestamp 1698175906
transform 1 0 37296 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_2
timestamp 1698175906
transform 1 0 1568 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_66
timestamp 1698175906
transform 1 0 8736 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_72
timestamp 1698175906
transform 1 0 9408 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_115
timestamp 1698175906
transform 1 0 14224 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_131
timestamp 1698175906
transform 1 0 16016 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_139
timestamp 1698175906
transform 1 0 16912 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_142
timestamp 1698175906
transform 1 0 17248 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_146
timestamp 1698175906
transform 1 0 17696 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_154
timestamp 1698175906
transform 1 0 18592 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_170
timestamp 1698175906
transform 1 0 20384 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_176
timestamp 1698175906
transform 1 0 21056 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_180
timestamp 1698175906
transform 1 0 21504 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_190
timestamp 1698175906
transform 1 0 22624 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_194
timestamp 1698175906
transform 1 0 23072 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_208
timestamp 1698175906
transform 1 0 24640 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_212
timestamp 1698175906
transform 1 0 25088 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_214
timestamp 1698175906
transform 1 0 25312 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_221
timestamp 1698175906
transform 1 0 26096 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_254
timestamp 1698175906
transform 1 0 29792 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_270
timestamp 1698175906
transform 1 0 31584 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_278
timestamp 1698175906
transform 1 0 32480 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_282
timestamp 1698175906
transform 1 0 32928 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_314
timestamp 1698175906
transform 1 0 36512 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_322
timestamp 1698175906
transform 1 0 37408 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_28
timestamp 1698175906
transform 1 0 4480 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_32
timestamp 1698175906
transform 1 0 4928 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698175906
transform 1 0 5152 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_37
timestamp 1698175906
transform 1 0 5488 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_69
timestamp 1698175906
transform 1 0 9072 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_73
timestamp 1698175906
transform 1 0 9520 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_75
timestamp 1698175906
transform 1 0 9744 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_112
timestamp 1698175906
transform 1 0 13888 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_116
timestamp 1698175906
transform 1 0 14336 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_124
timestamp 1698175906
transform 1 0 15232 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_128
timestamp 1698175906
transform 1 0 15680 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_147
timestamp 1698175906
transform 1 0 17808 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_160
timestamp 1698175906
transform 1 0 19264 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_168
timestamp 1698175906
transform 1 0 20160 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_172
timestamp 1698175906
transform 1 0 20608 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_174
timestamp 1698175906
transform 1 0 20832 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_177
timestamp 1698175906
transform 1 0 21168 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_181
timestamp 1698175906
transform 1 0 21616 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_211
timestamp 1698175906
transform 1 0 24976 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_215
timestamp 1698175906
transform 1 0 25424 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_228
timestamp 1698175906
transform 1 0 26880 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_230
timestamp 1698175906
transform 1 0 27104 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_236
timestamp 1698175906
transform 1 0 27776 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_244
timestamp 1698175906
transform 1 0 28672 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_247
timestamp 1698175906
transform 1 0 29008 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_311
timestamp 1698175906
transform 1 0 36176 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_317
timestamp 1698175906
transform 1 0 36848 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_321
timestamp 1698175906
transform 1 0 37296 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_28
timestamp 1698175906
transform 1 0 4480 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_60
timestamp 1698175906
transform 1 0 8064 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_68
timestamp 1698175906
transform 1 0 8960 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_72
timestamp 1698175906
transform 1 0 9408 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_104
timestamp 1698175906
transform 1 0 12992 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_108
timestamp 1698175906
transform 1 0 13440 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_110
timestamp 1698175906
transform 1 0 13664 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_142
timestamp 1698175906
transform 1 0 17248 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_162
timestamp 1698175906
transform 1 0 19488 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_178
timestamp 1698175906
transform 1 0 21280 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_182
timestamp 1698175906
transform 1 0 21728 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_193
timestamp 1698175906
transform 1 0 22960 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_209
timestamp 1698175906
transform 1 0 24752 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_212
timestamp 1698175906
transform 1 0 25088 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_225
timestamp 1698175906
transform 1 0 26544 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_257
timestamp 1698175906
transform 1 0 30128 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_273
timestamp 1698175906
transform 1 0 31920 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_277
timestamp 1698175906
transform 1 0 32368 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_279
timestamp 1698175906
transform 1 0 32592 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_282
timestamp 1698175906
transform 1 0 32928 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_346
timestamp 1698175906
transform 1 0 40096 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_348
timestamp 1698175906
transform 1 0 40320 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_2
timestamp 1698175906
transform 1 0 1568 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698175906
transform 1 0 5152 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_37
timestamp 1698175906
transform 1 0 5488 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_107
timestamp 1698175906
transform 1 0 13328 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_111
timestamp 1698175906
transform 1 0 13776 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_113
timestamp 1698175906
transform 1 0 14000 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_116
timestamp 1698175906
transform 1 0 14336 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_124
timestamp 1698175906
transform 1 0 15232 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_132
timestamp 1698175906
transform 1 0 16128 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_148
timestamp 1698175906
transform 1 0 17920 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_158
timestamp 1698175906
transform 1 0 19040 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_166
timestamp 1698175906
transform 1 0 19936 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_194
timestamp 1698175906
transform 1 0 23072 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_205
timestamp 1698175906
transform 1 0 24304 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_213
timestamp 1698175906
transform 1 0 25200 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_215
timestamp 1698175906
transform 1 0 25424 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_247
timestamp 1698175906
transform 1 0 29008 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_251
timestamp 1698175906
transform 1 0 29456 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_317
timestamp 1698175906
transform 1 0 36848 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_2
timestamp 1698175906
transform 1 0 1568 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_66
timestamp 1698175906
transform 1 0 8736 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_72
timestamp 1698175906
transform 1 0 9408 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_80
timestamp 1698175906
transform 1 0 10304 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_84
timestamp 1698175906
transform 1 0 10752 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_123
timestamp 1698175906
transform 1 0 15120 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_139
timestamp 1698175906
transform 1 0 16912 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_147
timestamp 1698175906
transform 1 0 17808 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_156
timestamp 1698175906
transform 1 0 18816 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_160
timestamp 1698175906
transform 1 0 19264 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_168
timestamp 1698175906
transform 1 0 20160 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_198
timestamp 1698175906
transform 1 0 23520 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_202
timestamp 1698175906
transform 1 0 23968 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_212
timestamp 1698175906
transform 1 0 25088 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_219
timestamp 1698175906
transform 1 0 25872 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_226
timestamp 1698175906
transform 1 0 26656 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_241
timestamp 1698175906
transform 1 0 28336 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_273
timestamp 1698175906
transform 1 0 31920 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_277
timestamp 1698175906
transform 1 0 32368 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_279
timestamp 1698175906
transform 1 0 32592 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_282
timestamp 1698175906
transform 1 0 32928 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_314
timestamp 1698175906
transform 1 0 36512 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_322
timestamp 1698175906
transform 1 0 37408 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_28
timestamp 1698175906
transform 1 0 4480 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_32
timestamp 1698175906
transform 1 0 4928 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698175906
transform 1 0 5152 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_37
timestamp 1698175906
transform 1 0 5488 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_101
timestamp 1698175906
transform 1 0 12656 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_111
timestamp 1698175906
transform 1 0 13776 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_124
timestamp 1698175906
transform 1 0 15232 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_168
timestamp 1698175906
transform 1 0 20160 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_172
timestamp 1698175906
transform 1 0 20608 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_174
timestamp 1698175906
transform 1 0 20832 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_177
timestamp 1698175906
transform 1 0 21168 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_181
timestamp 1698175906
transform 1 0 21616 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_240
timestamp 1698175906
transform 1 0 28224 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_244
timestamp 1698175906
transform 1 0 28672 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_247
timestamp 1698175906
transform 1 0 29008 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_311
timestamp 1698175906
transform 1 0 36176 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_317
timestamp 1698175906
transform 1 0 36848 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_321
timestamp 1698175906
transform 1 0 37296 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_28
timestamp 1698175906
transform 1 0 4480 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_60
timestamp 1698175906
transform 1 0 8064 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_68
timestamp 1698175906
transform 1 0 8960 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_72
timestamp 1698175906
transform 1 0 9408 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_88
timestamp 1698175906
transform 1 0 11200 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_127
timestamp 1698175906
transform 1 0 15568 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_131
timestamp 1698175906
transform 1 0 16016 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_139
timestamp 1698175906
transform 1 0 16912 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_142
timestamp 1698175906
transform 1 0 17248 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_150
timestamp 1698175906
transform 1 0 18144 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_154
timestamp 1698175906
transform 1 0 18592 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_159
timestamp 1698175906
transform 1 0 19152 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_167
timestamp 1698175906
transform 1 0 20048 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_199
timestamp 1698175906
transform 1 0 23632 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_207
timestamp 1698175906
transform 1 0 24528 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_209
timestamp 1698175906
transform 1 0 24752 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_212
timestamp 1698175906
transform 1 0 25088 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_216
timestamp 1698175906
transform 1 0 25536 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_282
timestamp 1698175906
transform 1 0 32928 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_314
timestamp 1698175906
transform 1 0 36512 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_322
timestamp 1698175906
transform 1 0 37408 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_28
timestamp 1698175906
transform 1 0 4480 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_32
timestamp 1698175906
transform 1 0 4928 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698175906
transform 1 0 5152 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_37
timestamp 1698175906
transform 1 0 5488 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_101
timestamp 1698175906
transform 1 0 12656 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_107
timestamp 1698175906
transform 1 0 13328 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_111
timestamp 1698175906
transform 1 0 13776 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_119
timestamp 1698175906
transform 1 0 14672 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_135
timestamp 1698175906
transform 1 0 16464 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_139
timestamp 1698175906
transform 1 0 16912 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_170
timestamp 1698175906
transform 1 0 20384 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_174
timestamp 1698175906
transform 1 0 20832 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_177
timestamp 1698175906
transform 1 0 21168 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_241
timestamp 1698175906
transform 1 0 28336 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_247
timestamp 1698175906
transform 1 0 29008 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_311
timestamp 1698175906
transform 1 0 36176 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_317
timestamp 1698175906
transform 1 0 36848 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_28
timestamp 1698175906
transform 1 0 4480 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_60
timestamp 1698175906
transform 1 0 8064 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_68
timestamp 1698175906
transform 1 0 8960 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_72
timestamp 1698175906
transform 1 0 9408 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_136
timestamp 1698175906
transform 1 0 16576 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_142
timestamp 1698175906
transform 1 0 17248 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_206
timestamp 1698175906
transform 1 0 24416 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_212
timestamp 1698175906
transform 1 0 25088 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_276
timestamp 1698175906
transform 1 0 32256 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_282
timestamp 1698175906
transform 1 0 32928 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_346
timestamp 1698175906
transform 1 0 40096 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_348
timestamp 1698175906
transform 1 0 40320 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_2
timestamp 1698175906
transform 1 0 1568 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698175906
transform 1 0 5152 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_37
timestamp 1698175906
transform 1 0 5488 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_101
timestamp 1698175906
transform 1 0 12656 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_107
timestamp 1698175906
transform 1 0 13328 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_171
timestamp 1698175906
transform 1 0 20496 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_177
timestamp 1698175906
transform 1 0 21168 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_241
timestamp 1698175906
transform 1 0 28336 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_247
timestamp 1698175906
transform 1 0 29008 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_311
timestamp 1698175906
transform 1 0 36176 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_317
timestamp 1698175906
transform 1 0 36848 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_2
timestamp 1698175906
transform 1 0 1568 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_66
timestamp 1698175906
transform 1 0 8736 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_72
timestamp 1698175906
transform 1 0 9408 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_136
timestamp 1698175906
transform 1 0 16576 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_142
timestamp 1698175906
transform 1 0 17248 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_206
timestamp 1698175906
transform 1 0 24416 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_212
timestamp 1698175906
transform 1 0 25088 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_276
timestamp 1698175906
transform 1 0 32256 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_282
timestamp 1698175906
transform 1 0 32928 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_346
timestamp 1698175906
transform 1 0 40096 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_348
timestamp 1698175906
transform 1 0 40320 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698175906
transform 1 0 1568 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698175906
transform 1 0 5152 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_37
timestamp 1698175906
transform 1 0 5488 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_101
timestamp 1698175906
transform 1 0 12656 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_107
timestamp 1698175906
transform 1 0 13328 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_171
timestamp 1698175906
transform 1 0 20496 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_177
timestamp 1698175906
transform 1 0 21168 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_241
timestamp 1698175906
transform 1 0 28336 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_247
timestamp 1698175906
transform 1 0 29008 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_311
timestamp 1698175906
transform 1 0 36176 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_317
timestamp 1698175906
transform 1 0 36848 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2
timestamp 1698175906
transform 1 0 1568 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_66
timestamp 1698175906
transform 1 0 8736 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_72
timestamp 1698175906
transform 1 0 9408 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_136
timestamp 1698175906
transform 1 0 16576 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_142
timestamp 1698175906
transform 1 0 17248 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_206
timestamp 1698175906
transform 1 0 24416 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_212
timestamp 1698175906
transform 1 0 25088 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_276
timestamp 1698175906
transform 1 0 32256 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_282
timestamp 1698175906
transform 1 0 32928 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_346
timestamp 1698175906
transform 1 0 40096 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_348
timestamp 1698175906
transform 1 0 40320 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_2
timestamp 1698175906
transform 1 0 1568 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698175906
transform 1 0 5152 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_37
timestamp 1698175906
transform 1 0 5488 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_101
timestamp 1698175906
transform 1 0 12656 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_107
timestamp 1698175906
transform 1 0 13328 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_171
timestamp 1698175906
transform 1 0 20496 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_177
timestamp 1698175906
transform 1 0 21168 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_241
timestamp 1698175906
transform 1 0 28336 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_247
timestamp 1698175906
transform 1 0 29008 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_311
timestamp 1698175906
transform 1 0 36176 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_317
timestamp 1698175906
transform 1 0 36848 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2
timestamp 1698175906
transform 1 0 1568 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_66
timestamp 1698175906
transform 1 0 8736 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_72
timestamp 1698175906
transform 1 0 9408 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_136
timestamp 1698175906
transform 1 0 16576 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_142
timestamp 1698175906
transform 1 0 17248 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_206
timestamp 1698175906
transform 1 0 24416 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_212
timestamp 1698175906
transform 1 0 25088 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_276
timestamp 1698175906
transform 1 0 32256 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_282
timestamp 1698175906
transform 1 0 32928 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_346
timestamp 1698175906
transform 1 0 40096 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_348
timestamp 1698175906
transform 1 0 40320 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698175906
transform 1 0 1568 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698175906
transform 1 0 5152 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_37
timestamp 1698175906
transform 1 0 5488 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_101
timestamp 1698175906
transform 1 0 12656 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_107
timestamp 1698175906
transform 1 0 13328 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_171
timestamp 1698175906
transform 1 0 20496 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_177
timestamp 1698175906
transform 1 0 21168 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_241
timestamp 1698175906
transform 1 0 28336 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_247
timestamp 1698175906
transform 1 0 29008 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_311
timestamp 1698175906
transform 1 0 36176 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_317
timestamp 1698175906
transform 1 0 36848 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_2
timestamp 1698175906
transform 1 0 1568 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_66
timestamp 1698175906
transform 1 0 8736 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_72
timestamp 1698175906
transform 1 0 9408 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_136
timestamp 1698175906
transform 1 0 16576 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_142
timestamp 1698175906
transform 1 0 17248 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_206
timestamp 1698175906
transform 1 0 24416 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_212
timestamp 1698175906
transform 1 0 25088 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_276
timestamp 1698175906
transform 1 0 32256 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_282
timestamp 1698175906
transform 1 0 32928 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_346
timestamp 1698175906
transform 1 0 40096 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_348
timestamp 1698175906
transform 1 0 40320 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698175906
transform 1 0 1568 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698175906
transform 1 0 5152 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_37
timestamp 1698175906
transform 1 0 5488 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_101
timestamp 1698175906
transform 1 0 12656 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_107
timestamp 1698175906
transform 1 0 13328 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_171
timestamp 1698175906
transform 1 0 20496 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_177
timestamp 1698175906
transform 1 0 21168 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_241
timestamp 1698175906
transform 1 0 28336 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_247
timestamp 1698175906
transform 1 0 29008 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_311
timestamp 1698175906
transform 1 0 36176 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_317
timestamp 1698175906
transform 1 0 36848 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2
timestamp 1698175906
transform 1 0 1568 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1698175906
transform 1 0 8736 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_72
timestamp 1698175906
transform 1 0 9408 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_136
timestamp 1698175906
transform 1 0 16576 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_142
timestamp 1698175906
transform 1 0 17248 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_206
timestamp 1698175906
transform 1 0 24416 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_212
timestamp 1698175906
transform 1 0 25088 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_276
timestamp 1698175906
transform 1 0 32256 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_282
timestamp 1698175906
transform 1 0 32928 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_346
timestamp 1698175906
transform 1 0 40096 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_348
timestamp 1698175906
transform 1 0 40320 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_2
timestamp 1698175906
transform 1 0 1568 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698175906
transform 1 0 5152 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_37
timestamp 1698175906
transform 1 0 5488 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_101
timestamp 1698175906
transform 1 0 12656 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_107
timestamp 1698175906
transform 1 0 13328 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_139
timestamp 1698175906
transform 1 0 16912 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_155
timestamp 1698175906
transform 1 0 18704 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_167
timestamp 1698175906
transform 1 0 20048 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_177
timestamp 1698175906
transform 1 0 21168 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_241
timestamp 1698175906
transform 1 0 28336 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_247
timestamp 1698175906
transform 1 0 29008 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_311
timestamp 1698175906
transform 1 0 36176 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_317
timestamp 1698175906
transform 1 0 36848 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_2
timestamp 1698175906
transform 1 0 1568 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_66
timestamp 1698175906
transform 1 0 8736 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_72
timestamp 1698175906
transform 1 0 9408 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_136
timestamp 1698175906
transform 1 0 16576 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_142
timestamp 1698175906
transform 1 0 17248 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_150
timestamp 1698175906
transform 1 0 18144 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_154
timestamp 1698175906
transform 1 0 18592 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_156
timestamp 1698175906
transform 1 0 18816 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_183
timestamp 1698175906
transform 1 0 21840 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_199
timestamp 1698175906
transform 1 0 23632 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_207
timestamp 1698175906
transform 1 0 24528 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_209
timestamp 1698175906
transform 1 0 24752 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_238
timestamp 1698175906
transform 1 0 28000 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_270
timestamp 1698175906
transform 1 0 31584 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_278
timestamp 1698175906
transform 1 0 32480 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_282
timestamp 1698175906
transform 1 0 32928 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_346
timestamp 1698175906
transform 1 0 40096 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_348
timestamp 1698175906
transform 1 0 40320 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_2
timestamp 1698175906
transform 1 0 1568 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_36
timestamp 1698175906
transform 1 0 5376 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_70
timestamp 1698175906
transform 1 0 9184 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_104
timestamp 1698175906
transform 1 0 12992 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_138
timestamp 1698175906
transform 1 0 16800 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_142
timestamp 1698175906
transform 1 0 17248 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_198
timestamp 1698175906
transform 1 0 23520 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_202
timestamp 1698175906
transform 1 0 23968 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_232
timestamp 1698175906
transform 1 0 27328 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_236
timestamp 1698175906
transform 1 0 27776 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_240
timestamp 1698175906
transform 1 0 28224 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_274
timestamp 1698175906
transform 1 0 32032 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_308
timestamp 1698175906
transform 1 0 35840 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_342
timestamp 1698175906
transform 1 0 39648 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_346
timestamp 1698175906
transform 1 0 40096 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_348
timestamp 1698175906
transform 1 0 40320 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita41_25 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 39984 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita41_26
timestamp 1698175906
transform -1 0 20048 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 37520 0 1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output2
timestamp 1698175906
transform -1 0 4480 0 1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output3
timestamp 1698175906
transform -1 0 4480 0 1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output4
timestamp 1698175906
transform 1 0 24416 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output5
timestamp 1698175906
transform -1 0 4480 0 -1 28224
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output6
timestamp 1698175906
transform 1 0 37520 0 -1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output7
timestamp 1698175906
transform -1 0 4480 0 -1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output8
timestamp 1698175906
transform 1 0 37520 0 -1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output9
timestamp 1698175906
transform 1 0 37520 0 1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output10
timestamp 1698175906
transform -1 0 20384 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output11
timestamp 1698175906
transform 1 0 20608 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output12
timestamp 1698175906
transform 1 0 18928 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output13
timestamp 1698175906
transform -1 0 4480 0 1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output14
timestamp 1698175906
transform 1 0 37520 0 1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output15
timestamp 1698175906
transform -1 0 4480 0 -1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output16
timestamp 1698175906
transform 1 0 24416 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output17
timestamp 1698175906
transform 1 0 37520 0 -1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output18
timestamp 1698175906
transform -1 0 24192 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output19
timestamp 1698175906
transform 1 0 37520 0 1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output20
timestamp 1698175906
transform 1 0 37520 0 -1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output21
timestamp 1698175906
transform 1 0 25088 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output22
timestamp 1698175906
transform 1 0 37520 0 -1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output23
timestamp 1698175906
transform -1 0 4480 0 1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output24
timestamp 1698175906
transform -1 0 4480 0 -1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_45 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698175906
transform -1 0 40656 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_46
timestamp 1698175906
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698175906
transform -1 0 40656 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_47
timestamp 1698175906
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698175906
transform -1 0 40656 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_48
timestamp 1698175906
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698175906
transform -1 0 40656 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_49
timestamp 1698175906
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698175906
transform -1 0 40656 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_50
timestamp 1698175906
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698175906
transform -1 0 40656 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_51
timestamp 1698175906
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698175906
transform -1 0 40656 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_52
timestamp 1698175906
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698175906
transform -1 0 40656 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_53
timestamp 1698175906
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698175906
transform -1 0 40656 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_54
timestamp 1698175906
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698175906
transform -1 0 40656 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_55
timestamp 1698175906
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698175906
transform -1 0 40656 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_56
timestamp 1698175906
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698175906
transform -1 0 40656 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_57
timestamp 1698175906
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698175906
transform -1 0 40656 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_58
timestamp 1698175906
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698175906
transform -1 0 40656 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_59
timestamp 1698175906
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698175906
transform -1 0 40656 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_60
timestamp 1698175906
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698175906
transform -1 0 40656 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_61
timestamp 1698175906
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698175906
transform -1 0 40656 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_62
timestamp 1698175906
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698175906
transform -1 0 40656 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_63
timestamp 1698175906
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698175906
transform -1 0 40656 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_64
timestamp 1698175906
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698175906
transform -1 0 40656 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_65
timestamp 1698175906
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698175906
transform -1 0 40656 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_66
timestamp 1698175906
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698175906
transform -1 0 40656 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_67
timestamp 1698175906
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698175906
transform -1 0 40656 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_68
timestamp 1698175906
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698175906
transform -1 0 40656 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_69
timestamp 1698175906
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698175906
transform -1 0 40656 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_70
timestamp 1698175906
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698175906
transform -1 0 40656 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_71
timestamp 1698175906
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698175906
transform -1 0 40656 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_72
timestamp 1698175906
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698175906
transform -1 0 40656 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_73
timestamp 1698175906
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698175906
transform -1 0 40656 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_74
timestamp 1698175906
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698175906
transform -1 0 40656 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_75
timestamp 1698175906
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698175906
transform -1 0 40656 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_76
timestamp 1698175906
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698175906
transform -1 0 40656 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_77
timestamp 1698175906
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698175906
transform -1 0 40656 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_78
timestamp 1698175906
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698175906
transform -1 0 40656 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_79
timestamp 1698175906
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698175906
transform -1 0 40656 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_80
timestamp 1698175906
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698175906
transform -1 0 40656 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_81
timestamp 1698175906
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698175906
transform -1 0 40656 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_82
timestamp 1698175906
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698175906
transform -1 0 40656 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_83
timestamp 1698175906
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698175906
transform -1 0 40656 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_84
timestamp 1698175906
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698175906
transform -1 0 40656 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_85
timestamp 1698175906
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698175906
transform -1 0 40656 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_86
timestamp 1698175906
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698175906
transform -1 0 40656 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_87
timestamp 1698175906
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698175906
transform -1 0 40656 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_88
timestamp 1698175906
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698175906
transform -1 0 40656 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_89
timestamp 1698175906
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698175906
transform -1 0 40656 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_90 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_91
timestamp 1698175906
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_92
timestamp 1698175906
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_93
timestamp 1698175906
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_94
timestamp 1698175906
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_95
timestamp 1698175906
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_96
timestamp 1698175906
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_97
timestamp 1698175906
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_98
timestamp 1698175906
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_99
timestamp 1698175906
transform 1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_100
timestamp 1698175906
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_101
timestamp 1698175906
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_102
timestamp 1698175906
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_103
timestamp 1698175906
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_104
timestamp 1698175906
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_105
timestamp 1698175906
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_106
timestamp 1698175906
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_107
timestamp 1698175906
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_108
timestamp 1698175906
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_109
timestamp 1698175906
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_110
timestamp 1698175906
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_111
timestamp 1698175906
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_112
timestamp 1698175906
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_113
timestamp 1698175906
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_114
timestamp 1698175906
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_115
timestamp 1698175906
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_116
timestamp 1698175906
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_117
timestamp 1698175906
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_118
timestamp 1698175906
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_119
timestamp 1698175906
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_120
timestamp 1698175906
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_121
timestamp 1698175906
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_122
timestamp 1698175906
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_123
timestamp 1698175906
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_124
timestamp 1698175906
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_125
timestamp 1698175906
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_126
timestamp 1698175906
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_127
timestamp 1698175906
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_128
timestamp 1698175906
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_129
timestamp 1698175906
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_130
timestamp 1698175906
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_131
timestamp 1698175906
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_132
timestamp 1698175906
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_133
timestamp 1698175906
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_134
timestamp 1698175906
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_135
timestamp 1698175906
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_136
timestamp 1698175906
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_137
timestamp 1698175906
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_138
timestamp 1698175906
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_139
timestamp 1698175906
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_140
timestamp 1698175906
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_141
timestamp 1698175906
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_142
timestamp 1698175906
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_143
timestamp 1698175906
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_144
timestamp 1698175906
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_145
timestamp 1698175906
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_146
timestamp 1698175906
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_147
timestamp 1698175906
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_148
timestamp 1698175906
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_149
timestamp 1698175906
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_150
timestamp 1698175906
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_151
timestamp 1698175906
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_152
timestamp 1698175906
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_153
timestamp 1698175906
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_154
timestamp 1698175906
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_155
timestamp 1698175906
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_156
timestamp 1698175906
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_157
timestamp 1698175906
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_158
timestamp 1698175906
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_159
timestamp 1698175906
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_160
timestamp 1698175906
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_161
timestamp 1698175906
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_162
timestamp 1698175906
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_163
timestamp 1698175906
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_164
timestamp 1698175906
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_165
timestamp 1698175906
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_166
timestamp 1698175906
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_167
timestamp 1698175906
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_168
timestamp 1698175906
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_169
timestamp 1698175906
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_170
timestamp 1698175906
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_171
timestamp 1698175906
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_172
timestamp 1698175906
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_173
timestamp 1698175906
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_174
timestamp 1698175906
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_175
timestamp 1698175906
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_176
timestamp 1698175906
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_177
timestamp 1698175906
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_178
timestamp 1698175906
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_179
timestamp 1698175906
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_180
timestamp 1698175906
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_181
timestamp 1698175906
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_182
timestamp 1698175906
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_183
timestamp 1698175906
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_184
timestamp 1698175906
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_185
timestamp 1698175906
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_186
timestamp 1698175906
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_187
timestamp 1698175906
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_188
timestamp 1698175906
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_189
timestamp 1698175906
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_190
timestamp 1698175906
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_191
timestamp 1698175906
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_192
timestamp 1698175906
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_193
timestamp 1698175906
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_194
timestamp 1698175906
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_195
timestamp 1698175906
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_196
timestamp 1698175906
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_197
timestamp 1698175906
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_198
timestamp 1698175906
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_199
timestamp 1698175906
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_200
timestamp 1698175906
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_201
timestamp 1698175906
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_202
timestamp 1698175906
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_203
timestamp 1698175906
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_204
timestamp 1698175906
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_205
timestamp 1698175906
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_206
timestamp 1698175906
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_207
timestamp 1698175906
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_208
timestamp 1698175906
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_209
timestamp 1698175906
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_210
timestamp 1698175906
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_211
timestamp 1698175906
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_212
timestamp 1698175906
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_213
timestamp 1698175906
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_214
timestamp 1698175906
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_215
timestamp 1698175906
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_216
timestamp 1698175906
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_217
timestamp 1698175906
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_218
timestamp 1698175906
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_219
timestamp 1698175906
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_220
timestamp 1698175906
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_221
timestamp 1698175906
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_222
timestamp 1698175906
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_223
timestamp 1698175906
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_224
timestamp 1698175906
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_225
timestamp 1698175906
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_226
timestamp 1698175906
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_227
timestamp 1698175906
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_228
timestamp 1698175906
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_229
timestamp 1698175906
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_230
timestamp 1698175906
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_231
timestamp 1698175906
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_232
timestamp 1698175906
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_233
timestamp 1698175906
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_234
timestamp 1698175906
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_235
timestamp 1698175906
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_236
timestamp 1698175906
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_237
timestamp 1698175906
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_238
timestamp 1698175906
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_239
timestamp 1698175906
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_240
timestamp 1698175906
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_241
timestamp 1698175906
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_242
timestamp 1698175906
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_243
timestamp 1698175906
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_244
timestamp 1698175906
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_245
timestamp 1698175906
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_246
timestamp 1698175906
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_247
timestamp 1698175906
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_248
timestamp 1698175906
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_249
timestamp 1698175906
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_250
timestamp 1698175906
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_251
timestamp 1698175906
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_252
timestamp 1698175906
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_253
timestamp 1698175906
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_254
timestamp 1698175906
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_255
timestamp 1698175906
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_256
timestamp 1698175906
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_257
timestamp 1698175906
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_258
timestamp 1698175906
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_259
timestamp 1698175906
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_260
timestamp 1698175906
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_261
timestamp 1698175906
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_262
timestamp 1698175906
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_263
timestamp 1698175906
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_264
timestamp 1698175906
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_265
timestamp 1698175906
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_266
timestamp 1698175906
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_267
timestamp 1698175906
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_268
timestamp 1698175906
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_269
timestamp 1698175906
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_270
timestamp 1698175906
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_271
timestamp 1698175906
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_272
timestamp 1698175906
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_273
timestamp 1698175906
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_274
timestamp 1698175906
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_275
timestamp 1698175906
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_276
timestamp 1698175906
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_277
timestamp 1698175906
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_278
timestamp 1698175906
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_279
timestamp 1698175906
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_280
timestamp 1698175906
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_281
timestamp 1698175906
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_282
timestamp 1698175906
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_283
timestamp 1698175906
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_284
timestamp 1698175906
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_285
timestamp 1698175906
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_286
timestamp 1698175906
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_287
timestamp 1698175906
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_288
timestamp 1698175906
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_289
timestamp 1698175906
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_290
timestamp 1698175906
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_291
timestamp 1698175906
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_292
timestamp 1698175906
transform 1 0 32704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_293
timestamp 1698175906
transform 1 0 5152 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_294
timestamp 1698175906
transform 1 0 8960 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_295
timestamp 1698175906
transform 1 0 12768 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_296
timestamp 1698175906
transform 1 0 16576 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_297
timestamp 1698175906
transform 1 0 20384 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_298
timestamp 1698175906
transform 1 0 24192 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_299
timestamp 1698175906
transform 1 0 28000 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_300
timestamp 1698175906
transform 1 0 31808 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_301
timestamp 1698175906
transform 1 0 35616 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_302
timestamp 1698175906
transform 1 0 39424 0 1 37632
box -86 -86 310 870
<< labels >>
flabel metal3 s 0 24192 800 24304 0 FreeSans 448 0 0 0 clk
port 0 nsew signal input
flabel metal3 s 41200 10080 42000 10192 0 FreeSans 448 0 0 0 segm[0]
port 1 nsew signal tristate
flabel metal3 s 41200 19488 42000 19600 0 FreeSans 448 0 0 0 segm[10]
port 2 nsew signal tristate
flabel metal3 s 0 17472 800 17584 0 FreeSans 448 0 0 0 segm[11]
port 3 nsew signal tristate
flabel metal3 s 0 22176 800 22288 0 FreeSans 448 0 0 0 segm[12]
port 4 nsew signal tristate
flabel metal2 s 22848 41200 22960 42000 0 FreeSans 448 90 0 0 segm[13]
port 5 nsew signal tristate
flabel metal3 s 0 26880 800 26992 0 FreeSans 448 0 0 0 segm[1]
port 6 nsew signal tristate
flabel metal3 s 41200 21504 42000 21616 0 FreeSans 448 0 0 0 segm[2]
port 7 nsew signal tristate
flabel metal2 s 19488 41200 19600 42000 0 FreeSans 448 90 0 0 segm[3]
port 8 nsew signal tristate
flabel metal3 s 0 25536 800 25648 0 FreeSans 448 0 0 0 segm[4]
port 9 nsew signal tristate
flabel metal3 s 41200 20160 42000 20272 0 FreeSans 448 0 0 0 segm[5]
port 10 nsew signal tristate
flabel metal3 s 41200 24864 42000 24976 0 FreeSans 448 0 0 0 segm[6]
port 11 nsew signal tristate
flabel metal2 s 18144 41200 18256 42000 0 FreeSans 448 90 0 0 segm[7]
port 12 nsew signal tristate
flabel metal2 s 20160 41200 20272 42000 0 FreeSans 448 90 0 0 segm[8]
port 13 nsew signal tristate
flabel metal2 s 18816 41200 18928 42000 0 FreeSans 448 90 0 0 segm[9]
port 14 nsew signal tristate
flabel metal3 s 0 24864 800 24976 0 FreeSans 448 0 0 0 sel[0]
port 15 nsew signal tristate
flabel metal3 s 41200 22176 42000 22288 0 FreeSans 448 0 0 0 sel[10]
port 16 nsew signal tristate
flabel metal3 s 0 16128 800 16240 0 FreeSans 448 0 0 0 sel[11]
port 17 nsew signal tristate
flabel metal2 s 22848 0 22960 800 0 FreeSans 448 90 0 0 sel[1]
port 18 nsew signal tristate
flabel metal3 s 41200 24192 42000 24304 0 FreeSans 448 0 0 0 sel[2]
port 19 nsew signal tristate
flabel metal2 s 22176 0 22288 800 0 FreeSans 448 90 0 0 sel[3]
port 20 nsew signal tristate
flabel metal3 s 41200 20832 42000 20944 0 FreeSans 448 0 0 0 sel[4]
port 21 nsew signal tristate
flabel metal3 s 41200 16128 42000 16240 0 FreeSans 448 0 0 0 sel[5]
port 22 nsew signal tristate
flabel metal2 s 24192 41200 24304 42000 0 FreeSans 448 90 0 0 sel[6]
port 23 nsew signal tristate
flabel metal3 s 41200 25536 42000 25648 0 FreeSans 448 0 0 0 sel[7]
port 24 nsew signal tristate
flabel metal3 s 0 26208 800 26320 0 FreeSans 448 0 0 0 sel[8]
port 25 nsew signal tristate
flabel metal3 s 0 22848 800 22960 0 FreeSans 448 0 0 0 sel[9]
port 26 nsew signal tristate
flabel metal4 s 4448 3076 4768 38476 0 FreeSans 1280 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 35168 3076 35488 38476 0 FreeSans 1280 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 19808 3076 20128 38476 0 FreeSans 1280 90 0 0 vss
port 28 nsew ground bidirectional
rlabel metal1 21000 38416 21000 38416 0 vdd
rlabel metal1 21000 37632 21000 37632 0 vss
rlabel metal2 15680 16184 15680 16184 0 _000_
rlabel metal2 22680 24696 22680 24696 0 _001_
rlabel metal2 22008 22008 22008 22008 0 _002_
rlabel metal2 14168 16240 14168 16240 0 _003_
rlabel metal3 16968 24920 16968 24920 0 _004_
rlabel metal2 16128 22456 16128 22456 0 _005_
rlabel metal2 25424 16184 25424 16184 0 _006_
rlabel metal2 20328 18704 20328 18704 0 _007_
rlabel metal3 12488 20552 12488 20552 0 _008_
rlabel metal2 16632 15456 16632 15456 0 _009_
rlabel metal2 27384 17192 27384 17192 0 _010_
rlabel metal2 20440 14840 20440 14840 0 _011_
rlabel metal2 26488 23576 26488 23576 0 _012_
rlabel metal2 21000 15512 21000 15512 0 _013_
rlabel metal2 12936 24360 12936 24360 0 _014_
rlabel metal2 13608 25928 13608 25928 0 _015_
rlabel metal2 19208 26236 19208 26236 0 _016_
rlabel metal2 25816 25144 25816 25144 0 _017_
rlabel metal2 26040 19320 26040 19320 0 _018_
rlabel metal3 12656 21784 12656 21784 0 _019_
rlabel metal2 21280 24584 21280 24584 0 _020_
rlabel metal2 28616 21224 28616 21224 0 _021_
rlabel metal2 23352 23800 23352 23800 0 _022_
rlabel metal3 25480 18984 25480 18984 0 _023_
rlabel metal3 25424 21672 25424 21672 0 _024_
rlabel metal3 27048 20664 27048 20664 0 _025_
rlabel metal2 21560 19544 21560 19544 0 _026_
rlabel metal2 14056 22120 14056 22120 0 _027_
rlabel metal2 22456 19712 22456 19712 0 _028_
rlabel metal3 24304 21336 24304 21336 0 _029_
rlabel metal2 21896 22568 21896 22568 0 _030_
rlabel metal2 22456 23576 22456 23576 0 _031_
rlabel metal2 26768 21000 26768 21000 0 _032_
rlabel metal2 27776 18984 27776 18984 0 _033_
rlabel metal2 17864 17136 17864 17136 0 _034_
rlabel metal3 21672 23912 21672 23912 0 _035_
rlabel metal3 23352 23800 23352 23800 0 _036_
rlabel metal3 21448 21560 21448 21560 0 _037_
rlabel metal2 22568 21504 22568 21504 0 _038_
rlabel metal2 15400 15736 15400 15736 0 _039_
rlabel metal2 17192 23408 17192 23408 0 _040_
rlabel metal3 18144 24808 18144 24808 0 _041_
rlabel metal2 18088 24024 18088 24024 0 _042_
rlabel metal3 16968 22232 16968 22232 0 _043_
rlabel metal3 25200 21560 25200 21560 0 _044_
rlabel metal3 26488 17528 26488 17528 0 _045_
rlabel metal2 15064 19152 15064 19152 0 _046_
rlabel metal2 21504 18424 21504 18424 0 _047_
rlabel metal2 21728 18424 21728 18424 0 _048_
rlabel metal2 22176 18200 22176 18200 0 _049_
rlabel metal2 21840 18984 21840 18984 0 _050_
rlabel metal3 27608 20776 27608 20776 0 _051_
rlabel metal2 14784 20552 14784 20552 0 _052_
rlabel metal2 24024 18816 24024 18816 0 _053_
rlabel metal2 14616 18872 14616 18872 0 _054_
rlabel metal2 13552 20328 13552 20328 0 _055_
rlabel metal2 17080 19488 17080 19488 0 _056_
rlabel metal2 24248 20860 24248 20860 0 _057_
rlabel metal3 21616 18200 21616 18200 0 _058_
rlabel metal2 20552 19208 20552 19208 0 _059_
rlabel metal3 15568 22232 15568 22232 0 _060_
rlabel metal2 15400 17528 15400 17528 0 _061_
rlabel metal3 23408 23128 23408 23128 0 _062_
rlabel metal3 24808 18200 24808 18200 0 _063_
rlabel metal2 26264 17920 26264 17920 0 _064_
rlabel metal2 20608 23912 20608 23912 0 _065_
rlabel metal2 18592 22120 18592 22120 0 _066_
rlabel metal2 19096 22680 19096 22680 0 _067_
rlabel metal2 20720 16296 20720 16296 0 _068_
rlabel metal2 21448 17304 21448 17304 0 _069_
rlabel metal3 21560 16072 21560 16072 0 _070_
rlabel metal2 20720 21000 20720 21000 0 _071_
rlabel metal3 25088 22344 25088 22344 0 _072_
rlabel metal2 26600 22624 26600 22624 0 _073_
rlabel metal2 21448 23800 21448 23800 0 _074_
rlabel metal2 26152 23856 26152 23856 0 _075_
rlabel metal2 21784 17192 21784 17192 0 _076_
rlabel metal2 21896 16352 21896 16352 0 _077_
rlabel metal2 18648 23352 18648 23352 0 _078_
rlabel metal3 21056 24024 21056 24024 0 _079_
rlabel metal2 20216 23576 20216 23576 0 _080_
rlabel metal2 12824 24304 12824 24304 0 _081_
rlabel metal3 14112 25592 14112 25592 0 _082_
rlabel metal2 19992 25424 19992 25424 0 _083_
rlabel metal2 25928 24696 25928 24696 0 _084_
rlabel metal3 23576 21784 23576 21784 0 _085_
rlabel metal2 24584 22400 24584 22400 0 _086_
rlabel metal3 2478 24248 2478 24248 0 clk
rlabel metal3 22288 20776 22288 20776 0 clknet_0_clk
rlabel metal2 12936 22232 12936 22232 0 clknet_1_0__leaf_clk
rlabel metal3 21224 25480 21224 25480 0 clknet_1_1__leaf_clk
rlabel metal2 14504 19208 14504 19208 0 dut41.count\[0\]
rlabel metal2 14392 20440 14392 20440 0 dut41.count\[1\]
rlabel metal2 18536 16016 18536 16016 0 dut41.count\[2\]
rlabel metal2 24808 17416 24808 17416 0 dut41.count\[3\]
rlabel metal3 28056 19880 28056 19880 0 net1
rlabel metal2 18536 25256 18536 25256 0 net10
rlabel metal3 20328 26488 20328 26488 0 net11
rlabel metal3 19208 26936 19208 26936 0 net12
rlabel metal2 4312 25032 4312 25032 0 net13
rlabel metal2 24808 22176 24808 22176 0 net14
rlabel metal2 12040 16016 12040 16016 0 net15
rlabel metal2 24584 5964 24584 5964 0 net16
rlabel metal2 28616 24304 28616 24304 0 net17
rlabel metal2 22568 13552 22568 13552 0 net18
rlabel metal3 31108 20552 31108 20552 0 net19
rlabel metal2 13496 16912 13496 16912 0 net2
rlabel metal2 27048 17360 27048 17360 0 net20
rlabel metal2 24808 26208 24808 26208 0 net21
rlabel metal2 37912 25536 37912 25536 0 net22
rlabel metal2 15064 26768 15064 26768 0 net23
rlabel metal2 13944 23072 13944 23072 0 net24
rlabel metal2 40264 10416 40264 10416 0 net25
rlabel metal2 19544 39942 19544 39942 0 net26
rlabel metal3 6356 22344 6356 22344 0 net3
rlabel metal3 23968 24584 23968 24584 0 net4
rlabel metal2 14168 27384 14168 27384 0 net5
rlabel metal3 29624 20496 29624 20496 0 net6
rlabel metal2 11816 26208 11816 26208 0 net7
rlabel metal3 29680 20776 29680 20776 0 net8
rlabel metal2 28056 25480 28056 25480 0 net9
rlabel metal2 40040 19488 40040 19488 0 segm[10]
rlabel metal3 1358 17528 1358 17528 0 segm[11]
rlabel metal3 1358 22232 1358 22232 0 segm[12]
rlabel metal3 24248 38248 24248 38248 0 segm[13]
rlabel metal3 1358 26936 1358 26936 0 segm[1]
rlabel metal2 40040 21504 40040 21504 0 segm[2]
rlabel metal3 1358 25592 1358 25592 0 segm[4]
rlabel metal3 40642 20216 40642 20216 0 segm[5]
rlabel metal2 40040 25256 40040 25256 0 segm[6]
rlabel metal2 18200 39690 18200 39690 0 segm[7]
rlabel metal3 21000 38248 21000 38248 0 segm[8]
rlabel metal3 19488 37464 19488 37464 0 segm[9]
rlabel metal3 1414 24920 1414 24920 0 sel[0]
rlabel metal2 40040 22344 40040 22344 0 sel[10]
rlabel metal3 1358 16184 1358 16184 0 sel[11]
rlabel metal2 22904 2198 22904 2198 0 sel[1]
rlabel metal2 40040 24360 40040 24360 0 sel[2]
rlabel metal2 22232 2086 22232 2086 0 sel[3]
rlabel metal3 40642 20888 40642 20888 0 sel[4]
rlabel metal2 40040 16408 40040 16408 0 sel[5]
rlabel metal3 25256 37464 25256 37464 0 sel[6]
rlabel metal2 39928 25872 39928 25872 0 sel[7]
rlabel metal3 1414 26264 1414 26264 0 sel[8]
rlabel metal3 1358 22904 1358 22904 0 sel[9]
<< properties >>
string FIXED_BBOX 0 0 42000 42000
<< end >>
