magic
tech gf180mcuD
magscale 1 5
timestamp 1699641407
<< metal1 >>
rect 672 19221 20328 19238
rect 672 19195 2239 19221
rect 2265 19195 2291 19221
rect 2317 19195 2343 19221
rect 2369 19195 17599 19221
rect 17625 19195 17651 19221
rect 17677 19195 17703 19221
rect 17729 19195 20328 19221
rect 672 19178 20328 19195
rect 12783 19137 12809 19143
rect 12783 19105 12809 19111
rect 9081 19055 9087 19081
rect 9113 19055 9119 19081
rect 11097 19055 11103 19081
rect 11129 19055 11135 19081
rect 9865 18999 9871 19025
rect 9897 18999 9903 19025
rect 11993 18999 11999 19025
rect 12025 18999 12031 19025
rect 12273 18999 12279 19025
rect 12305 18999 12311 19025
rect 5839 18969 5865 18975
rect 5839 18937 5865 18943
rect 17599 18969 17625 18975
rect 17599 18937 17625 18943
rect 672 18829 20328 18846
rect 672 18803 9919 18829
rect 9945 18803 9971 18829
rect 9997 18803 10023 18829
rect 10049 18803 20328 18829
rect 672 18786 20328 18803
rect 11047 18745 11073 18751
rect 11047 18713 11073 18719
rect 14071 18745 14097 18751
rect 14071 18713 14097 18719
rect 10537 18607 10543 18633
rect 10569 18607 10575 18633
rect 13561 18607 13567 18633
rect 13593 18607 13599 18633
rect 672 18437 20328 18454
rect 672 18411 2239 18437
rect 2265 18411 2291 18437
rect 2317 18411 2343 18437
rect 2369 18411 17599 18437
rect 17625 18411 17651 18437
rect 17677 18411 17703 18437
rect 17729 18411 20328 18437
rect 672 18394 20328 18411
rect 11159 18353 11185 18359
rect 11159 18321 11185 18327
rect 10649 18215 10655 18241
rect 10681 18215 10687 18241
rect 855 18185 881 18191
rect 855 18153 881 18159
rect 672 18045 20328 18062
rect 672 18019 9919 18045
rect 9945 18019 9971 18045
rect 9997 18019 10023 18045
rect 10049 18019 20328 18045
rect 672 18002 20328 18019
rect 672 17653 20328 17670
rect 672 17627 2239 17653
rect 2265 17627 2291 17653
rect 2317 17627 2343 17653
rect 2369 17627 17599 17653
rect 17625 17627 17651 17653
rect 17677 17627 17703 17653
rect 17729 17627 20328 17653
rect 672 17610 20328 17627
rect 672 17261 20328 17278
rect 672 17235 9919 17261
rect 9945 17235 9971 17261
rect 9997 17235 10023 17261
rect 10049 17235 20328 17261
rect 672 17218 20328 17235
rect 672 16869 20328 16886
rect 672 16843 2239 16869
rect 2265 16843 2291 16869
rect 2317 16843 2343 16869
rect 2369 16843 17599 16869
rect 17625 16843 17651 16869
rect 17677 16843 17703 16869
rect 17729 16843 20328 16869
rect 672 16826 20328 16843
rect 672 16477 20328 16494
rect 672 16451 9919 16477
rect 9945 16451 9971 16477
rect 9997 16451 10023 16477
rect 10049 16451 20328 16477
rect 672 16434 20328 16451
rect 672 16085 20328 16102
rect 672 16059 2239 16085
rect 2265 16059 2291 16085
rect 2317 16059 2343 16085
rect 2369 16059 17599 16085
rect 17625 16059 17651 16085
rect 17677 16059 17703 16085
rect 17729 16059 20328 16085
rect 672 16042 20328 16059
rect 672 15693 20328 15710
rect 672 15667 9919 15693
rect 9945 15667 9971 15693
rect 9997 15667 10023 15693
rect 10049 15667 20328 15693
rect 672 15650 20328 15667
rect 672 15301 20328 15318
rect 672 15275 2239 15301
rect 2265 15275 2291 15301
rect 2317 15275 2343 15301
rect 2369 15275 17599 15301
rect 17625 15275 17651 15301
rect 17677 15275 17703 15301
rect 17729 15275 20328 15301
rect 672 15258 20328 15275
rect 672 14909 20328 14926
rect 672 14883 9919 14909
rect 9945 14883 9971 14909
rect 9997 14883 10023 14909
rect 10049 14883 20328 14909
rect 672 14866 20328 14883
rect 672 14517 20328 14534
rect 672 14491 2239 14517
rect 2265 14491 2291 14517
rect 2317 14491 2343 14517
rect 2369 14491 17599 14517
rect 17625 14491 17651 14517
rect 17677 14491 17703 14517
rect 17729 14491 20328 14517
rect 672 14474 20328 14491
rect 10039 14321 10065 14327
rect 10039 14289 10065 14295
rect 10151 14265 10177 14271
rect 10151 14233 10177 14239
rect 10207 14265 10233 14271
rect 10207 14233 10233 14239
rect 672 14125 20328 14142
rect 672 14099 9919 14125
rect 9945 14099 9971 14125
rect 9997 14099 10023 14125
rect 10049 14099 20328 14125
rect 672 14082 20328 14099
rect 9815 14041 9841 14047
rect 12951 14041 12977 14047
rect 9977 14015 9983 14041
rect 10009 14015 10015 14041
rect 9815 14009 9841 14015
rect 12951 14009 12977 14015
rect 9255 13985 9281 13991
rect 9255 13953 9281 13959
rect 9311 13985 9337 13991
rect 9311 13953 9337 13959
rect 9143 13929 9169 13935
rect 13007 13929 13033 13935
rect 10201 13903 10207 13929
rect 10233 13903 10239 13929
rect 9143 13897 9169 13903
rect 13007 13897 13033 13903
rect 11887 13873 11913 13879
rect 10537 13847 10543 13873
rect 10569 13847 10575 13873
rect 11601 13847 11607 13873
rect 11633 13847 11639 13873
rect 11887 13841 11913 13847
rect 12951 13817 12977 13823
rect 12951 13785 12977 13791
rect 672 13733 20328 13750
rect 672 13707 2239 13733
rect 2265 13707 2291 13733
rect 2317 13707 2343 13733
rect 2369 13707 17599 13733
rect 17625 13707 17651 13733
rect 17677 13707 17703 13733
rect 17729 13707 20328 13733
rect 672 13690 20328 13707
rect 20007 13593 20033 13599
rect 8633 13567 8639 13593
rect 8665 13567 8671 13593
rect 9193 13567 9199 13593
rect 9225 13567 9231 13593
rect 10257 13567 10263 13593
rect 10289 13567 10295 13593
rect 13449 13567 13455 13593
rect 13481 13567 13487 13593
rect 20007 13561 20033 13567
rect 10655 13537 10681 13543
rect 7177 13511 7183 13537
rect 7209 13511 7215 13537
rect 8801 13511 8807 13537
rect 8833 13511 8839 13537
rect 10655 13505 10681 13511
rect 11159 13537 11185 13543
rect 12049 13511 12055 13537
rect 12081 13511 12087 13537
rect 18825 13511 18831 13537
rect 18857 13511 18863 13537
rect 11159 13505 11185 13511
rect 10823 13481 10849 13487
rect 7569 13455 7575 13481
rect 7601 13455 7607 13481
rect 10823 13449 10849 13455
rect 10991 13481 11017 13487
rect 10991 13449 11017 13455
rect 11103 13481 11129 13487
rect 12385 13455 12391 13481
rect 12417 13455 12423 13481
rect 11103 13449 11129 13455
rect 10767 13425 10793 13431
rect 10767 13393 10793 13399
rect 11831 13425 11857 13431
rect 11831 13393 11857 13399
rect 672 13341 20328 13358
rect 672 13315 9919 13341
rect 9945 13315 9971 13341
rect 9997 13315 10023 13341
rect 10049 13315 20328 13341
rect 672 13298 20328 13315
rect 8975 13257 9001 13263
rect 8975 13225 9001 13231
rect 9591 13257 9617 13263
rect 10369 13231 10375 13257
rect 10401 13231 10407 13257
rect 9591 13225 9617 13231
rect 9031 13201 9057 13207
rect 9031 13169 9057 13175
rect 12279 13201 12305 13207
rect 12279 13169 12305 13175
rect 12335 13201 12361 13207
rect 12335 13169 12361 13175
rect 9143 13145 9169 13151
rect 9143 13113 9169 13119
rect 9255 13145 9281 13151
rect 9255 13113 9281 13119
rect 9367 13145 9393 13151
rect 9367 13113 9393 13119
rect 9479 13145 9505 13151
rect 9479 13113 9505 13119
rect 9647 13145 9673 13151
rect 10481 13119 10487 13145
rect 10513 13119 10519 13145
rect 12609 13119 12615 13145
rect 12641 13119 12647 13145
rect 9647 13113 9673 13119
rect 8751 13089 8777 13095
rect 8751 13057 8777 13063
rect 10767 13089 10793 13095
rect 10767 13057 10793 13063
rect 12055 13089 12081 13095
rect 13001 13063 13007 13089
rect 13033 13063 13039 13089
rect 14065 13063 14071 13089
rect 14097 13063 14103 13089
rect 12055 13057 12081 13063
rect 12279 13033 12305 13039
rect 12279 13001 12305 13007
rect 672 12949 20328 12966
rect 672 12923 2239 12949
rect 2265 12923 2291 12949
rect 2317 12923 2343 12949
rect 2369 12923 17599 12949
rect 17625 12923 17651 12949
rect 17677 12923 17703 12949
rect 17729 12923 20328 12949
rect 672 12906 20328 12923
rect 12951 12865 12977 12871
rect 12951 12833 12977 12839
rect 12335 12809 12361 12815
rect 12105 12783 12111 12809
rect 12137 12783 12143 12809
rect 12335 12777 12361 12783
rect 13175 12753 13201 12759
rect 10649 12727 10655 12753
rect 10681 12727 10687 12753
rect 13175 12721 13201 12727
rect 13007 12697 13033 12703
rect 11041 12671 11047 12697
rect 11073 12671 11079 12697
rect 13007 12665 13033 12671
rect 13231 12697 13257 12703
rect 13231 12665 13257 12671
rect 12951 12641 12977 12647
rect 12951 12609 12977 12615
rect 13343 12641 13369 12647
rect 13343 12609 13369 12615
rect 672 12557 20328 12574
rect 672 12531 9919 12557
rect 9945 12531 9971 12557
rect 9997 12531 10023 12557
rect 10049 12531 20328 12557
rect 672 12514 20328 12531
rect 10823 12473 10849 12479
rect 10823 12441 10849 12447
rect 7233 12391 7239 12417
rect 7265 12391 7271 12417
rect 7407 12361 7433 12367
rect 2137 12335 2143 12361
rect 2169 12335 2175 12361
rect 7065 12335 7071 12361
rect 7097 12335 7103 12361
rect 7407 12329 7433 12335
rect 10767 12361 10793 12367
rect 10767 12329 10793 12335
rect 7631 12305 7657 12311
rect 5609 12279 5615 12305
rect 5641 12279 5647 12305
rect 6673 12279 6679 12305
rect 6705 12279 6711 12305
rect 7631 12273 7657 12279
rect 967 12249 993 12255
rect 967 12217 993 12223
rect 10823 12249 10849 12255
rect 10823 12217 10849 12223
rect 672 12165 20328 12182
rect 672 12139 2239 12165
rect 2265 12139 2291 12165
rect 2317 12139 2343 12165
rect 2369 12139 17599 12165
rect 17625 12139 17651 12165
rect 17677 12139 17703 12165
rect 17729 12139 20328 12165
rect 672 12122 20328 12139
rect 11047 12081 11073 12087
rect 11047 12049 11073 12055
rect 11103 12081 11129 12087
rect 11103 12049 11129 12055
rect 9927 12025 9953 12031
rect 9361 11999 9367 12025
rect 9393 11999 9399 12025
rect 9927 11993 9953 11999
rect 20007 12025 20033 12031
rect 20007 11993 20033 11999
rect 6679 11969 6705 11975
rect 6679 11937 6705 11943
rect 7127 11969 7153 11975
rect 10711 11969 10737 11975
rect 7961 11943 7967 11969
rect 7993 11943 7999 11969
rect 7127 11937 7153 11943
rect 10711 11937 10737 11943
rect 10823 11969 10849 11975
rect 10823 11937 10849 11943
rect 11047 11969 11073 11975
rect 18825 11943 18831 11969
rect 18857 11943 18863 11969
rect 11047 11937 11073 11943
rect 6847 11913 6873 11919
rect 9535 11913 9561 11919
rect 8297 11887 8303 11913
rect 8329 11887 8335 11913
rect 6847 11881 6873 11887
rect 9535 11881 9561 11887
rect 9703 11913 9729 11919
rect 9703 11881 9729 11887
rect 13455 11913 13481 11919
rect 13455 11881 13481 11887
rect 13511 11913 13537 11919
rect 13511 11881 13537 11887
rect 6791 11857 6817 11863
rect 6791 11825 6817 11831
rect 6959 11857 6985 11863
rect 6959 11825 6985 11831
rect 7071 11857 7097 11863
rect 7071 11825 7097 11831
rect 13343 11857 13369 11863
rect 13343 11825 13369 11831
rect 672 11773 20328 11790
rect 672 11747 9919 11773
rect 9945 11747 9971 11773
rect 9997 11747 10023 11773
rect 10049 11747 20328 11773
rect 672 11730 20328 11747
rect 8751 11689 8777 11695
rect 8751 11657 8777 11663
rect 9311 11633 9337 11639
rect 10929 11607 10935 11633
rect 10961 11607 10967 11633
rect 14625 11607 14631 11633
rect 14657 11607 14663 11633
rect 9311 11601 9337 11607
rect 8359 11577 8385 11583
rect 6729 11551 6735 11577
rect 6761 11551 6767 11577
rect 8359 11545 8385 11551
rect 8695 11577 8721 11583
rect 8695 11545 8721 11551
rect 8807 11577 8833 11583
rect 8807 11545 8833 11551
rect 9031 11577 9057 11583
rect 9031 11545 9057 11551
rect 9143 11577 9169 11583
rect 9753 11551 9759 11577
rect 9785 11551 9791 11577
rect 12833 11551 12839 11577
rect 12865 11551 12871 11577
rect 14513 11551 14519 11577
rect 14545 11551 14551 11577
rect 18825 11551 18831 11577
rect 18857 11551 18863 11577
rect 9143 11545 9169 11551
rect 12671 11521 12697 11527
rect 7065 11495 7071 11521
rect 7097 11495 7103 11521
rect 8129 11495 8135 11521
rect 8161 11495 8167 11521
rect 13225 11495 13231 11521
rect 13257 11495 13263 11521
rect 14289 11495 14295 11521
rect 14321 11495 14327 11521
rect 12671 11489 12697 11495
rect 8415 11465 8441 11471
rect 8415 11433 8441 11439
rect 20007 11465 20033 11471
rect 20007 11433 20033 11439
rect 672 11381 20328 11398
rect 672 11355 2239 11381
rect 2265 11355 2291 11381
rect 2317 11355 2343 11381
rect 2369 11355 17599 11381
rect 17625 11355 17651 11381
rect 17677 11355 17703 11381
rect 17729 11355 20328 11381
rect 672 11338 20328 11355
rect 8471 11297 8497 11303
rect 8471 11265 8497 11271
rect 7967 11241 7993 11247
rect 7967 11209 7993 11215
rect 8247 11241 8273 11247
rect 12783 11241 12809 11247
rect 13455 11241 13481 11247
rect 10873 11215 10879 11241
rect 10905 11215 10911 11241
rect 13057 11215 13063 11241
rect 13089 11215 13095 11241
rect 8247 11209 8273 11215
rect 12783 11209 12809 11215
rect 13455 11209 13481 11215
rect 20007 11241 20033 11247
rect 20007 11209 20033 11215
rect 7687 11185 7713 11191
rect 9367 11185 9393 11191
rect 10319 11185 10345 11191
rect 12559 11185 12585 11191
rect 9025 11159 9031 11185
rect 9057 11159 9063 11185
rect 10089 11159 10095 11185
rect 10121 11159 10127 11185
rect 12273 11159 12279 11185
rect 12305 11159 12311 11185
rect 7687 11153 7713 11159
rect 9367 11153 9393 11159
rect 10319 11153 10345 11159
rect 12559 11153 12585 11159
rect 12895 11185 12921 11191
rect 12895 11153 12921 11159
rect 13343 11185 13369 11191
rect 13343 11153 13369 11159
rect 13511 11185 13537 11191
rect 18825 11159 18831 11185
rect 18857 11159 18863 11185
rect 13511 11153 13537 11159
rect 8415 11129 8441 11135
rect 8415 11097 8441 11103
rect 9199 11129 9225 11135
rect 9199 11097 9225 11103
rect 10655 11129 10681 11135
rect 10655 11097 10681 11103
rect 10711 11129 10737 11135
rect 13231 11129 13257 11135
rect 11937 11103 11943 11129
rect 11969 11103 11975 11129
rect 10711 11097 10737 11103
rect 13231 11097 13257 11103
rect 7911 11073 7937 11079
rect 7911 11041 7937 11047
rect 8023 11073 8049 11079
rect 8023 11041 8049 11047
rect 8471 11073 8497 11079
rect 8863 11073 8889 11079
rect 8689 11047 8695 11073
rect 8721 11047 8727 11073
rect 8471 11041 8497 11047
rect 8863 11041 8889 11047
rect 9143 11073 9169 11079
rect 9703 11073 9729 11079
rect 9529 11047 9535 11073
rect 9561 11047 9567 11073
rect 9865 11047 9871 11073
rect 9897 11047 9903 11073
rect 9143 11041 9169 11047
rect 9703 11041 9729 11047
rect 672 10989 20328 11006
rect 672 10963 9919 10989
rect 9945 10963 9971 10989
rect 9997 10963 10023 10989
rect 10049 10963 20328 10989
rect 672 10946 20328 10963
rect 6399 10905 6425 10911
rect 6399 10873 6425 10879
rect 6791 10905 6817 10911
rect 6791 10873 6817 10879
rect 8135 10905 8161 10911
rect 8135 10873 8161 10879
rect 8247 10905 8273 10911
rect 8247 10873 8273 10879
rect 11943 10905 11969 10911
rect 11943 10873 11969 10879
rect 12335 10905 12361 10911
rect 12335 10873 12361 10879
rect 6511 10849 6537 10855
rect 6511 10817 6537 10823
rect 8807 10849 8833 10855
rect 8807 10817 8833 10823
rect 9535 10849 9561 10855
rect 9535 10817 9561 10823
rect 10263 10849 10289 10855
rect 10263 10817 10289 10823
rect 10319 10849 10345 10855
rect 11383 10849 11409 10855
rect 10817 10823 10823 10849
rect 10849 10823 10855 10849
rect 11545 10823 11551 10849
rect 11577 10823 11583 10849
rect 10319 10817 10345 10823
rect 11383 10817 11409 10823
rect 6567 10793 6593 10799
rect 2137 10767 2143 10793
rect 2169 10767 2175 10793
rect 6567 10761 6593 10767
rect 6847 10793 6873 10799
rect 6847 10761 6873 10767
rect 8303 10793 8329 10799
rect 8303 10761 8329 10767
rect 8919 10793 8945 10799
rect 8919 10761 8945 10767
rect 9031 10793 9057 10799
rect 10431 10793 10457 10799
rect 11271 10793 11297 10799
rect 11775 10793 11801 10799
rect 9137 10767 9143 10793
rect 9169 10767 9175 10793
rect 10033 10767 10039 10793
rect 10065 10767 10071 10793
rect 10705 10767 10711 10793
rect 10737 10767 10743 10793
rect 11489 10767 11495 10793
rect 11521 10767 11527 10793
rect 9031 10761 9057 10767
rect 10431 10761 10457 10767
rect 11271 10761 11297 10767
rect 11775 10761 11801 10767
rect 11943 10793 11969 10799
rect 11943 10761 11969 10767
rect 12055 10793 12081 10799
rect 12833 10767 12839 10793
rect 12865 10767 12871 10793
rect 18825 10767 18831 10793
rect 18857 10767 18863 10793
rect 12055 10761 12081 10767
rect 7071 10737 7097 10743
rect 9647 10737 9673 10743
rect 9081 10711 9087 10737
rect 9113 10711 9119 10737
rect 9473 10711 9479 10737
rect 9505 10711 9511 10737
rect 7071 10705 7097 10711
rect 9647 10705 9673 10711
rect 9815 10737 9841 10743
rect 20007 10737 20033 10743
rect 11657 10711 11663 10737
rect 11689 10711 11695 10737
rect 13169 10711 13175 10737
rect 13201 10711 13207 10737
rect 14233 10711 14239 10737
rect 14265 10711 14271 10737
rect 9815 10705 9841 10711
rect 20007 10705 20033 10711
rect 967 10681 993 10687
rect 967 10649 993 10655
rect 6791 10681 6817 10687
rect 6791 10649 6817 10655
rect 672 10597 20328 10614
rect 672 10571 2239 10597
rect 2265 10571 2291 10597
rect 2317 10571 2343 10597
rect 2369 10571 17599 10597
rect 17625 10571 17651 10597
rect 17677 10571 17703 10597
rect 17729 10571 20328 10597
rect 672 10554 20328 10571
rect 9535 10513 9561 10519
rect 9535 10481 9561 10487
rect 13007 10457 13033 10463
rect 1017 10431 1023 10457
rect 1049 10431 1055 10457
rect 4993 10431 4999 10457
rect 5025 10431 5031 10457
rect 6057 10431 6063 10457
rect 6089 10431 6095 10457
rect 8801 10431 8807 10457
rect 8833 10431 8839 10457
rect 12217 10431 12223 10457
rect 12249 10431 12255 10457
rect 13007 10425 13033 10431
rect 13455 10457 13481 10463
rect 13455 10425 13481 10431
rect 6959 10401 6985 10407
rect 10935 10401 10961 10407
rect 2137 10375 2143 10401
rect 2169 10375 2175 10401
rect 6449 10375 6455 10401
rect 6481 10375 6487 10401
rect 9473 10375 9479 10401
rect 9505 10375 9511 10401
rect 9977 10375 9983 10401
rect 10009 10375 10015 10401
rect 6959 10369 6985 10375
rect 10935 10369 10961 10375
rect 10991 10401 11017 10407
rect 10991 10369 11017 10375
rect 11271 10401 11297 10407
rect 11271 10369 11297 10375
rect 11551 10401 11577 10407
rect 11551 10369 11577 10375
rect 12895 10401 12921 10407
rect 12895 10369 12921 10375
rect 13119 10401 13145 10407
rect 13119 10369 13145 10375
rect 13175 10401 13201 10407
rect 13175 10369 13201 10375
rect 13343 10401 13369 10407
rect 13505 10375 13511 10401
rect 13537 10375 13543 10401
rect 13343 10369 13369 10375
rect 7239 10345 7265 10351
rect 7239 10313 7265 10319
rect 7463 10345 7489 10351
rect 9031 10345 9057 10351
rect 11047 10345 11073 10351
rect 8969 10319 8975 10345
rect 9001 10319 9007 10345
rect 9865 10319 9871 10345
rect 9897 10319 9903 10345
rect 10201 10319 10207 10345
rect 10233 10319 10239 10345
rect 7463 10313 7489 10319
rect 9031 10313 9057 10319
rect 11047 10313 11073 10319
rect 11607 10345 11633 10351
rect 11607 10313 11633 10319
rect 11663 10345 11689 10351
rect 12055 10345 12081 10351
rect 11713 10319 11719 10345
rect 11745 10319 11751 10345
rect 11663 10313 11689 10319
rect 12055 10313 12081 10319
rect 12167 10345 12193 10351
rect 12167 10313 12193 10319
rect 13623 10345 13649 10351
rect 13623 10313 13649 10319
rect 7015 10289 7041 10295
rect 7015 10257 7041 10263
rect 7071 10289 7097 10295
rect 7071 10257 7097 10263
rect 7127 10289 7153 10295
rect 7127 10257 7153 10263
rect 7407 10289 7433 10295
rect 7407 10257 7433 10263
rect 9087 10289 9113 10295
rect 9087 10257 9113 10263
rect 9199 10289 9225 10295
rect 9199 10257 9225 10263
rect 9591 10289 9617 10295
rect 9591 10257 9617 10263
rect 9703 10289 9729 10295
rect 9703 10257 9729 10263
rect 10375 10289 10401 10295
rect 10375 10257 10401 10263
rect 11383 10289 11409 10295
rect 11383 10257 11409 10263
rect 11495 10289 11521 10295
rect 11495 10257 11521 10263
rect 672 10205 20328 10222
rect 672 10179 9919 10205
rect 9945 10179 9971 10205
rect 9997 10179 10023 10205
rect 10049 10179 20328 10205
rect 672 10162 20328 10179
rect 7183 10121 7209 10127
rect 7183 10089 7209 10095
rect 8415 10065 8441 10071
rect 6561 10039 6567 10065
rect 6593 10039 6599 10065
rect 8241 10039 8247 10065
rect 8273 10039 8279 10065
rect 8415 10033 8441 10039
rect 9087 10065 9113 10071
rect 9087 10033 9113 10039
rect 9143 10065 9169 10071
rect 9143 10033 9169 10039
rect 8807 10009 8833 10015
rect 6953 9983 6959 10009
rect 6985 9983 6991 10009
rect 8969 9983 8975 10009
rect 9001 9983 9007 10009
rect 9305 9983 9311 10009
rect 9337 9983 9343 10009
rect 18825 9983 18831 10009
rect 18857 9983 18863 10009
rect 8807 9977 8833 9983
rect 12223 9953 12249 9959
rect 5497 9927 5503 9953
rect 5529 9927 5535 9953
rect 10313 9927 10319 9953
rect 10345 9927 10351 9953
rect 12223 9921 12249 9927
rect 20007 9897 20033 9903
rect 20007 9865 20033 9871
rect 672 9813 20328 9830
rect 672 9787 2239 9813
rect 2265 9787 2291 9813
rect 2317 9787 2343 9813
rect 2369 9787 17599 9813
rect 17625 9787 17651 9813
rect 17677 9787 17703 9813
rect 17729 9787 20328 9813
rect 672 9770 20328 9787
rect 11943 9729 11969 9735
rect 11943 9697 11969 9703
rect 8857 9647 8863 9673
rect 8889 9647 8895 9673
rect 13729 9647 13735 9673
rect 13761 9647 13767 9673
rect 7799 9617 7825 9623
rect 9087 9617 9113 9623
rect 8801 9591 8807 9617
rect 8833 9591 8839 9617
rect 7799 9585 7825 9591
rect 9087 9585 9113 9591
rect 9647 9617 9673 9623
rect 10369 9591 10375 9617
rect 10401 9591 10407 9617
rect 11601 9591 11607 9617
rect 11633 9591 11639 9617
rect 12273 9591 12279 9617
rect 12305 9591 12311 9617
rect 9647 9585 9673 9591
rect 8135 9561 8161 9567
rect 8135 9529 8161 9535
rect 8975 9561 9001 9567
rect 8975 9529 9001 9535
rect 9367 9561 9393 9567
rect 9367 9529 9393 9535
rect 9591 9561 9617 9567
rect 11775 9561 11801 9567
rect 9921 9535 9927 9561
rect 9953 9535 9959 9561
rect 10201 9535 10207 9561
rect 10233 9535 10239 9561
rect 11321 9535 11327 9561
rect 11353 9535 11359 9561
rect 11545 9535 11551 9561
rect 11577 9535 11583 9561
rect 9591 9529 9617 9535
rect 11775 9529 11801 9535
rect 11887 9561 11913 9567
rect 12665 9535 12671 9561
rect 12697 9535 12703 9561
rect 11887 9529 11913 9535
rect 7855 9505 7881 9511
rect 7855 9473 7881 9479
rect 7967 9505 7993 9511
rect 7967 9473 7993 9479
rect 8079 9505 8105 9511
rect 8079 9473 8105 9479
rect 9255 9505 9281 9511
rect 9255 9473 9281 9479
rect 9423 9505 9449 9511
rect 9423 9473 9449 9479
rect 9479 9505 9505 9511
rect 10033 9479 10039 9505
rect 10065 9479 10071 9505
rect 11097 9479 11103 9505
rect 11129 9479 11135 9505
rect 9479 9473 9505 9479
rect 672 9421 20328 9438
rect 672 9395 9919 9421
rect 9945 9395 9971 9421
rect 9997 9395 10023 9421
rect 10049 9395 20328 9421
rect 672 9378 20328 9395
rect 8191 9337 8217 9343
rect 8191 9305 8217 9311
rect 12055 9337 12081 9343
rect 12055 9305 12081 9311
rect 6617 9255 6623 9281
rect 6649 9255 6655 9281
rect 7625 9255 7631 9281
rect 7657 9255 7663 9281
rect 8857 9255 8863 9281
rect 8889 9255 8895 9281
rect 10425 9255 10431 9281
rect 10457 9255 10463 9281
rect 7463 9225 7489 9231
rect 8247 9225 8273 9231
rect 7009 9199 7015 9225
rect 7041 9199 7047 9225
rect 8129 9199 8135 9225
rect 8161 9199 8167 9225
rect 7463 9193 7489 9199
rect 8247 9193 8273 9199
rect 8695 9225 8721 9231
rect 8695 9193 8721 9199
rect 9255 9225 9281 9231
rect 9255 9193 9281 9199
rect 9871 9225 9897 9231
rect 9871 9193 9897 9199
rect 10151 9225 10177 9231
rect 10151 9193 10177 9199
rect 10263 9225 10289 9231
rect 11271 9225 11297 9231
rect 10593 9199 10599 9225
rect 10625 9199 10631 9225
rect 11153 9199 11159 9225
rect 11185 9199 11191 9225
rect 10263 9193 10289 9199
rect 11271 9193 11297 9199
rect 11943 9225 11969 9231
rect 11943 9193 11969 9199
rect 7239 9169 7265 9175
rect 5553 9143 5559 9169
rect 5585 9143 5591 9169
rect 7239 9137 7265 9143
rect 9143 9169 9169 9175
rect 10543 9169 10569 9175
rect 9417 9143 9423 9169
rect 9449 9143 9455 9169
rect 10089 9143 10095 9169
rect 10121 9143 10127 9169
rect 11489 9143 11495 9169
rect 11521 9143 11527 9169
rect 12105 9143 12111 9169
rect 12137 9143 12143 9169
rect 9143 9137 9169 9143
rect 10543 9137 10569 9143
rect 9983 9113 10009 9119
rect 9983 9081 10009 9087
rect 672 9029 20328 9046
rect 672 9003 2239 9029
rect 2265 9003 2291 9029
rect 2317 9003 2343 9029
rect 2369 9003 17599 9029
rect 17625 9003 17651 9029
rect 17677 9003 17703 9029
rect 17729 9003 20328 9029
rect 672 8986 20328 9003
rect 11999 8945 12025 8951
rect 11999 8913 12025 8919
rect 9927 8889 9953 8895
rect 6729 8863 6735 8889
rect 6761 8863 6767 8889
rect 7793 8863 7799 8889
rect 7825 8863 7831 8889
rect 9927 8857 9953 8863
rect 10711 8889 10737 8895
rect 10711 8857 10737 8863
rect 11887 8889 11913 8895
rect 20007 8889 20033 8895
rect 13673 8863 13679 8889
rect 13705 8863 13711 8889
rect 11887 8857 11913 8863
rect 20007 8857 20033 8863
rect 8527 8833 8553 8839
rect 9591 8833 9617 8839
rect 8185 8807 8191 8833
rect 8217 8807 8223 8833
rect 8913 8807 8919 8833
rect 8945 8807 8951 8833
rect 8527 8801 8553 8807
rect 9591 8801 9617 8807
rect 9759 8833 9785 8839
rect 9759 8801 9785 8807
rect 9871 8833 9897 8839
rect 10655 8833 10681 8839
rect 11831 8833 11857 8839
rect 10257 8807 10263 8833
rect 10289 8807 10295 8833
rect 10873 8807 10879 8833
rect 10905 8807 10911 8833
rect 11041 8807 11047 8833
rect 11073 8807 11079 8833
rect 11321 8807 11327 8833
rect 11353 8807 11359 8833
rect 12217 8807 12223 8833
rect 12249 8807 12255 8833
rect 13897 8807 13903 8833
rect 13929 8807 13935 8833
rect 18825 8807 18831 8833
rect 18857 8807 18863 8833
rect 9871 8801 9897 8807
rect 10655 8801 10681 8807
rect 11831 8801 11857 8807
rect 8695 8777 8721 8783
rect 8695 8745 8721 8751
rect 9647 8777 9673 8783
rect 9647 8745 9673 8751
rect 9983 8777 10009 8783
rect 9983 8745 10009 8751
rect 10039 8777 10065 8783
rect 10039 8745 10065 8751
rect 10767 8777 10793 8783
rect 10767 8745 10793 8751
rect 12055 8777 12081 8783
rect 12609 8751 12615 8777
rect 12641 8751 12647 8777
rect 12055 8745 12081 8751
rect 11607 8721 11633 8727
rect 9025 8695 9031 8721
rect 9057 8695 9063 8721
rect 11209 8695 11215 8721
rect 11241 8695 11247 8721
rect 14009 8695 14015 8721
rect 14041 8695 14047 8721
rect 11607 8689 11633 8695
rect 672 8637 20328 8654
rect 672 8611 9919 8637
rect 9945 8611 9971 8637
rect 9997 8611 10023 8637
rect 10049 8611 20328 8637
rect 672 8594 20328 8611
rect 7967 8553 7993 8559
rect 7967 8521 7993 8527
rect 9143 8497 9169 8503
rect 11601 8471 11607 8497
rect 11633 8471 11639 8497
rect 9143 8465 9169 8471
rect 7575 8441 7601 8447
rect 7401 8415 7407 8441
rect 7433 8415 7439 8441
rect 7575 8409 7601 8415
rect 7631 8441 7657 8447
rect 7631 8409 7657 8415
rect 7799 8441 7825 8447
rect 7799 8409 7825 8415
rect 8303 8441 8329 8447
rect 9809 8415 9815 8441
rect 9841 8415 9847 8441
rect 12777 8415 12783 8441
rect 12809 8415 12815 8441
rect 18937 8415 18943 8441
rect 18969 8415 18975 8441
rect 8303 8409 8329 8415
rect 12671 8385 12697 8391
rect 12671 8353 12697 8359
rect 20007 8385 20033 8391
rect 20007 8353 20033 8359
rect 9199 8329 9225 8335
rect 9199 8297 9225 8303
rect 12615 8329 12641 8335
rect 12615 8297 12641 8303
rect 672 8245 20328 8262
rect 672 8219 2239 8245
rect 2265 8219 2291 8245
rect 2317 8219 2343 8245
rect 2369 8219 17599 8245
rect 17625 8219 17651 8245
rect 17677 8219 17703 8245
rect 17729 8219 20328 8245
rect 672 8202 20328 8219
rect 12223 8161 12249 8167
rect 12223 8129 12249 8135
rect 967 8105 993 8111
rect 12559 8105 12585 8111
rect 12385 8079 12391 8105
rect 12417 8079 12423 8105
rect 967 8073 993 8079
rect 12559 8073 12585 8079
rect 6735 8049 6761 8055
rect 2137 8023 2143 8049
rect 2169 8023 2175 8049
rect 6735 8017 6761 8023
rect 9927 8049 9953 8055
rect 10705 8023 10711 8049
rect 10737 8023 10743 8049
rect 9927 8017 9953 8023
rect 9759 7993 9785 7999
rect 9759 7961 9785 7967
rect 9815 7993 9841 7999
rect 12671 7993 12697 7999
rect 10817 7967 10823 7993
rect 10849 7967 10855 7993
rect 9815 7961 9841 7967
rect 12671 7961 12697 7967
rect 6791 7937 6817 7943
rect 6791 7905 6817 7911
rect 6903 7937 6929 7943
rect 6903 7905 6929 7911
rect 12335 7937 12361 7943
rect 12335 7905 12361 7911
rect 12615 7937 12641 7943
rect 12615 7905 12641 7911
rect 672 7853 20328 7870
rect 672 7827 9919 7853
rect 9945 7827 9971 7853
rect 9997 7827 10023 7853
rect 10049 7827 20328 7853
rect 672 7810 20328 7827
rect 8191 7769 8217 7775
rect 8191 7737 8217 7743
rect 10431 7769 10457 7775
rect 10431 7737 10457 7743
rect 10655 7769 10681 7775
rect 10655 7737 10681 7743
rect 10767 7769 10793 7775
rect 10767 7737 10793 7743
rect 6847 7713 6873 7719
rect 6847 7681 6873 7687
rect 6903 7713 6929 7719
rect 6903 7681 6929 7687
rect 8023 7713 8049 7719
rect 9809 7687 9815 7713
rect 9841 7687 9847 7713
rect 8023 7681 8049 7687
rect 7015 7657 7041 7663
rect 6281 7631 6287 7657
rect 6313 7631 6319 7657
rect 6673 7631 6679 7657
rect 6705 7631 6711 7657
rect 7015 7625 7041 7631
rect 8191 7657 8217 7663
rect 8191 7625 8217 7631
rect 8303 7657 8329 7663
rect 8303 7625 8329 7631
rect 9087 7657 9113 7663
rect 9087 7625 9113 7631
rect 9311 7657 9337 7663
rect 9311 7625 9337 7631
rect 9423 7657 9449 7663
rect 9423 7625 9449 7631
rect 9647 7657 9673 7663
rect 9647 7625 9673 7631
rect 10319 7657 10345 7663
rect 10319 7625 10345 7631
rect 10487 7657 10513 7663
rect 10487 7625 10513 7631
rect 10991 7657 11017 7663
rect 10991 7625 11017 7631
rect 7183 7601 7209 7607
rect 5217 7575 5223 7601
rect 5249 7575 5255 7601
rect 7183 7569 7209 7575
rect 10711 7601 10737 7607
rect 10711 7569 10737 7575
rect 9031 7545 9057 7551
rect 9031 7513 9057 7519
rect 9087 7545 9113 7551
rect 9087 7513 9113 7519
rect 672 7461 20328 7478
rect 672 7435 2239 7461
rect 2265 7435 2291 7461
rect 2317 7435 2343 7461
rect 2369 7435 17599 7461
rect 17625 7435 17651 7461
rect 17677 7435 17703 7461
rect 17729 7435 20328 7461
rect 672 7418 20328 7435
rect 11159 7377 11185 7383
rect 11159 7345 11185 7351
rect 11663 7321 11689 7327
rect 9473 7295 9479 7321
rect 9505 7295 9511 7321
rect 12217 7295 12223 7321
rect 12249 7295 12255 7321
rect 13281 7295 13287 7321
rect 13313 7295 13319 7321
rect 11663 7289 11689 7295
rect 7687 7265 7713 7271
rect 9703 7265 9729 7271
rect 8073 7239 8079 7265
rect 8105 7239 8111 7265
rect 7687 7233 7713 7239
rect 9703 7233 9729 7239
rect 10431 7265 10457 7271
rect 10431 7233 10457 7239
rect 10599 7265 10625 7271
rect 10599 7233 10625 7239
rect 10823 7265 10849 7271
rect 10823 7233 10849 7239
rect 10935 7265 10961 7271
rect 11825 7239 11831 7265
rect 11857 7239 11863 7265
rect 10935 7233 10961 7239
rect 7631 7209 7657 7215
rect 10263 7209 10289 7215
rect 8409 7183 8415 7209
rect 8441 7183 8447 7209
rect 7631 7177 7657 7183
rect 10263 7177 10289 7183
rect 11103 7209 11129 7215
rect 11103 7177 11129 7183
rect 7519 7153 7545 7159
rect 7519 7121 7545 7127
rect 10319 7153 10345 7159
rect 10319 7121 10345 7127
rect 10879 7153 10905 7159
rect 10879 7121 10905 7127
rect 11159 7153 11185 7159
rect 11159 7121 11185 7127
rect 672 7069 20328 7086
rect 672 7043 9919 7069
rect 9945 7043 9971 7069
rect 9997 7043 10023 7069
rect 10049 7043 20328 7069
rect 672 7026 20328 7043
rect 8751 6985 8777 6991
rect 8751 6953 8777 6959
rect 9031 6985 9057 6991
rect 9031 6953 9057 6959
rect 11831 6985 11857 6991
rect 11831 6953 11857 6959
rect 9143 6929 9169 6935
rect 7233 6903 7239 6929
rect 7265 6903 7271 6929
rect 9143 6897 9169 6903
rect 9199 6929 9225 6935
rect 10537 6903 10543 6929
rect 10569 6903 10575 6929
rect 9199 6897 9225 6903
rect 6897 6847 6903 6873
rect 6929 6847 6935 6873
rect 10201 6847 10207 6873
rect 10233 6847 10239 6873
rect 8297 6791 8303 6817
rect 8329 6791 8335 6817
rect 11601 6791 11607 6817
rect 11633 6791 11639 6817
rect 672 6677 20328 6694
rect 672 6651 2239 6677
rect 2265 6651 2291 6677
rect 2317 6651 2343 6677
rect 2369 6651 17599 6677
rect 17625 6651 17651 6677
rect 17677 6651 17703 6677
rect 17729 6651 20328 6677
rect 672 6634 20328 6651
rect 672 6285 20328 6302
rect 672 6259 9919 6285
rect 9945 6259 9971 6285
rect 9997 6259 10023 6285
rect 10049 6259 20328 6285
rect 672 6242 20328 6259
rect 11439 6201 11465 6207
rect 11439 6169 11465 6175
rect 10817 6119 10823 6145
rect 10849 6119 10855 6145
rect 11209 6063 11215 6089
rect 11241 6063 11247 6089
rect 9753 6007 9759 6033
rect 9785 6007 9791 6033
rect 672 5893 20328 5910
rect 672 5867 2239 5893
rect 2265 5867 2291 5893
rect 2317 5867 2343 5893
rect 2369 5867 17599 5893
rect 17625 5867 17651 5893
rect 17677 5867 17703 5893
rect 17729 5867 20328 5893
rect 672 5850 20328 5867
rect 672 5501 20328 5518
rect 672 5475 9919 5501
rect 9945 5475 9971 5501
rect 9997 5475 10023 5501
rect 10049 5475 20328 5501
rect 672 5458 20328 5475
rect 672 5109 20328 5126
rect 672 5083 2239 5109
rect 2265 5083 2291 5109
rect 2317 5083 2343 5109
rect 2369 5083 17599 5109
rect 17625 5083 17651 5109
rect 17677 5083 17703 5109
rect 17729 5083 20328 5109
rect 672 5066 20328 5083
rect 672 4717 20328 4734
rect 672 4691 9919 4717
rect 9945 4691 9971 4717
rect 9997 4691 10023 4717
rect 10049 4691 20328 4717
rect 672 4674 20328 4691
rect 672 4325 20328 4342
rect 672 4299 2239 4325
rect 2265 4299 2291 4325
rect 2317 4299 2343 4325
rect 2369 4299 17599 4325
rect 17625 4299 17651 4325
rect 17677 4299 17703 4325
rect 17729 4299 20328 4325
rect 672 4282 20328 4299
rect 672 3933 20328 3950
rect 672 3907 9919 3933
rect 9945 3907 9971 3933
rect 9997 3907 10023 3933
rect 10049 3907 20328 3933
rect 672 3890 20328 3907
rect 672 3541 20328 3558
rect 672 3515 2239 3541
rect 2265 3515 2291 3541
rect 2317 3515 2343 3541
rect 2369 3515 17599 3541
rect 17625 3515 17651 3541
rect 17677 3515 17703 3541
rect 17729 3515 20328 3541
rect 672 3498 20328 3515
rect 672 3149 20328 3166
rect 672 3123 9919 3149
rect 9945 3123 9971 3149
rect 9997 3123 10023 3149
rect 10049 3123 20328 3149
rect 672 3106 20328 3123
rect 672 2757 20328 2774
rect 672 2731 2239 2757
rect 2265 2731 2291 2757
rect 2317 2731 2343 2757
rect 2369 2731 17599 2757
rect 17625 2731 17651 2757
rect 17677 2731 17703 2757
rect 17729 2731 20328 2757
rect 672 2714 20328 2731
rect 672 2365 20328 2382
rect 672 2339 9919 2365
rect 9945 2339 9971 2365
rect 9997 2339 10023 2365
rect 10049 2339 20328 2365
rect 672 2322 20328 2339
rect 9529 2143 9535 2169
rect 9561 2143 9567 2169
rect 12609 2143 12615 2169
rect 12641 2143 12647 2169
rect 10039 2057 10065 2063
rect 10039 2025 10065 2031
rect 13119 2057 13145 2063
rect 13119 2025 13145 2031
rect 672 1973 20328 1990
rect 672 1947 2239 1973
rect 2265 1947 2291 1973
rect 2317 1947 2343 1973
rect 2369 1947 17599 1973
rect 17625 1947 17651 1973
rect 17677 1947 17703 1973
rect 17729 1947 20328 1973
rect 672 1930 20328 1947
rect 12783 1833 12809 1839
rect 12783 1801 12809 1807
rect 8521 1751 8527 1777
rect 8553 1751 8559 1777
rect 10705 1751 10711 1777
rect 10737 1751 10743 1777
rect 12273 1751 12279 1777
rect 12305 1751 12311 1777
rect 9031 1665 9057 1671
rect 9031 1633 9057 1639
rect 11215 1665 11241 1671
rect 11215 1633 11241 1639
rect 672 1581 20328 1598
rect 672 1555 9919 1581
rect 9945 1555 9971 1581
rect 9997 1555 10023 1581
rect 10049 1555 20328 1581
rect 672 1538 20328 1555
<< via1 >>
rect 2239 19195 2265 19221
rect 2291 19195 2317 19221
rect 2343 19195 2369 19221
rect 17599 19195 17625 19221
rect 17651 19195 17677 19221
rect 17703 19195 17729 19221
rect 12783 19111 12809 19137
rect 9087 19055 9113 19081
rect 11103 19055 11129 19081
rect 9871 18999 9897 19025
rect 11999 18999 12025 19025
rect 12279 18999 12305 19025
rect 5839 18943 5865 18969
rect 17599 18943 17625 18969
rect 9919 18803 9945 18829
rect 9971 18803 9997 18829
rect 10023 18803 10049 18829
rect 11047 18719 11073 18745
rect 14071 18719 14097 18745
rect 10543 18607 10569 18633
rect 13567 18607 13593 18633
rect 2239 18411 2265 18437
rect 2291 18411 2317 18437
rect 2343 18411 2369 18437
rect 17599 18411 17625 18437
rect 17651 18411 17677 18437
rect 17703 18411 17729 18437
rect 11159 18327 11185 18353
rect 10655 18215 10681 18241
rect 855 18159 881 18185
rect 9919 18019 9945 18045
rect 9971 18019 9997 18045
rect 10023 18019 10049 18045
rect 2239 17627 2265 17653
rect 2291 17627 2317 17653
rect 2343 17627 2369 17653
rect 17599 17627 17625 17653
rect 17651 17627 17677 17653
rect 17703 17627 17729 17653
rect 9919 17235 9945 17261
rect 9971 17235 9997 17261
rect 10023 17235 10049 17261
rect 2239 16843 2265 16869
rect 2291 16843 2317 16869
rect 2343 16843 2369 16869
rect 17599 16843 17625 16869
rect 17651 16843 17677 16869
rect 17703 16843 17729 16869
rect 9919 16451 9945 16477
rect 9971 16451 9997 16477
rect 10023 16451 10049 16477
rect 2239 16059 2265 16085
rect 2291 16059 2317 16085
rect 2343 16059 2369 16085
rect 17599 16059 17625 16085
rect 17651 16059 17677 16085
rect 17703 16059 17729 16085
rect 9919 15667 9945 15693
rect 9971 15667 9997 15693
rect 10023 15667 10049 15693
rect 2239 15275 2265 15301
rect 2291 15275 2317 15301
rect 2343 15275 2369 15301
rect 17599 15275 17625 15301
rect 17651 15275 17677 15301
rect 17703 15275 17729 15301
rect 9919 14883 9945 14909
rect 9971 14883 9997 14909
rect 10023 14883 10049 14909
rect 2239 14491 2265 14517
rect 2291 14491 2317 14517
rect 2343 14491 2369 14517
rect 17599 14491 17625 14517
rect 17651 14491 17677 14517
rect 17703 14491 17729 14517
rect 10039 14295 10065 14321
rect 10151 14239 10177 14265
rect 10207 14239 10233 14265
rect 9919 14099 9945 14125
rect 9971 14099 9997 14125
rect 10023 14099 10049 14125
rect 9815 14015 9841 14041
rect 9983 14015 10009 14041
rect 12951 14015 12977 14041
rect 9255 13959 9281 13985
rect 9311 13959 9337 13985
rect 9143 13903 9169 13929
rect 10207 13903 10233 13929
rect 13007 13903 13033 13929
rect 10543 13847 10569 13873
rect 11607 13847 11633 13873
rect 11887 13847 11913 13873
rect 12951 13791 12977 13817
rect 2239 13707 2265 13733
rect 2291 13707 2317 13733
rect 2343 13707 2369 13733
rect 17599 13707 17625 13733
rect 17651 13707 17677 13733
rect 17703 13707 17729 13733
rect 8639 13567 8665 13593
rect 9199 13567 9225 13593
rect 10263 13567 10289 13593
rect 13455 13567 13481 13593
rect 20007 13567 20033 13593
rect 7183 13511 7209 13537
rect 8807 13511 8833 13537
rect 10655 13511 10681 13537
rect 11159 13511 11185 13537
rect 12055 13511 12081 13537
rect 18831 13511 18857 13537
rect 7575 13455 7601 13481
rect 10823 13455 10849 13481
rect 10991 13455 11017 13481
rect 11103 13455 11129 13481
rect 12391 13455 12417 13481
rect 10767 13399 10793 13425
rect 11831 13399 11857 13425
rect 9919 13315 9945 13341
rect 9971 13315 9997 13341
rect 10023 13315 10049 13341
rect 8975 13231 9001 13257
rect 9591 13231 9617 13257
rect 10375 13231 10401 13257
rect 9031 13175 9057 13201
rect 12279 13175 12305 13201
rect 12335 13175 12361 13201
rect 9143 13119 9169 13145
rect 9255 13119 9281 13145
rect 9367 13119 9393 13145
rect 9479 13119 9505 13145
rect 9647 13119 9673 13145
rect 10487 13119 10513 13145
rect 12615 13119 12641 13145
rect 8751 13063 8777 13089
rect 10767 13063 10793 13089
rect 12055 13063 12081 13089
rect 13007 13063 13033 13089
rect 14071 13063 14097 13089
rect 12279 13007 12305 13033
rect 2239 12923 2265 12949
rect 2291 12923 2317 12949
rect 2343 12923 2369 12949
rect 17599 12923 17625 12949
rect 17651 12923 17677 12949
rect 17703 12923 17729 12949
rect 12951 12839 12977 12865
rect 12111 12783 12137 12809
rect 12335 12783 12361 12809
rect 10655 12727 10681 12753
rect 13175 12727 13201 12753
rect 11047 12671 11073 12697
rect 13007 12671 13033 12697
rect 13231 12671 13257 12697
rect 12951 12615 12977 12641
rect 13343 12615 13369 12641
rect 9919 12531 9945 12557
rect 9971 12531 9997 12557
rect 10023 12531 10049 12557
rect 10823 12447 10849 12473
rect 7239 12391 7265 12417
rect 2143 12335 2169 12361
rect 7071 12335 7097 12361
rect 7407 12335 7433 12361
rect 10767 12335 10793 12361
rect 5615 12279 5641 12305
rect 6679 12279 6705 12305
rect 7631 12279 7657 12305
rect 967 12223 993 12249
rect 10823 12223 10849 12249
rect 2239 12139 2265 12165
rect 2291 12139 2317 12165
rect 2343 12139 2369 12165
rect 17599 12139 17625 12165
rect 17651 12139 17677 12165
rect 17703 12139 17729 12165
rect 11047 12055 11073 12081
rect 11103 12055 11129 12081
rect 9367 11999 9393 12025
rect 9927 11999 9953 12025
rect 20007 11999 20033 12025
rect 6679 11943 6705 11969
rect 7127 11943 7153 11969
rect 7967 11943 7993 11969
rect 10711 11943 10737 11969
rect 10823 11943 10849 11969
rect 11047 11943 11073 11969
rect 18831 11943 18857 11969
rect 6847 11887 6873 11913
rect 8303 11887 8329 11913
rect 9535 11887 9561 11913
rect 9703 11887 9729 11913
rect 13455 11887 13481 11913
rect 13511 11887 13537 11913
rect 6791 11831 6817 11857
rect 6959 11831 6985 11857
rect 7071 11831 7097 11857
rect 13343 11831 13369 11857
rect 9919 11747 9945 11773
rect 9971 11747 9997 11773
rect 10023 11747 10049 11773
rect 8751 11663 8777 11689
rect 9311 11607 9337 11633
rect 10935 11607 10961 11633
rect 14631 11607 14657 11633
rect 6735 11551 6761 11577
rect 8359 11551 8385 11577
rect 8695 11551 8721 11577
rect 8807 11551 8833 11577
rect 9031 11551 9057 11577
rect 9143 11551 9169 11577
rect 9759 11551 9785 11577
rect 12839 11551 12865 11577
rect 14519 11551 14545 11577
rect 18831 11551 18857 11577
rect 7071 11495 7097 11521
rect 8135 11495 8161 11521
rect 12671 11495 12697 11521
rect 13231 11495 13257 11521
rect 14295 11495 14321 11521
rect 8415 11439 8441 11465
rect 20007 11439 20033 11465
rect 2239 11355 2265 11381
rect 2291 11355 2317 11381
rect 2343 11355 2369 11381
rect 17599 11355 17625 11381
rect 17651 11355 17677 11381
rect 17703 11355 17729 11381
rect 8471 11271 8497 11297
rect 7967 11215 7993 11241
rect 8247 11215 8273 11241
rect 10879 11215 10905 11241
rect 12783 11215 12809 11241
rect 13063 11215 13089 11241
rect 13455 11215 13481 11241
rect 20007 11215 20033 11241
rect 7687 11159 7713 11185
rect 9031 11159 9057 11185
rect 9367 11159 9393 11185
rect 10095 11159 10121 11185
rect 10319 11159 10345 11185
rect 12279 11159 12305 11185
rect 12559 11159 12585 11185
rect 12895 11159 12921 11185
rect 13343 11159 13369 11185
rect 13511 11159 13537 11185
rect 18831 11159 18857 11185
rect 8415 11103 8441 11129
rect 9199 11103 9225 11129
rect 10655 11103 10681 11129
rect 10711 11103 10737 11129
rect 11943 11103 11969 11129
rect 13231 11103 13257 11129
rect 7911 11047 7937 11073
rect 8023 11047 8049 11073
rect 8471 11047 8497 11073
rect 8695 11047 8721 11073
rect 8863 11047 8889 11073
rect 9143 11047 9169 11073
rect 9535 11047 9561 11073
rect 9703 11047 9729 11073
rect 9871 11047 9897 11073
rect 9919 10963 9945 10989
rect 9971 10963 9997 10989
rect 10023 10963 10049 10989
rect 6399 10879 6425 10905
rect 6791 10879 6817 10905
rect 8135 10879 8161 10905
rect 8247 10879 8273 10905
rect 11943 10879 11969 10905
rect 12335 10879 12361 10905
rect 6511 10823 6537 10849
rect 8807 10823 8833 10849
rect 9535 10823 9561 10849
rect 10263 10823 10289 10849
rect 10319 10823 10345 10849
rect 10823 10823 10849 10849
rect 11383 10823 11409 10849
rect 11551 10823 11577 10849
rect 2143 10767 2169 10793
rect 6567 10767 6593 10793
rect 6847 10767 6873 10793
rect 8303 10767 8329 10793
rect 8919 10767 8945 10793
rect 9031 10767 9057 10793
rect 9143 10767 9169 10793
rect 10039 10767 10065 10793
rect 10431 10767 10457 10793
rect 10711 10767 10737 10793
rect 11271 10767 11297 10793
rect 11495 10767 11521 10793
rect 11775 10767 11801 10793
rect 11943 10767 11969 10793
rect 12055 10767 12081 10793
rect 12839 10767 12865 10793
rect 18831 10767 18857 10793
rect 7071 10711 7097 10737
rect 9087 10711 9113 10737
rect 9479 10711 9505 10737
rect 9647 10711 9673 10737
rect 9815 10711 9841 10737
rect 11663 10711 11689 10737
rect 13175 10711 13201 10737
rect 14239 10711 14265 10737
rect 20007 10711 20033 10737
rect 967 10655 993 10681
rect 6791 10655 6817 10681
rect 2239 10571 2265 10597
rect 2291 10571 2317 10597
rect 2343 10571 2369 10597
rect 17599 10571 17625 10597
rect 17651 10571 17677 10597
rect 17703 10571 17729 10597
rect 9535 10487 9561 10513
rect 1023 10431 1049 10457
rect 4999 10431 5025 10457
rect 6063 10431 6089 10457
rect 8807 10431 8833 10457
rect 12223 10431 12249 10457
rect 13007 10431 13033 10457
rect 13455 10431 13481 10457
rect 2143 10375 2169 10401
rect 6455 10375 6481 10401
rect 6959 10375 6985 10401
rect 9479 10375 9505 10401
rect 9983 10375 10009 10401
rect 10935 10375 10961 10401
rect 10991 10375 11017 10401
rect 11271 10375 11297 10401
rect 11551 10375 11577 10401
rect 12895 10375 12921 10401
rect 13119 10375 13145 10401
rect 13175 10375 13201 10401
rect 13343 10375 13369 10401
rect 13511 10375 13537 10401
rect 7239 10319 7265 10345
rect 7463 10319 7489 10345
rect 8975 10319 9001 10345
rect 9031 10319 9057 10345
rect 9871 10319 9897 10345
rect 10207 10319 10233 10345
rect 11047 10319 11073 10345
rect 11607 10319 11633 10345
rect 11663 10319 11689 10345
rect 11719 10319 11745 10345
rect 12055 10319 12081 10345
rect 12167 10319 12193 10345
rect 13623 10319 13649 10345
rect 7015 10263 7041 10289
rect 7071 10263 7097 10289
rect 7127 10263 7153 10289
rect 7407 10263 7433 10289
rect 9087 10263 9113 10289
rect 9199 10263 9225 10289
rect 9591 10263 9617 10289
rect 9703 10263 9729 10289
rect 10375 10263 10401 10289
rect 11383 10263 11409 10289
rect 11495 10263 11521 10289
rect 9919 10179 9945 10205
rect 9971 10179 9997 10205
rect 10023 10179 10049 10205
rect 7183 10095 7209 10121
rect 6567 10039 6593 10065
rect 8247 10039 8273 10065
rect 8415 10039 8441 10065
rect 9087 10039 9113 10065
rect 9143 10039 9169 10065
rect 6959 9983 6985 10009
rect 8807 9983 8833 10009
rect 8975 9983 9001 10009
rect 9311 9983 9337 10009
rect 18831 9983 18857 10009
rect 5503 9927 5529 9953
rect 10319 9927 10345 9953
rect 12223 9927 12249 9953
rect 20007 9871 20033 9897
rect 2239 9787 2265 9813
rect 2291 9787 2317 9813
rect 2343 9787 2369 9813
rect 17599 9787 17625 9813
rect 17651 9787 17677 9813
rect 17703 9787 17729 9813
rect 11943 9703 11969 9729
rect 8863 9647 8889 9673
rect 13735 9647 13761 9673
rect 7799 9591 7825 9617
rect 8807 9591 8833 9617
rect 9087 9591 9113 9617
rect 9647 9591 9673 9617
rect 10375 9591 10401 9617
rect 11607 9591 11633 9617
rect 12279 9591 12305 9617
rect 8135 9535 8161 9561
rect 8975 9535 9001 9561
rect 9367 9535 9393 9561
rect 9591 9535 9617 9561
rect 9927 9535 9953 9561
rect 10207 9535 10233 9561
rect 11327 9535 11353 9561
rect 11551 9535 11577 9561
rect 11775 9535 11801 9561
rect 11887 9535 11913 9561
rect 12671 9535 12697 9561
rect 7855 9479 7881 9505
rect 7967 9479 7993 9505
rect 8079 9479 8105 9505
rect 9255 9479 9281 9505
rect 9423 9479 9449 9505
rect 9479 9479 9505 9505
rect 10039 9479 10065 9505
rect 11103 9479 11129 9505
rect 9919 9395 9945 9421
rect 9971 9395 9997 9421
rect 10023 9395 10049 9421
rect 8191 9311 8217 9337
rect 12055 9311 12081 9337
rect 6623 9255 6649 9281
rect 7631 9255 7657 9281
rect 8863 9255 8889 9281
rect 10431 9255 10457 9281
rect 7015 9199 7041 9225
rect 7463 9199 7489 9225
rect 8135 9199 8161 9225
rect 8247 9199 8273 9225
rect 8695 9199 8721 9225
rect 9255 9199 9281 9225
rect 9871 9199 9897 9225
rect 10151 9199 10177 9225
rect 10263 9199 10289 9225
rect 10599 9199 10625 9225
rect 11159 9199 11185 9225
rect 11271 9199 11297 9225
rect 11943 9199 11969 9225
rect 5559 9143 5585 9169
rect 7239 9143 7265 9169
rect 9143 9143 9169 9169
rect 9423 9143 9449 9169
rect 10095 9143 10121 9169
rect 10543 9143 10569 9169
rect 11495 9143 11521 9169
rect 12111 9143 12137 9169
rect 9983 9087 10009 9113
rect 2239 9003 2265 9029
rect 2291 9003 2317 9029
rect 2343 9003 2369 9029
rect 17599 9003 17625 9029
rect 17651 9003 17677 9029
rect 17703 9003 17729 9029
rect 11999 8919 12025 8945
rect 6735 8863 6761 8889
rect 7799 8863 7825 8889
rect 9927 8863 9953 8889
rect 10711 8863 10737 8889
rect 11887 8863 11913 8889
rect 13679 8863 13705 8889
rect 20007 8863 20033 8889
rect 8191 8807 8217 8833
rect 8527 8807 8553 8833
rect 8919 8807 8945 8833
rect 9591 8807 9617 8833
rect 9759 8807 9785 8833
rect 9871 8807 9897 8833
rect 10263 8807 10289 8833
rect 10655 8807 10681 8833
rect 10879 8807 10905 8833
rect 11047 8807 11073 8833
rect 11327 8807 11353 8833
rect 11831 8807 11857 8833
rect 12223 8807 12249 8833
rect 13903 8807 13929 8833
rect 18831 8807 18857 8833
rect 8695 8751 8721 8777
rect 9647 8751 9673 8777
rect 9983 8751 10009 8777
rect 10039 8751 10065 8777
rect 10767 8751 10793 8777
rect 12055 8751 12081 8777
rect 12615 8751 12641 8777
rect 9031 8695 9057 8721
rect 11215 8695 11241 8721
rect 11607 8695 11633 8721
rect 14015 8695 14041 8721
rect 9919 8611 9945 8637
rect 9971 8611 9997 8637
rect 10023 8611 10049 8637
rect 7967 8527 7993 8553
rect 9143 8471 9169 8497
rect 11607 8471 11633 8497
rect 7407 8415 7433 8441
rect 7575 8415 7601 8441
rect 7631 8415 7657 8441
rect 7799 8415 7825 8441
rect 8303 8415 8329 8441
rect 9815 8415 9841 8441
rect 12783 8415 12809 8441
rect 18943 8415 18969 8441
rect 12671 8359 12697 8385
rect 20007 8359 20033 8385
rect 9199 8303 9225 8329
rect 12615 8303 12641 8329
rect 2239 8219 2265 8245
rect 2291 8219 2317 8245
rect 2343 8219 2369 8245
rect 17599 8219 17625 8245
rect 17651 8219 17677 8245
rect 17703 8219 17729 8245
rect 12223 8135 12249 8161
rect 967 8079 993 8105
rect 12391 8079 12417 8105
rect 12559 8079 12585 8105
rect 2143 8023 2169 8049
rect 6735 8023 6761 8049
rect 9927 8023 9953 8049
rect 10711 8023 10737 8049
rect 9759 7967 9785 7993
rect 9815 7967 9841 7993
rect 10823 7967 10849 7993
rect 12671 7967 12697 7993
rect 6791 7911 6817 7937
rect 6903 7911 6929 7937
rect 12335 7911 12361 7937
rect 12615 7911 12641 7937
rect 9919 7827 9945 7853
rect 9971 7827 9997 7853
rect 10023 7827 10049 7853
rect 8191 7743 8217 7769
rect 10431 7743 10457 7769
rect 10655 7743 10681 7769
rect 10767 7743 10793 7769
rect 6847 7687 6873 7713
rect 6903 7687 6929 7713
rect 8023 7687 8049 7713
rect 9815 7687 9841 7713
rect 6287 7631 6313 7657
rect 6679 7631 6705 7657
rect 7015 7631 7041 7657
rect 8191 7631 8217 7657
rect 8303 7631 8329 7657
rect 9087 7631 9113 7657
rect 9311 7631 9337 7657
rect 9423 7631 9449 7657
rect 9647 7631 9673 7657
rect 10319 7631 10345 7657
rect 10487 7631 10513 7657
rect 10991 7631 11017 7657
rect 5223 7575 5249 7601
rect 7183 7575 7209 7601
rect 10711 7575 10737 7601
rect 9031 7519 9057 7545
rect 9087 7519 9113 7545
rect 2239 7435 2265 7461
rect 2291 7435 2317 7461
rect 2343 7435 2369 7461
rect 17599 7435 17625 7461
rect 17651 7435 17677 7461
rect 17703 7435 17729 7461
rect 11159 7351 11185 7377
rect 9479 7295 9505 7321
rect 11663 7295 11689 7321
rect 12223 7295 12249 7321
rect 13287 7295 13313 7321
rect 7687 7239 7713 7265
rect 8079 7239 8105 7265
rect 9703 7239 9729 7265
rect 10431 7239 10457 7265
rect 10599 7239 10625 7265
rect 10823 7239 10849 7265
rect 10935 7239 10961 7265
rect 11831 7239 11857 7265
rect 7631 7183 7657 7209
rect 8415 7183 8441 7209
rect 10263 7183 10289 7209
rect 11103 7183 11129 7209
rect 7519 7127 7545 7153
rect 10319 7127 10345 7153
rect 10879 7127 10905 7153
rect 11159 7127 11185 7153
rect 9919 7043 9945 7069
rect 9971 7043 9997 7069
rect 10023 7043 10049 7069
rect 8751 6959 8777 6985
rect 9031 6959 9057 6985
rect 11831 6959 11857 6985
rect 7239 6903 7265 6929
rect 9143 6903 9169 6929
rect 9199 6903 9225 6929
rect 10543 6903 10569 6929
rect 6903 6847 6929 6873
rect 10207 6847 10233 6873
rect 8303 6791 8329 6817
rect 11607 6791 11633 6817
rect 2239 6651 2265 6677
rect 2291 6651 2317 6677
rect 2343 6651 2369 6677
rect 17599 6651 17625 6677
rect 17651 6651 17677 6677
rect 17703 6651 17729 6677
rect 9919 6259 9945 6285
rect 9971 6259 9997 6285
rect 10023 6259 10049 6285
rect 11439 6175 11465 6201
rect 10823 6119 10849 6145
rect 11215 6063 11241 6089
rect 9759 6007 9785 6033
rect 2239 5867 2265 5893
rect 2291 5867 2317 5893
rect 2343 5867 2369 5893
rect 17599 5867 17625 5893
rect 17651 5867 17677 5893
rect 17703 5867 17729 5893
rect 9919 5475 9945 5501
rect 9971 5475 9997 5501
rect 10023 5475 10049 5501
rect 2239 5083 2265 5109
rect 2291 5083 2317 5109
rect 2343 5083 2369 5109
rect 17599 5083 17625 5109
rect 17651 5083 17677 5109
rect 17703 5083 17729 5109
rect 9919 4691 9945 4717
rect 9971 4691 9997 4717
rect 10023 4691 10049 4717
rect 2239 4299 2265 4325
rect 2291 4299 2317 4325
rect 2343 4299 2369 4325
rect 17599 4299 17625 4325
rect 17651 4299 17677 4325
rect 17703 4299 17729 4325
rect 9919 3907 9945 3933
rect 9971 3907 9997 3933
rect 10023 3907 10049 3933
rect 2239 3515 2265 3541
rect 2291 3515 2317 3541
rect 2343 3515 2369 3541
rect 17599 3515 17625 3541
rect 17651 3515 17677 3541
rect 17703 3515 17729 3541
rect 9919 3123 9945 3149
rect 9971 3123 9997 3149
rect 10023 3123 10049 3149
rect 2239 2731 2265 2757
rect 2291 2731 2317 2757
rect 2343 2731 2369 2757
rect 17599 2731 17625 2757
rect 17651 2731 17677 2757
rect 17703 2731 17729 2757
rect 9919 2339 9945 2365
rect 9971 2339 9997 2365
rect 10023 2339 10049 2365
rect 9535 2143 9561 2169
rect 12615 2143 12641 2169
rect 10039 2031 10065 2057
rect 13119 2031 13145 2057
rect 2239 1947 2265 1973
rect 2291 1947 2317 1973
rect 2343 1947 2369 1973
rect 17599 1947 17625 1973
rect 17651 1947 17677 1973
rect 17703 1947 17729 1973
rect 12783 1807 12809 1833
rect 8527 1751 8553 1777
rect 10711 1751 10737 1777
rect 12279 1751 12305 1777
rect 9031 1639 9057 1665
rect 11215 1639 11241 1665
rect 9919 1555 9945 1581
rect 9971 1555 9997 1581
rect 10023 1555 10049 1581
<< metal2 >>
rect 5712 20600 5768 21000
rect 9072 20600 9128 21000
rect 10080 20600 10136 21000
rect 10416 20600 10472 21000
rect 11088 20600 11144 21000
rect 11424 20600 11480 21000
rect 13440 20600 13496 21000
rect 17472 20600 17528 21000
rect 2238 19222 2370 19227
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2238 19189 2370 19194
rect 5726 18970 5754 20600
rect 9086 19081 9114 20600
rect 9086 19055 9087 19081
rect 9113 19055 9114 19081
rect 9086 19049 9114 19055
rect 9870 19026 9898 19031
rect 9590 19025 9898 19026
rect 9590 18999 9871 19025
rect 9897 18999 9898 19025
rect 9590 18998 9898 18999
rect 5838 18970 5866 18975
rect 5726 18969 5866 18970
rect 5726 18943 5839 18969
rect 5865 18943 5866 18969
rect 5726 18942 5866 18943
rect 5838 18937 5866 18942
rect 2238 18438 2370 18443
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2238 18405 2370 18410
rect 854 18186 882 18191
rect 854 18139 882 18158
rect 2238 17654 2370 17659
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2238 17621 2370 17626
rect 2238 16870 2370 16875
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2238 16837 2370 16842
rect 2238 16086 2370 16091
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2238 16053 2370 16058
rect 2238 15302 2370 15307
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2238 15269 2370 15274
rect 2238 14518 2370 14523
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2238 14485 2370 14490
rect 9310 14322 9338 14327
rect 9254 13985 9282 13991
rect 9254 13959 9255 13985
rect 9281 13959 9282 13985
rect 9142 13930 9170 13935
rect 9142 13929 9226 13930
rect 9142 13903 9143 13929
rect 9169 13903 9226 13929
rect 9142 13902 9226 13903
rect 9142 13897 9170 13902
rect 2086 13818 2114 13823
rect 966 12250 994 12255
rect 966 12203 994 12222
rect 966 10681 994 10687
rect 966 10655 967 10681
rect 993 10655 994 10681
rect 966 10458 994 10655
rect 966 10425 994 10430
rect 1022 10457 1050 10463
rect 1022 10431 1023 10457
rect 1049 10431 1050 10457
rect 1022 10122 1050 10431
rect 1022 10089 1050 10094
rect 2086 9954 2114 13790
rect 2238 13734 2370 13739
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2238 13701 2370 13706
rect 8638 13594 8666 13599
rect 8638 13547 8666 13566
rect 9198 13593 9226 13902
rect 9198 13567 9199 13593
rect 9225 13567 9226 13593
rect 9198 13561 9226 13567
rect 7182 13537 7210 13543
rect 8806 13538 8834 13543
rect 7182 13511 7183 13537
rect 7209 13511 7210 13537
rect 2238 12950 2370 12955
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2238 12917 2370 12922
rect 2142 12362 2170 12367
rect 2142 12315 2170 12334
rect 5614 12362 5642 12367
rect 5614 12305 5642 12334
rect 6958 12362 6986 12367
rect 7070 12362 7098 12367
rect 7182 12362 7210 13511
rect 8750 13537 8834 13538
rect 8750 13511 8807 13537
rect 8833 13511 8834 13537
rect 8750 13510 8834 13511
rect 7574 13481 7602 13487
rect 7574 13455 7575 13481
rect 7601 13455 7602 13481
rect 7574 13258 7602 13455
rect 7574 13225 7602 13230
rect 8750 13089 8778 13510
rect 8806 13505 8834 13510
rect 9254 13454 9282 13959
rect 9310 13985 9338 14294
rect 9310 13959 9311 13985
rect 9337 13959 9338 13985
rect 9310 13953 9338 13959
rect 9590 13594 9618 18998
rect 9870 18993 9898 18998
rect 9918 18830 10050 18835
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 9918 18797 10050 18802
rect 10094 18354 10122 20600
rect 10430 18746 10458 20600
rect 11102 19081 11130 20600
rect 11438 19138 11466 20600
rect 11438 19105 11466 19110
rect 12782 19138 12810 19143
rect 12782 19091 12810 19110
rect 11102 19055 11103 19081
rect 11129 19055 11130 19081
rect 11102 19049 11130 19055
rect 11998 19025 12026 19031
rect 11998 18999 11999 19025
rect 12025 18999 12026 19025
rect 10430 18713 10458 18718
rect 11046 18746 11074 18751
rect 11046 18699 11074 18718
rect 10094 18321 10122 18326
rect 10542 18633 10570 18639
rect 10542 18607 10543 18633
rect 10569 18607 10570 18633
rect 10150 18242 10178 18247
rect 9918 18046 10050 18051
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 9918 18013 10050 18018
rect 9918 17262 10050 17267
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 9918 17229 10050 17234
rect 9918 16478 10050 16483
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 9918 16445 10050 16450
rect 9918 15694 10050 15699
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 9918 15661 10050 15666
rect 9918 14910 10050 14915
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 9918 14877 10050 14882
rect 10038 14322 10066 14327
rect 10038 14275 10066 14294
rect 9870 14266 9898 14271
rect 9814 14238 9870 14266
rect 9814 14041 9842 14238
rect 9870 14233 9898 14238
rect 10150 14266 10178 18214
rect 10150 14154 10178 14238
rect 10206 14265 10234 14271
rect 10206 14239 10207 14265
rect 10233 14239 10234 14265
rect 10206 14210 10234 14239
rect 10206 14182 10346 14210
rect 9918 14126 10050 14131
rect 10150 14126 10290 14154
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 9918 14093 10050 14098
rect 9814 14015 9815 14041
rect 9841 14015 9842 14041
rect 9814 14009 9842 14015
rect 9982 14042 10010 14047
rect 9982 13995 10010 14014
rect 9254 13426 9338 13454
rect 8974 13258 9002 13263
rect 8974 13211 9002 13230
rect 9030 13202 9058 13207
rect 9030 13155 9058 13174
rect 8750 13063 8751 13089
rect 8777 13063 8778 13089
rect 6986 12334 7042 12362
rect 6958 12329 6986 12334
rect 5614 12279 5615 12305
rect 5641 12279 5642 12305
rect 5614 12273 5642 12279
rect 6678 12305 6706 12311
rect 6678 12279 6679 12305
rect 6705 12279 6706 12305
rect 2238 12166 2370 12171
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2238 12133 2370 12138
rect 6678 11969 6706 12279
rect 6678 11943 6679 11969
rect 6705 11943 6706 11969
rect 6678 11937 6706 11943
rect 6734 11970 6762 11975
rect 6734 11577 6762 11942
rect 6846 11914 6874 11919
rect 6846 11867 6874 11886
rect 6790 11857 6818 11863
rect 6790 11831 6791 11857
rect 6817 11831 6818 11857
rect 6790 11802 6818 11831
rect 6958 11857 6986 11863
rect 6958 11831 6959 11857
rect 6985 11831 6986 11857
rect 6958 11802 6986 11831
rect 7014 11858 7042 12334
rect 7070 12361 7210 12362
rect 7070 12335 7071 12361
rect 7097 12335 7210 12361
rect 7070 12334 7210 12335
rect 7238 12417 7266 12423
rect 7238 12391 7239 12417
rect 7265 12391 7266 12417
rect 7070 12306 7098 12334
rect 7070 11970 7098 12278
rect 7238 12026 7266 12391
rect 7406 12362 7434 12367
rect 7406 12315 7434 12334
rect 7630 12306 7658 12311
rect 7630 12259 7658 12278
rect 7966 12306 7994 12311
rect 7070 11937 7098 11942
rect 7126 11998 7266 12026
rect 7126 11969 7154 11998
rect 7126 11943 7127 11969
rect 7153 11943 7154 11969
rect 7070 11858 7098 11863
rect 7014 11857 7098 11858
rect 7014 11831 7071 11857
rect 7097 11831 7098 11857
rect 7014 11830 7098 11831
rect 7070 11825 7098 11830
rect 6790 11774 6986 11802
rect 6734 11551 6735 11577
rect 6761 11551 6762 11577
rect 2238 11382 2370 11387
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2238 11349 2370 11354
rect 6398 10906 6426 10911
rect 6398 10859 6426 10878
rect 4998 10850 5026 10855
rect 2142 10794 2170 10799
rect 2142 10747 2170 10766
rect 2238 10598 2370 10603
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2238 10565 2370 10570
rect 4998 10457 5026 10822
rect 6510 10850 6538 10855
rect 6510 10803 6538 10822
rect 6566 10794 6594 10799
rect 6566 10747 6594 10766
rect 4998 10431 4999 10457
rect 5025 10431 5026 10457
rect 4998 10425 5026 10431
rect 6062 10682 6090 10687
rect 6062 10457 6090 10654
rect 6062 10431 6063 10457
rect 6089 10431 6090 10457
rect 6062 10425 6090 10431
rect 2142 10402 2170 10407
rect 2142 10355 2170 10374
rect 6454 10402 6482 10407
rect 6454 10355 6482 10374
rect 6734 10402 6762 11551
rect 7070 11522 7098 11527
rect 7070 11475 7098 11494
rect 6790 10906 6818 10911
rect 6790 10859 6818 10878
rect 6846 10793 6874 10799
rect 6846 10767 6847 10793
rect 6873 10767 6874 10793
rect 6790 10682 6818 10687
rect 6790 10635 6818 10654
rect 6846 10514 6874 10767
rect 6846 10481 6874 10486
rect 6958 10794 6986 10799
rect 6958 10402 6986 10766
rect 7126 10794 7154 11943
rect 7966 11970 7994 12278
rect 8750 12306 8778 13063
rect 8750 12273 8778 12278
rect 9142 13145 9170 13151
rect 9142 13119 9143 13145
rect 9169 13119 9170 13145
rect 8470 12026 8498 12031
rect 7966 11969 8218 11970
rect 7966 11943 7967 11969
rect 7993 11943 8218 11969
rect 7966 11942 8218 11943
rect 7966 11937 7994 11942
rect 7686 11746 7714 11751
rect 7686 11186 7714 11718
rect 8134 11578 8162 11583
rect 7966 11522 7994 11527
rect 7966 11241 7994 11494
rect 8134 11521 8162 11550
rect 8134 11495 8135 11521
rect 8161 11495 8162 11521
rect 8134 11489 8162 11495
rect 7966 11215 7967 11241
rect 7993 11215 7994 11241
rect 7966 11209 7994 11215
rect 8190 11242 8218 11942
rect 8302 11913 8330 11919
rect 8302 11887 8303 11913
rect 8329 11887 8330 11913
rect 8302 11690 8330 11887
rect 8302 11657 8330 11662
rect 8358 11578 8386 11583
rect 8358 11531 8386 11550
rect 8414 11466 8442 11471
rect 8414 11419 8442 11438
rect 8470 11297 8498 11998
rect 9030 12026 9058 12031
rect 8750 11690 8778 11695
rect 8750 11643 8778 11662
rect 8694 11578 8722 11583
rect 8470 11271 8471 11297
rect 8497 11271 8498 11297
rect 8470 11265 8498 11271
rect 8638 11577 8722 11578
rect 8638 11551 8695 11577
rect 8721 11551 8722 11577
rect 8638 11550 8722 11551
rect 8246 11242 8274 11247
rect 8190 11241 8274 11242
rect 8190 11215 8247 11241
rect 8273 11215 8274 11241
rect 8190 11214 8274 11215
rect 8246 11209 8274 11214
rect 7686 11139 7714 11158
rect 8134 11186 8162 11191
rect 7910 11074 7938 11079
rect 7910 11027 7938 11046
rect 8022 11073 8050 11079
rect 8022 11047 8023 11073
rect 8049 11047 8050 11073
rect 8022 11018 8050 11047
rect 8022 10985 8050 10990
rect 8134 10905 8162 11158
rect 8414 11129 8442 11135
rect 8414 11103 8415 11129
rect 8441 11103 8442 11129
rect 8134 10879 8135 10905
rect 8161 10879 8162 10905
rect 8134 10873 8162 10879
rect 8246 11074 8274 11079
rect 8246 10905 8274 11046
rect 8246 10879 8247 10905
rect 8273 10879 8274 10905
rect 8246 10873 8274 10879
rect 7126 10761 7154 10766
rect 8302 10794 8330 10799
rect 8302 10747 8330 10766
rect 6734 10369 6762 10374
rect 6846 10401 6986 10402
rect 6846 10375 6959 10401
rect 6985 10375 6986 10401
rect 6846 10374 6986 10375
rect 2086 9921 2114 9926
rect 5502 10234 5530 10239
rect 5502 9953 5530 10206
rect 6566 10122 6594 10127
rect 6566 10065 6594 10094
rect 6566 10039 6567 10065
rect 6593 10039 6594 10065
rect 6566 10033 6594 10039
rect 5502 9927 5503 9953
rect 5529 9927 5530 9953
rect 5502 9921 5530 9927
rect 2238 9814 2370 9819
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2238 9781 2370 9786
rect 6622 9282 6650 9287
rect 6622 9235 6650 9254
rect 5558 9170 5586 9175
rect 5558 9123 5586 9142
rect 2238 9030 2370 9035
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2238 8997 2370 9002
rect 6734 8890 6762 8895
rect 6734 8843 6762 8862
rect 2238 8246 2370 8251
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2238 8213 2370 8218
rect 966 8105 994 8111
rect 966 8079 967 8105
rect 993 8079 994 8105
rect 966 7770 994 8079
rect 2142 8050 2170 8055
rect 2142 8003 2170 8022
rect 5222 8050 5250 8055
rect 966 7737 994 7742
rect 5222 7938 5250 8022
rect 6734 8050 6762 8055
rect 6846 8050 6874 10374
rect 6958 10369 6986 10374
rect 7070 10737 7098 10743
rect 7070 10711 7071 10737
rect 7097 10711 7098 10737
rect 7070 10402 7098 10711
rect 7098 10374 7210 10402
rect 7070 10369 7098 10374
rect 6958 10290 6986 10295
rect 6958 10009 6986 10262
rect 7014 10289 7042 10295
rect 7014 10263 7015 10289
rect 7041 10263 7042 10289
rect 7014 10234 7042 10263
rect 7070 10290 7098 10295
rect 7070 10243 7098 10262
rect 7126 10289 7154 10295
rect 7126 10263 7127 10289
rect 7153 10263 7154 10289
rect 7014 10201 7042 10206
rect 7126 10178 7154 10263
rect 7126 10145 7154 10150
rect 7182 10121 7210 10374
rect 7182 10095 7183 10121
rect 7209 10095 7210 10121
rect 7182 10089 7210 10095
rect 7238 10345 7266 10351
rect 7238 10319 7239 10345
rect 7265 10319 7266 10345
rect 6958 9983 6959 10009
rect 6985 9983 6986 10009
rect 6958 9977 6986 9983
rect 7238 9618 7266 10319
rect 7462 10345 7490 10351
rect 7462 10319 7463 10345
rect 7489 10319 7490 10345
rect 7406 10289 7434 10295
rect 7406 10263 7407 10289
rect 7433 10263 7434 10289
rect 7406 10122 7434 10263
rect 7462 10290 7490 10319
rect 7462 10257 7490 10262
rect 7406 10089 7434 10094
rect 7798 10178 7826 10183
rect 8414 10178 8442 11103
rect 8470 11074 8498 11079
rect 8638 11074 8666 11550
rect 8694 11545 8722 11550
rect 8806 11577 8834 11583
rect 8806 11551 8807 11577
rect 8833 11551 8834 11577
rect 8806 11242 8834 11551
rect 9030 11577 9058 11998
rect 9142 11858 9170 13119
rect 9254 13145 9282 13151
rect 9254 13119 9255 13145
rect 9281 13119 9282 13145
rect 9198 11858 9226 11863
rect 9142 11830 9198 11858
rect 9198 11825 9226 11830
rect 9254 11746 9282 13119
rect 9310 12026 9338 13426
rect 9590 13257 9618 13566
rect 10206 13929 10234 13935
rect 10206 13903 10207 13929
rect 10233 13903 10234 13929
rect 10206 13454 10234 13903
rect 10262 13593 10290 14126
rect 10262 13567 10263 13593
rect 10289 13567 10290 13593
rect 10262 13561 10290 13567
rect 10318 13538 10346 14182
rect 10542 14042 10570 18607
rect 11158 18354 11186 18359
rect 11158 18307 11186 18326
rect 10654 18242 10682 18247
rect 10654 18195 10682 18214
rect 11998 15974 12026 18999
rect 12278 19025 12306 19031
rect 12278 18999 12279 19025
rect 12305 18999 12306 19025
rect 11998 15946 12138 15974
rect 10542 14009 10570 14014
rect 10542 13874 10570 13879
rect 11102 13874 11130 13879
rect 10542 13873 10682 13874
rect 10542 13847 10543 13873
rect 10569 13847 10682 13873
rect 10542 13846 10682 13847
rect 10542 13841 10570 13846
rect 10374 13538 10402 13543
rect 10318 13510 10374 13538
rect 10094 13426 10234 13454
rect 9918 13342 10050 13347
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 9918 13309 10050 13314
rect 9590 13231 9591 13257
rect 9617 13231 9618 13257
rect 9590 13225 9618 13231
rect 9366 13146 9394 13151
rect 9478 13146 9506 13151
rect 9366 13145 9506 13146
rect 9366 13119 9367 13145
rect 9393 13119 9479 13145
rect 9505 13119 9506 13145
rect 9366 13118 9506 13119
rect 9366 13113 9394 13118
rect 9478 13113 9506 13118
rect 9646 13145 9674 13151
rect 9646 13119 9647 13145
rect 9673 13119 9674 13145
rect 9646 12362 9674 13119
rect 10094 12754 10122 13426
rect 10374 13257 10402 13510
rect 10654 13537 10682 13846
rect 10654 13511 10655 13537
rect 10681 13511 10682 13537
rect 10654 13505 10682 13511
rect 10822 13482 10850 13487
rect 10990 13482 11018 13487
rect 10822 13481 11018 13482
rect 10822 13455 10823 13481
rect 10849 13455 10991 13481
rect 11017 13455 11018 13481
rect 10822 13454 11018 13455
rect 10822 13449 10850 13454
rect 10990 13449 11018 13454
rect 11102 13481 11130 13846
rect 11606 13874 11634 13879
rect 11606 13827 11634 13846
rect 11886 13873 11914 13879
rect 11886 13847 11887 13873
rect 11913 13847 11914 13873
rect 11158 13538 11186 13543
rect 11158 13491 11186 13510
rect 11102 13455 11103 13481
rect 11129 13455 11130 13481
rect 11102 13449 11130 13455
rect 11886 13454 11914 13847
rect 10374 13231 10375 13257
rect 10401 13231 10402 13257
rect 10374 13225 10402 13231
rect 10766 13425 10794 13431
rect 10766 13399 10767 13425
rect 10793 13399 10794 13425
rect 10766 13202 10794 13399
rect 11830 13426 11914 13454
rect 12054 13537 12082 13543
rect 12054 13511 12055 13537
rect 12081 13511 12082 13537
rect 11830 13425 11858 13426
rect 11830 13399 11831 13425
rect 11857 13399 11858 13425
rect 10794 13174 10906 13202
rect 10766 13169 10794 13174
rect 9918 12558 10050 12563
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 9918 12525 10050 12530
rect 10094 12474 10122 12726
rect 10038 12446 10122 12474
rect 10486 13145 10514 13151
rect 10486 13119 10487 13145
rect 10513 13119 10514 13145
rect 9702 12362 9730 12367
rect 9646 12334 9702 12362
rect 9310 11993 9338 11998
rect 9366 12026 9394 12031
rect 9366 12025 9450 12026
rect 9366 11999 9367 12025
rect 9393 11999 9450 12025
rect 9366 11998 9450 11999
rect 9366 11993 9394 11998
rect 9030 11551 9031 11577
rect 9057 11551 9058 11577
rect 9030 11545 9058 11551
rect 9086 11718 9282 11746
rect 8806 11209 8834 11214
rect 9030 11466 9058 11471
rect 9030 11186 9058 11438
rect 9030 11139 9058 11158
rect 8470 11073 8666 11074
rect 8470 11047 8471 11073
rect 8497 11047 8666 11073
rect 8470 11046 8666 11047
rect 8694 11074 8722 11079
rect 8722 11046 8834 11074
rect 8470 11018 8498 11046
rect 8694 11027 8722 11046
rect 8470 10738 8498 10990
rect 8806 10906 8834 11046
rect 8862 11073 8890 11079
rect 8862 11047 8863 11073
rect 8889 11047 8890 11073
rect 8862 11018 8890 11047
rect 8862 10985 8890 10990
rect 8806 10878 9002 10906
rect 8806 10849 8834 10878
rect 8806 10823 8807 10849
rect 8833 10823 8834 10849
rect 8806 10817 8834 10823
rect 8470 10705 8498 10710
rect 8862 10794 8890 10799
rect 8918 10794 8946 10799
rect 8890 10793 8946 10794
rect 8890 10767 8919 10793
rect 8945 10767 8946 10793
rect 8890 10766 8946 10767
rect 8806 10514 8834 10519
rect 8806 10457 8834 10486
rect 8806 10431 8807 10457
rect 8833 10431 8834 10457
rect 8806 10425 8834 10431
rect 7238 9585 7266 9590
rect 7798 9618 7826 10150
rect 8358 10150 8442 10178
rect 8246 10066 8274 10071
rect 8358 10066 8386 10150
rect 8246 10065 8386 10066
rect 8246 10039 8247 10065
rect 8273 10039 8386 10065
rect 8246 10038 8386 10039
rect 8414 10066 8442 10071
rect 8246 9730 8274 10038
rect 8414 10019 8442 10038
rect 8806 10010 8834 10015
rect 8806 9963 8834 9982
rect 8078 9702 8274 9730
rect 8078 9618 8106 9702
rect 7798 9617 8106 9618
rect 7798 9591 7799 9617
rect 7825 9591 8106 9617
rect 7798 9590 8106 9591
rect 8806 9674 8834 9679
rect 8806 9617 8834 9646
rect 8862 9673 8890 10766
rect 8918 10761 8946 10766
rect 8918 10346 8946 10351
rect 8918 10234 8946 10318
rect 8974 10345 9002 10878
rect 9030 10793 9058 10799
rect 9030 10767 9031 10793
rect 9057 10767 9058 10793
rect 9030 10458 9058 10767
rect 9086 10737 9114 11718
rect 9310 11633 9338 11639
rect 9310 11607 9311 11633
rect 9337 11607 9338 11633
rect 9142 11578 9170 11583
rect 9142 11531 9170 11550
rect 9254 11298 9282 11303
rect 9198 11130 9226 11135
rect 9198 11083 9226 11102
rect 9142 11073 9170 11079
rect 9142 11047 9143 11073
rect 9169 11047 9170 11073
rect 9142 10962 9170 11047
rect 9254 10962 9282 11270
rect 9142 10934 9282 10962
rect 9142 10794 9170 10799
rect 9142 10747 9170 10766
rect 9086 10711 9087 10737
rect 9113 10711 9114 10737
rect 9086 10705 9114 10711
rect 9030 10425 9058 10430
rect 9142 10682 9170 10687
rect 8974 10319 8975 10345
rect 9001 10319 9002 10345
rect 8974 10313 9002 10319
rect 9030 10345 9058 10351
rect 9030 10319 9031 10345
rect 9057 10319 9058 10345
rect 9030 10290 9058 10319
rect 9030 10257 9058 10262
rect 9086 10289 9114 10295
rect 9086 10263 9087 10289
rect 9113 10263 9114 10289
rect 8918 10206 9002 10234
rect 8862 9647 8863 9673
rect 8889 9647 8890 9673
rect 8862 9641 8890 9647
rect 8918 10122 8946 10127
rect 8806 9591 8807 9617
rect 8833 9591 8834 9617
rect 7798 9585 7826 9590
rect 7854 9505 7882 9511
rect 7854 9479 7855 9505
rect 7881 9479 7882 9505
rect 7630 9281 7658 9287
rect 7630 9255 7631 9281
rect 7657 9255 7658 9281
rect 7014 9225 7042 9231
rect 7014 9199 7015 9225
rect 7041 9199 7042 9225
rect 7014 9170 7042 9199
rect 7462 9225 7490 9231
rect 7462 9199 7463 9225
rect 7489 9199 7490 9225
rect 7238 9170 7266 9175
rect 7462 9170 7490 9199
rect 7014 9169 7266 9170
rect 7014 9143 7239 9169
rect 7265 9143 7266 9169
rect 7014 9142 7266 9143
rect 6734 8049 6874 8050
rect 6734 8023 6735 8049
rect 6761 8023 6874 8049
rect 6734 8022 6874 8023
rect 6734 8017 6762 8022
rect 5222 7601 5250 7910
rect 6790 7938 6818 7943
rect 6902 7938 6930 7943
rect 6790 7891 6818 7910
rect 6846 7937 6930 7938
rect 6846 7911 6903 7937
rect 6929 7911 6930 7937
rect 6846 7910 6930 7911
rect 6846 7713 6874 7910
rect 6902 7905 6930 7910
rect 6846 7687 6847 7713
rect 6873 7687 6874 7713
rect 6846 7681 6874 7687
rect 6902 7714 6930 7719
rect 6902 7667 6930 7686
rect 6286 7658 6314 7663
rect 6286 7611 6314 7630
rect 6678 7658 6706 7663
rect 7014 7658 7042 7663
rect 6678 7657 6762 7658
rect 6678 7631 6679 7657
rect 6705 7631 6762 7657
rect 6678 7630 6762 7631
rect 6678 7625 6706 7630
rect 5222 7575 5223 7601
rect 5249 7575 5250 7601
rect 5222 7569 5250 7575
rect 2238 7462 2370 7467
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2238 7429 2370 7434
rect 6734 7266 6762 7630
rect 7014 7611 7042 7630
rect 7182 7602 7210 7607
rect 7238 7602 7266 9142
rect 7406 9142 7462 9170
rect 7406 8441 7434 9142
rect 7462 9137 7490 9142
rect 7630 9170 7658 9255
rect 7630 9137 7658 9142
rect 7406 8415 7407 8441
rect 7433 8415 7434 8441
rect 7406 8409 7434 8415
rect 7574 8890 7602 8895
rect 7574 8441 7602 8862
rect 7798 8890 7826 8895
rect 7854 8890 7882 9479
rect 7966 9506 7994 9511
rect 7966 9459 7994 9478
rect 7798 8889 7994 8890
rect 7798 8863 7799 8889
rect 7825 8863 7994 8889
rect 7798 8862 7994 8863
rect 7798 8857 7826 8862
rect 7966 8553 7994 8862
rect 7966 8527 7967 8553
rect 7993 8527 7994 8553
rect 7966 8521 7994 8527
rect 7574 8415 7575 8441
rect 7601 8415 7602 8441
rect 7574 8409 7602 8415
rect 7630 8442 7658 8447
rect 7798 8442 7826 8447
rect 7630 8441 7826 8442
rect 7630 8415 7631 8441
rect 7657 8415 7799 8441
rect 7825 8415 7826 8441
rect 7630 8414 7826 8415
rect 7630 8409 7658 8414
rect 7798 8409 7826 8414
rect 8022 7713 8050 9590
rect 8806 9585 8834 9591
rect 8134 9561 8162 9567
rect 8134 9535 8135 9561
rect 8161 9535 8162 9561
rect 8078 9506 8106 9511
rect 8078 9282 8106 9478
rect 8078 9249 8106 9254
rect 8134 9225 8162 9535
rect 8190 9337 8218 9343
rect 8190 9311 8191 9337
rect 8217 9311 8218 9337
rect 8190 9282 8218 9311
rect 8190 9249 8218 9254
rect 8862 9282 8890 9287
rect 8918 9282 8946 10094
rect 8974 10009 9002 10206
rect 9086 10178 9114 10263
rect 9030 10150 9114 10178
rect 9030 10122 9058 10150
rect 9030 10089 9058 10094
rect 8974 9983 8975 10009
rect 9001 9983 9002 10009
rect 8974 9977 9002 9983
rect 9086 10066 9114 10071
rect 9086 9617 9114 10038
rect 9142 10065 9170 10654
rect 9142 10039 9143 10065
rect 9169 10039 9170 10065
rect 9142 10033 9170 10039
rect 9198 10289 9226 10295
rect 9198 10263 9199 10289
rect 9225 10263 9226 10289
rect 9086 9591 9087 9617
rect 9113 9591 9114 9617
rect 9086 9585 9114 9591
rect 8974 9561 9002 9567
rect 8974 9535 8975 9561
rect 9001 9535 9002 9561
rect 8974 9506 9002 9535
rect 8974 9473 9002 9478
rect 8862 9281 8946 9282
rect 8862 9255 8863 9281
rect 8889 9255 8946 9281
rect 8862 9254 8946 9255
rect 8134 9199 8135 9225
rect 8161 9199 8162 9225
rect 8134 9170 8162 9199
rect 8246 9226 8274 9231
rect 8246 9179 8274 9198
rect 8526 9226 8554 9231
rect 8134 9137 8162 9142
rect 8526 8890 8554 9198
rect 8694 9226 8722 9231
rect 8694 9179 8722 9198
rect 8862 9114 8890 9254
rect 8862 9081 8890 9086
rect 9086 9170 9114 9175
rect 9142 9170 9170 9175
rect 9114 9169 9170 9170
rect 9114 9143 9143 9169
rect 9169 9143 9170 9169
rect 9114 9142 9170 9143
rect 8190 8833 8218 8839
rect 8190 8807 8191 8833
rect 8217 8807 8218 8833
rect 8190 8442 8218 8807
rect 8526 8833 8554 8862
rect 8526 8807 8527 8833
rect 8553 8807 8554 8833
rect 8526 8801 8554 8807
rect 8694 8834 8722 8839
rect 8694 8777 8722 8806
rect 8918 8834 8946 8839
rect 9086 8834 9114 9142
rect 9142 9137 9170 9142
rect 9198 8946 9226 10263
rect 9254 9898 9282 10934
rect 9310 10346 9338 11607
rect 9366 11186 9394 11191
rect 9366 11139 9394 11158
rect 9422 11074 9450 11998
rect 9534 11913 9562 11919
rect 9534 11887 9535 11913
rect 9561 11887 9562 11913
rect 9534 11298 9562 11887
rect 9702 11913 9730 12334
rect 9702 11887 9703 11913
rect 9729 11887 9730 11913
rect 9702 11881 9730 11887
rect 9926 12306 9954 12311
rect 10038 12306 10066 12446
rect 10486 12362 10514 13119
rect 10766 13090 10794 13095
rect 10654 12754 10682 12759
rect 10766 12754 10794 13062
rect 10682 12726 10794 12754
rect 10654 12707 10682 12726
rect 10822 12474 10850 12479
rect 10822 12427 10850 12446
rect 10486 12329 10514 12334
rect 10766 12362 10794 12367
rect 10766 12315 10794 12334
rect 9954 12278 10066 12306
rect 9926 12025 9954 12278
rect 10822 12250 10850 12255
rect 10878 12250 10906 13174
rect 11830 13090 11858 13399
rect 11830 13057 11858 13062
rect 12054 13090 12082 13511
rect 12054 12810 12082 13062
rect 12054 12777 12082 12782
rect 12110 12809 12138 15946
rect 12278 13874 12306 18999
rect 13454 18746 13482 20600
rect 17486 18970 17514 20600
rect 17598 19222 17730 19227
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17598 19189 17730 19194
rect 17598 18970 17626 18975
rect 17486 18969 17626 18970
rect 17486 18943 17599 18969
rect 17625 18943 17626 18969
rect 17486 18942 17626 18943
rect 17598 18937 17626 18942
rect 13454 18713 13482 18718
rect 14070 18746 14098 18751
rect 14070 18699 14098 18718
rect 13566 18633 13594 18639
rect 13566 18607 13567 18633
rect 13593 18607 13594 18633
rect 13566 15974 13594 18607
rect 17598 18438 17730 18443
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17598 18405 17730 18410
rect 17598 17654 17730 17659
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17598 17621 17730 17626
rect 17598 16870 17730 16875
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17598 16837 17730 16842
rect 17598 16086 17730 16091
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17598 16053 17730 16058
rect 13454 15946 13594 15974
rect 12950 14042 12978 14047
rect 12950 13995 12978 14014
rect 13454 14042 13482 15946
rect 17598 15302 17730 15307
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17598 15269 17730 15274
rect 17598 14518 17730 14523
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17598 14485 17730 14490
rect 13006 13930 13034 13935
rect 13006 13929 13090 13930
rect 13006 13903 13007 13929
rect 13033 13903 13090 13929
rect 13006 13902 13090 13903
rect 13006 13897 13034 13902
rect 12278 13841 12306 13846
rect 12334 13818 12362 13823
rect 12278 13202 12306 13207
rect 12110 12783 12111 12809
rect 12137 12783 12138 12809
rect 11046 12697 11074 12703
rect 11046 12671 11047 12697
rect 11073 12671 11074 12697
rect 10878 12222 11018 12250
rect 10822 12203 10850 12222
rect 9926 11999 9927 12025
rect 9953 11999 9954 12025
rect 9926 11858 9954 11999
rect 10710 11970 10738 11975
rect 10822 11970 10850 11975
rect 10710 11969 10794 11970
rect 10710 11943 10711 11969
rect 10737 11943 10794 11969
rect 10710 11942 10794 11943
rect 10710 11937 10738 11942
rect 9926 11825 9954 11830
rect 9918 11774 10050 11779
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 9918 11741 10050 11746
rect 9646 11690 9674 11695
rect 9534 11265 9562 11270
rect 9590 11662 9646 11690
rect 9478 11074 9506 11079
rect 9422 11046 9478 11074
rect 9478 11041 9506 11046
rect 9534 11073 9562 11079
rect 9534 11047 9535 11073
rect 9561 11047 9562 11073
rect 9534 11018 9562 11047
rect 9534 10849 9562 10990
rect 9534 10823 9535 10849
rect 9561 10823 9562 10849
rect 9478 10794 9506 10799
rect 9478 10737 9506 10766
rect 9478 10711 9479 10737
rect 9505 10711 9506 10737
rect 9310 10313 9338 10318
rect 9366 10458 9394 10463
rect 9366 10122 9394 10430
rect 9478 10401 9506 10711
rect 9534 10626 9562 10823
rect 9590 10794 9618 11662
rect 9646 11657 9674 11662
rect 9758 11577 9786 11583
rect 9758 11551 9759 11577
rect 9785 11551 9786 11577
rect 9702 11074 9730 11079
rect 9590 10761 9618 10766
rect 9646 10906 9674 10911
rect 9646 10737 9674 10878
rect 9646 10711 9647 10737
rect 9673 10711 9674 10737
rect 9646 10705 9674 10711
rect 9702 10682 9730 11046
rect 9702 10649 9730 10654
rect 9534 10598 9618 10626
rect 9534 10514 9562 10519
rect 9534 10467 9562 10486
rect 9590 10402 9618 10598
rect 9478 10375 9479 10401
rect 9505 10375 9506 10401
rect 9478 10369 9506 10375
rect 9534 10374 9618 10402
rect 9646 10514 9674 10519
rect 9310 10010 9338 10015
rect 9310 9963 9338 9982
rect 9254 9870 9338 9898
rect 9198 8913 9226 8918
rect 9254 9505 9282 9511
rect 9254 9479 9255 9505
rect 9281 9479 9282 9505
rect 9254 9225 9282 9479
rect 9310 9450 9338 9870
rect 9366 9562 9394 10094
rect 9366 9515 9394 9534
rect 9422 10290 9450 10295
rect 9422 9505 9450 10262
rect 9534 9562 9562 10374
rect 9590 10289 9618 10295
rect 9590 10263 9591 10289
rect 9617 10263 9618 10289
rect 9590 10178 9618 10263
rect 9590 10145 9618 10150
rect 9646 9617 9674 10486
rect 9702 10289 9730 10295
rect 9702 10263 9703 10289
rect 9729 10263 9730 10289
rect 9702 10122 9730 10263
rect 9702 10089 9730 10094
rect 9758 9954 9786 11551
rect 10094 11185 10122 11191
rect 10094 11159 10095 11185
rect 10121 11159 10122 11185
rect 10094 11130 10122 11159
rect 10318 11186 10346 11191
rect 10318 11139 10346 11158
rect 10654 11130 10682 11135
rect 10122 11102 10290 11130
rect 10094 11097 10122 11102
rect 9870 11074 9898 11079
rect 9814 11073 9898 11074
rect 9814 11047 9871 11073
rect 9897 11047 9898 11073
rect 9814 11046 9898 11047
rect 9814 10906 9842 11046
rect 9870 11041 9898 11046
rect 9918 10990 10050 10995
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 9918 10957 10050 10962
rect 9870 10906 9898 10911
rect 9814 10878 9870 10906
rect 9870 10873 9898 10878
rect 10262 10849 10290 11102
rect 10654 11083 10682 11102
rect 10710 11129 10738 11135
rect 10710 11103 10711 11129
rect 10737 11103 10738 11129
rect 10710 11074 10738 11103
rect 10710 11041 10738 11046
rect 10262 10823 10263 10849
rect 10289 10823 10290 10849
rect 10262 10817 10290 10823
rect 10318 10850 10346 10855
rect 10318 10803 10346 10822
rect 10710 10850 10738 10855
rect 9870 10794 9898 10799
rect 9814 10737 9842 10743
rect 9814 10711 9815 10737
rect 9841 10711 9842 10737
rect 9814 10514 9842 10711
rect 9814 10481 9842 10486
rect 9870 10346 9898 10766
rect 10038 10793 10066 10799
rect 10038 10767 10039 10793
rect 10065 10767 10066 10793
rect 10038 10682 10066 10767
rect 10038 10649 10066 10654
rect 10206 10794 10234 10799
rect 9814 10345 9898 10346
rect 9814 10319 9871 10345
rect 9897 10319 9898 10345
rect 9814 10318 9898 10319
rect 9814 10234 9842 10318
rect 9870 10313 9898 10318
rect 9982 10401 10010 10407
rect 9982 10375 9983 10401
rect 10009 10375 10010 10401
rect 9926 10290 9954 10295
rect 9982 10290 10010 10375
rect 10206 10345 10234 10766
rect 10430 10793 10458 10799
rect 10430 10767 10431 10793
rect 10457 10767 10458 10793
rect 10430 10402 10458 10767
rect 10430 10369 10458 10374
rect 10710 10793 10738 10822
rect 10710 10767 10711 10793
rect 10737 10767 10738 10793
rect 10206 10319 10207 10345
rect 10233 10319 10234 10345
rect 10206 10313 10234 10319
rect 10710 10346 10738 10767
rect 9954 10262 10010 10290
rect 10374 10290 10402 10295
rect 9926 10257 9954 10262
rect 10374 10243 10402 10262
rect 10542 10290 10570 10295
rect 9814 10201 9842 10206
rect 9918 10206 10050 10211
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 9918 10173 10050 10178
rect 10038 10122 10066 10127
rect 9814 9954 9842 9959
rect 9758 9926 9814 9954
rect 9646 9591 9647 9617
rect 9673 9591 9674 9617
rect 9590 9562 9618 9567
rect 9534 9534 9590 9562
rect 9590 9515 9618 9534
rect 9422 9479 9423 9505
rect 9449 9479 9450 9505
rect 9310 9422 9394 9450
rect 9254 9199 9255 9225
rect 9281 9199 9282 9225
rect 9254 8834 9282 9199
rect 8918 8833 9114 8834
rect 8918 8807 8919 8833
rect 8945 8807 9114 8833
rect 8918 8806 9114 8807
rect 9142 8806 9254 8834
rect 8918 8801 8946 8806
rect 8694 8751 8695 8777
rect 8721 8751 8722 8777
rect 8694 8745 8722 8751
rect 9030 8722 9058 8727
rect 8302 8442 8330 8447
rect 8190 8441 8386 8442
rect 8190 8415 8303 8441
rect 8329 8415 8386 8441
rect 8190 8414 8386 8415
rect 8302 8409 8330 8414
rect 8190 7770 8218 7775
rect 8022 7687 8023 7713
rect 8049 7687 8050 7713
rect 8022 7681 8050 7687
rect 8078 7769 8218 7770
rect 8078 7743 8191 7769
rect 8217 7743 8218 7769
rect 8078 7742 8218 7743
rect 7182 7601 7266 7602
rect 7182 7575 7183 7601
rect 7209 7575 7266 7601
rect 7182 7574 7266 7575
rect 7630 7602 7658 7607
rect 6902 7266 6930 7271
rect 6734 7238 6902 7266
rect 6902 6873 6930 7238
rect 7182 7266 7210 7574
rect 7182 7233 7210 7238
rect 7630 7209 7658 7574
rect 8078 7434 8106 7742
rect 8190 7737 8218 7742
rect 7686 7406 8106 7434
rect 8190 7657 8218 7663
rect 8190 7631 8191 7657
rect 8217 7631 8218 7657
rect 7686 7265 7714 7406
rect 7686 7239 7687 7265
rect 7713 7239 7714 7265
rect 7686 7233 7714 7239
rect 8078 7266 8106 7271
rect 8078 7219 8106 7238
rect 7630 7183 7631 7209
rect 7657 7183 7658 7209
rect 7630 7177 7658 7183
rect 7518 7154 7546 7159
rect 7238 7153 7546 7154
rect 7238 7127 7519 7153
rect 7545 7127 7546 7153
rect 7238 7126 7546 7127
rect 7238 6929 7266 7126
rect 7518 7121 7546 7126
rect 7238 6903 7239 6929
rect 7265 6903 7266 6929
rect 7238 6897 7266 6903
rect 6902 6847 6903 6873
rect 6929 6847 6930 6873
rect 6902 6841 6930 6847
rect 8190 6818 8218 7631
rect 8302 7658 8330 7663
rect 8302 7611 8330 7630
rect 8302 7266 8330 7271
rect 8358 7266 8386 8414
rect 9030 7658 9058 8694
rect 9142 8497 9170 8806
rect 9254 8801 9282 8806
rect 9142 8471 9143 8497
rect 9169 8471 9170 8497
rect 9142 8465 9170 8471
rect 9198 8330 9226 8335
rect 9198 8329 9338 8330
rect 9198 8303 9199 8329
rect 9225 8303 9338 8329
rect 9198 8302 9338 8303
rect 9198 8297 9226 8302
rect 9310 7994 9338 8302
rect 9086 7658 9114 7663
rect 9030 7657 9114 7658
rect 9030 7631 9087 7657
rect 9113 7631 9114 7657
rect 9030 7630 9114 7631
rect 9086 7625 9114 7630
rect 9254 7658 9282 7663
rect 9030 7545 9058 7551
rect 9030 7519 9031 7545
rect 9057 7519 9058 7545
rect 8330 7238 8386 7266
rect 8750 7266 8778 7271
rect 8302 7233 8330 7238
rect 8414 7210 8442 7215
rect 8414 7163 8442 7182
rect 8750 6985 8778 7238
rect 8750 6959 8751 6985
rect 8777 6959 8778 6985
rect 8750 6953 8778 6959
rect 9030 6985 9058 7519
rect 9086 7545 9114 7551
rect 9086 7519 9087 7545
rect 9113 7519 9114 7545
rect 9086 7210 9114 7519
rect 9086 7177 9114 7182
rect 9030 6959 9031 6985
rect 9057 6959 9058 6985
rect 9030 6953 9058 6959
rect 9142 6930 9170 6935
rect 9142 6883 9170 6902
rect 9198 6930 9226 6935
rect 9254 6930 9282 7630
rect 9310 7657 9338 7966
rect 9310 7631 9311 7657
rect 9337 7631 9338 7657
rect 9310 7625 9338 7631
rect 9366 7574 9394 9422
rect 9422 9394 9450 9479
rect 9478 9506 9506 9511
rect 9478 9505 9562 9506
rect 9478 9479 9479 9505
rect 9505 9479 9562 9505
rect 9478 9478 9562 9479
rect 9478 9473 9506 9478
rect 9422 9366 9506 9394
rect 9422 9170 9450 9175
rect 9422 9123 9450 9142
rect 9422 8946 9450 8951
rect 9422 7657 9450 8918
rect 9478 8890 9506 9366
rect 9534 9002 9562 9478
rect 9646 9338 9674 9591
rect 9646 9305 9674 9310
rect 9758 9506 9786 9511
rect 9534 8969 9562 8974
rect 9646 9226 9674 9231
rect 9534 8890 9562 8895
rect 9478 8862 9534 8890
rect 9534 8857 9562 8862
rect 9590 8834 9618 8839
rect 9590 8787 9618 8806
rect 9646 8777 9674 9198
rect 9758 8833 9786 9478
rect 9758 8807 9759 8833
rect 9785 8807 9786 8833
rect 9758 8801 9786 8807
rect 9646 8751 9647 8777
rect 9673 8751 9674 8777
rect 9646 8722 9674 8751
rect 9674 8694 9730 8722
rect 9646 8689 9674 8694
rect 9702 8330 9730 8694
rect 9814 8441 9842 9926
rect 9926 9562 9954 9567
rect 9926 9515 9954 9534
rect 10038 9505 10066 10094
rect 10318 9954 10346 9959
rect 10318 9907 10346 9926
rect 10374 9842 10402 9847
rect 10374 9617 10402 9814
rect 10374 9591 10375 9617
rect 10401 9591 10402 9617
rect 10038 9479 10039 9505
rect 10065 9479 10066 9505
rect 10038 9473 10066 9479
rect 10206 9561 10234 9567
rect 10206 9535 10207 9561
rect 10233 9535 10234 9561
rect 9918 9422 10050 9427
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 9918 9389 10050 9394
rect 9870 9338 9898 9343
rect 9870 9225 9898 9310
rect 10206 9338 10234 9535
rect 10206 9305 10234 9310
rect 10318 9562 10346 9567
rect 9870 9199 9871 9225
rect 9897 9199 9898 9225
rect 9870 9193 9898 9199
rect 10150 9226 10178 9231
rect 10150 9179 10178 9198
rect 10262 9226 10290 9231
rect 10262 9179 10290 9198
rect 10094 9169 10122 9175
rect 10094 9143 10095 9169
rect 10121 9143 10122 9169
rect 9982 9114 10010 9119
rect 9926 9058 9954 9063
rect 9870 8946 9898 8951
rect 9870 8833 9898 8918
rect 9926 8889 9954 9030
rect 9926 8863 9927 8889
rect 9953 8863 9954 8889
rect 9926 8857 9954 8863
rect 9870 8807 9871 8833
rect 9897 8807 9898 8833
rect 9870 8801 9898 8807
rect 9982 8777 10010 9086
rect 10094 8834 10122 9143
rect 9982 8751 9983 8777
rect 10009 8751 10010 8777
rect 9982 8745 10010 8751
rect 10038 8806 10122 8834
rect 10262 8834 10290 8839
rect 10318 8834 10346 9534
rect 10374 9282 10402 9591
rect 10374 9249 10402 9254
rect 10430 9281 10458 9287
rect 10430 9255 10431 9281
rect 10457 9255 10458 9281
rect 10262 8833 10346 8834
rect 10262 8807 10263 8833
rect 10289 8807 10346 8833
rect 10262 8806 10346 8807
rect 10038 8777 10066 8806
rect 10262 8801 10290 8806
rect 10038 8751 10039 8777
rect 10065 8751 10066 8777
rect 10038 8745 10066 8751
rect 9918 8638 10050 8643
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 9918 8605 10050 8610
rect 9814 8415 9815 8441
rect 9841 8415 9842 8441
rect 9814 8409 9842 8415
rect 10430 8330 10458 9255
rect 10542 9170 10570 10262
rect 10710 10234 10738 10318
rect 10710 10201 10738 10206
rect 10598 9338 10626 9343
rect 10598 9225 10626 9310
rect 10598 9199 10599 9225
rect 10625 9199 10626 9225
rect 10598 9193 10626 9199
rect 10542 9123 10570 9142
rect 10654 9002 10682 9007
rect 10654 8833 10682 8974
rect 10710 8890 10738 8895
rect 10766 8890 10794 11942
rect 10822 11969 10906 11970
rect 10822 11943 10823 11969
rect 10849 11943 10906 11969
rect 10822 11942 10906 11943
rect 10822 11937 10850 11942
rect 10878 11466 10906 11942
rect 10934 11746 10962 11751
rect 10934 11633 10962 11718
rect 10934 11607 10935 11633
rect 10961 11607 10962 11633
rect 10934 11601 10962 11607
rect 10878 11438 10962 11466
rect 10878 11241 10906 11247
rect 10878 11215 10879 11241
rect 10905 11215 10906 11241
rect 10878 11074 10906 11215
rect 10878 11041 10906 11046
rect 10934 10906 10962 11438
rect 10934 10873 10962 10878
rect 10822 10850 10850 10855
rect 10822 10803 10850 10822
rect 10934 10402 10962 10407
rect 10766 8862 10850 8890
rect 10710 8843 10738 8862
rect 10654 8807 10655 8833
rect 10681 8807 10682 8833
rect 10654 8801 10682 8807
rect 10766 8777 10794 8783
rect 10766 8751 10767 8777
rect 10793 8751 10794 8777
rect 9702 8302 9842 8330
rect 9758 7994 9786 7999
rect 9758 7947 9786 7966
rect 9814 7993 9842 8302
rect 9926 8050 9954 8055
rect 9926 8003 9954 8022
rect 10430 7994 10458 8302
rect 9814 7967 9815 7993
rect 9841 7967 9842 7993
rect 9814 7961 9842 7967
rect 10374 7966 10458 7994
rect 10654 8722 10682 8727
rect 9918 7854 10050 7859
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 9918 7821 10050 7826
rect 9814 7713 9842 7719
rect 9814 7687 9815 7713
rect 9841 7687 9842 7713
rect 9422 7631 9423 7657
rect 9449 7631 9450 7657
rect 9422 7625 9450 7631
rect 9646 7657 9674 7663
rect 9646 7631 9647 7657
rect 9673 7631 9674 7657
rect 9646 7574 9674 7631
rect 9366 7546 9674 7574
rect 9814 7658 9842 7687
rect 9198 6929 9282 6930
rect 9198 6903 9199 6929
rect 9225 6903 9282 6929
rect 9198 6902 9282 6903
rect 9478 7321 9506 7327
rect 9478 7295 9479 7321
rect 9505 7295 9506 7321
rect 9478 6930 9506 7295
rect 9814 7322 9842 7630
rect 10318 7657 10346 7663
rect 10318 7631 10319 7657
rect 10345 7631 10346 7657
rect 10318 7602 10346 7631
rect 10374 7658 10402 7966
rect 10430 7770 10458 7775
rect 10430 7723 10458 7742
rect 10654 7769 10682 8694
rect 10710 8050 10738 8055
rect 10766 8050 10794 8751
rect 10738 8022 10794 8050
rect 10710 8003 10738 8022
rect 10822 7994 10850 8862
rect 10878 8834 10906 8853
rect 10878 8801 10906 8806
rect 10878 8722 10906 8727
rect 10934 8722 10962 10374
rect 10990 10401 11018 12222
rect 11046 12081 11074 12671
rect 12110 12474 12138 12783
rect 12110 12441 12138 12446
rect 12222 13201 12306 13202
rect 12222 13175 12279 13201
rect 12305 13175 12306 13201
rect 12222 13174 12306 13175
rect 11046 12055 11047 12081
rect 11073 12055 11074 12081
rect 11046 12049 11074 12055
rect 11102 12250 11130 12255
rect 11102 12081 11130 12222
rect 11102 12055 11103 12081
rect 11129 12055 11130 12081
rect 11102 12049 11130 12055
rect 11046 11969 11074 11975
rect 11046 11943 11047 11969
rect 11073 11943 11074 11969
rect 11046 10850 11074 11943
rect 12222 11690 12250 13174
rect 12278 13169 12306 13174
rect 12334 13201 12362 13790
rect 12950 13818 12978 13823
rect 12950 13771 12978 13790
rect 13062 13538 13090 13902
rect 13454 13593 13482 14014
rect 17598 13734 17730 13739
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17598 13701 17730 13706
rect 13454 13567 13455 13593
rect 13481 13567 13482 13593
rect 13454 13561 13482 13567
rect 20006 13593 20034 13599
rect 20006 13567 20007 13593
rect 20033 13567 20034 13593
rect 12334 13175 12335 13201
rect 12361 13175 12362 13201
rect 12334 13169 12362 13175
rect 12390 13481 12418 13487
rect 12390 13455 12391 13481
rect 12417 13455 12418 13481
rect 12278 13034 12306 13039
rect 12390 13034 12418 13455
rect 13062 13454 13090 13510
rect 18830 13537 18858 13543
rect 18830 13511 18831 13537
rect 18857 13511 18858 13537
rect 13062 13426 13202 13454
rect 12278 13033 12418 13034
rect 12278 13007 12279 13033
rect 12305 13007 12418 13033
rect 12278 13006 12418 13007
rect 12614 13145 12642 13151
rect 12614 13119 12615 13145
rect 12641 13119 12642 13145
rect 12278 13001 12306 13006
rect 12334 12810 12362 12815
rect 12334 12763 12362 12782
rect 12614 12810 12642 13119
rect 13006 13090 13034 13095
rect 12950 13089 13034 13090
rect 12950 13063 13007 13089
rect 13033 13063 13034 13089
rect 12950 13062 13034 13063
rect 12950 12865 12978 13062
rect 13006 13057 13034 13062
rect 12950 12839 12951 12865
rect 12977 12839 12978 12865
rect 12950 12833 12978 12839
rect 12614 12777 12642 12782
rect 13174 12753 13202 13426
rect 13174 12727 13175 12753
rect 13201 12727 13202 12753
rect 13174 12721 13202 12727
rect 13230 13090 13258 13095
rect 13006 12697 13034 12703
rect 13006 12671 13007 12697
rect 13033 12671 13034 12697
rect 12950 12641 12978 12647
rect 12950 12615 12951 12641
rect 12977 12615 12978 12641
rect 12222 11410 12250 11662
rect 12222 11377 12250 11382
rect 12278 11746 12306 11751
rect 11046 10817 11074 10822
rect 11102 11186 11130 11191
rect 10990 10375 10991 10401
rect 11017 10375 11018 10401
rect 10990 10122 11018 10375
rect 10990 10089 11018 10094
rect 11046 10345 11074 10351
rect 11046 10319 11047 10345
rect 11073 10319 11074 10345
rect 11046 9562 11074 10319
rect 11102 9674 11130 11158
rect 12278 11186 12306 11718
rect 12838 11577 12866 11583
rect 12838 11551 12839 11577
rect 12865 11551 12866 11577
rect 12670 11522 12698 11527
rect 12838 11522 12866 11551
rect 12670 11521 12866 11522
rect 12670 11495 12671 11521
rect 12697 11495 12866 11521
rect 12670 11494 12866 11495
rect 12558 11186 12586 11191
rect 12670 11186 12698 11494
rect 12782 11410 12810 11415
rect 12782 11241 12810 11382
rect 12782 11215 12783 11241
rect 12809 11215 12810 11241
rect 12782 11209 12810 11215
rect 12278 11185 12698 11186
rect 12278 11159 12279 11185
rect 12305 11159 12559 11185
rect 12585 11159 12698 11185
rect 12278 11158 12698 11159
rect 12278 11153 12306 11158
rect 11942 11129 11970 11135
rect 11942 11103 11943 11129
rect 11969 11103 11970 11129
rect 11494 11074 11522 11079
rect 11382 10906 11410 10911
rect 11382 10849 11410 10878
rect 11382 10823 11383 10849
rect 11409 10823 11410 10849
rect 11270 10794 11298 10799
rect 11270 10747 11298 10766
rect 11382 10682 11410 10823
rect 11494 10793 11522 11046
rect 11942 10905 11970 11103
rect 11942 10879 11943 10905
rect 11969 10879 11970 10905
rect 11942 10873 11970 10879
rect 12334 10905 12362 11158
rect 12558 11153 12586 11158
rect 12334 10879 12335 10905
rect 12361 10879 12362 10905
rect 12334 10873 12362 10879
rect 11550 10850 11578 10855
rect 11550 10803 11578 10822
rect 11494 10767 11495 10793
rect 11521 10767 11522 10793
rect 11494 10761 11522 10767
rect 11774 10793 11802 10799
rect 11774 10767 11775 10793
rect 11801 10767 11802 10793
rect 11662 10738 11690 10743
rect 11774 10738 11802 10767
rect 11662 10737 11802 10738
rect 11662 10711 11663 10737
rect 11689 10711 11802 10737
rect 11662 10710 11802 10711
rect 11942 10793 11970 10799
rect 11942 10767 11943 10793
rect 11969 10767 11970 10793
rect 11662 10705 11690 10710
rect 11382 10654 11634 10682
rect 11270 10402 11298 10407
rect 11550 10402 11578 10407
rect 11270 10401 11578 10402
rect 11270 10375 11271 10401
rect 11297 10375 11551 10401
rect 11577 10375 11578 10401
rect 11270 10374 11578 10375
rect 11270 10369 11298 10374
rect 11550 10369 11578 10374
rect 11606 10345 11634 10654
rect 11942 10570 11970 10767
rect 11942 10537 11970 10542
rect 12054 10793 12082 10799
rect 12054 10767 12055 10793
rect 12081 10767 12082 10793
rect 12054 10458 12082 10767
rect 12838 10793 12866 11494
rect 12838 10767 12839 10793
rect 12865 10767 12866 10793
rect 12838 10761 12866 10767
rect 12894 11186 12922 11191
rect 12950 11186 12978 12615
rect 13006 12642 13034 12671
rect 13230 12697 13258 13062
rect 14070 13090 14098 13095
rect 14070 13043 14098 13062
rect 18830 13090 18858 13511
rect 20006 13146 20034 13567
rect 20006 13113 20034 13118
rect 18830 13057 18858 13062
rect 17598 12950 17730 12955
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17598 12917 17730 12922
rect 13230 12671 13231 12697
rect 13257 12671 13258 12697
rect 13230 12665 13258 12671
rect 13342 12642 13370 12647
rect 13006 12614 13202 12642
rect 13174 12586 13202 12614
rect 13286 12641 13370 12642
rect 13286 12615 13343 12641
rect 13369 12615 13370 12641
rect 13286 12614 13370 12615
rect 13286 12586 13314 12614
rect 13342 12609 13370 12614
rect 13174 12558 13314 12586
rect 17598 12166 17730 12171
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17598 12133 17730 12138
rect 20006 12025 20034 12031
rect 20006 11999 20007 12025
rect 20033 11999 20034 12025
rect 13454 11970 13482 11975
rect 13454 11913 13482 11942
rect 14518 11970 14546 11975
rect 13454 11887 13455 11913
rect 13481 11887 13482 11913
rect 13454 11881 13482 11887
rect 13510 11914 13538 11919
rect 13510 11913 13594 11914
rect 13510 11887 13511 11913
rect 13537 11887 13594 11913
rect 13510 11886 13594 11887
rect 13510 11881 13538 11886
rect 13342 11857 13370 11863
rect 13342 11831 13343 11857
rect 13369 11831 13370 11857
rect 13342 11634 13370 11831
rect 13342 11606 13538 11634
rect 13230 11522 13258 11527
rect 13230 11521 13482 11522
rect 13230 11495 13231 11521
rect 13257 11495 13482 11521
rect 13230 11494 13482 11495
rect 13230 11489 13258 11494
rect 13062 11242 13090 11247
rect 13062 11241 13370 11242
rect 13062 11215 13063 11241
rect 13089 11215 13370 11241
rect 13062 11214 13370 11215
rect 13062 11209 13090 11214
rect 12894 11185 12978 11186
rect 12894 11159 12895 11185
rect 12921 11159 12978 11185
rect 12894 11158 12978 11159
rect 13342 11185 13370 11214
rect 13454 11241 13482 11494
rect 13454 11215 13455 11241
rect 13481 11215 13482 11241
rect 13454 11209 13482 11215
rect 13342 11159 13343 11185
rect 13369 11159 13370 11185
rect 12894 10514 12922 11158
rect 13342 11153 13370 11159
rect 13510 11185 13538 11606
rect 13510 11159 13511 11185
rect 13537 11159 13538 11185
rect 13510 11153 13538 11159
rect 13230 11129 13258 11135
rect 13230 11103 13231 11129
rect 13257 11103 13258 11129
rect 13174 10738 13202 10743
rect 12838 10486 12922 10514
rect 13006 10737 13202 10738
rect 13006 10711 13175 10737
rect 13201 10711 13202 10737
rect 13006 10710 13202 10711
rect 11942 10430 12082 10458
rect 12222 10458 12250 10463
rect 11886 10402 11914 10407
rect 11606 10319 11607 10345
rect 11633 10319 11634 10345
rect 11606 10313 11634 10319
rect 11662 10346 11690 10351
rect 11662 10299 11690 10318
rect 11718 10345 11746 10351
rect 11718 10319 11719 10345
rect 11745 10319 11746 10345
rect 11382 10289 11410 10295
rect 11382 10263 11383 10289
rect 11409 10263 11410 10289
rect 11270 10234 11298 10239
rect 11102 9641 11130 9646
rect 11158 10178 11186 10183
rect 11046 9529 11074 9534
rect 11102 9506 11130 9511
rect 11158 9506 11186 10150
rect 11102 9505 11186 9506
rect 11102 9479 11103 9505
rect 11129 9479 11186 9505
rect 11102 9478 11186 9479
rect 10906 8694 10962 8722
rect 10990 8946 11018 8951
rect 10990 8722 11018 8918
rect 11046 8834 11074 8839
rect 11102 8834 11130 9478
rect 11158 9226 11186 9231
rect 11158 9114 11186 9198
rect 11270 9225 11298 10206
rect 11270 9199 11271 9225
rect 11297 9199 11298 9225
rect 11270 9193 11298 9199
rect 11326 10122 11354 10127
rect 11326 9561 11354 10094
rect 11326 9535 11327 9561
rect 11353 9535 11354 9561
rect 11326 9170 11354 9535
rect 11382 9282 11410 10263
rect 11494 10290 11522 10295
rect 11494 10243 11522 10262
rect 11718 10122 11746 10319
rect 11718 10089 11746 10094
rect 11606 9842 11634 9847
rect 11382 9249 11410 9254
rect 11550 9674 11578 9679
rect 11550 9561 11578 9646
rect 11606 9617 11634 9814
rect 11606 9591 11607 9617
rect 11633 9591 11634 9617
rect 11606 9585 11634 9591
rect 11550 9535 11551 9561
rect 11577 9535 11578 9561
rect 11494 9170 11522 9175
rect 11326 9169 11522 9170
rect 11326 9143 11495 9169
rect 11521 9143 11522 9169
rect 11326 9142 11522 9143
rect 11326 9114 11354 9142
rect 11494 9137 11522 9142
rect 11158 9086 11354 9114
rect 11046 8833 11130 8834
rect 11046 8807 11047 8833
rect 11073 8807 11130 8833
rect 11046 8806 11130 8807
rect 11326 9002 11354 9007
rect 11326 8833 11354 8974
rect 11326 8807 11327 8833
rect 11353 8807 11354 8833
rect 11046 8801 11074 8806
rect 11326 8801 11354 8807
rect 11214 8722 11242 8727
rect 10990 8721 11242 8722
rect 10990 8695 11215 8721
rect 11241 8695 11242 8721
rect 10990 8694 11242 8695
rect 10878 8689 10906 8694
rect 10990 8554 11018 8694
rect 11214 8689 11242 8694
rect 11550 8610 11578 9535
rect 11774 9561 11802 9567
rect 11774 9535 11775 9561
rect 11801 9535 11802 9561
rect 11774 9506 11802 9535
rect 11886 9561 11914 10374
rect 11942 9730 11970 10430
rect 12222 10411 12250 10430
rect 12166 10402 12194 10407
rect 12054 10345 12082 10351
rect 12054 10319 12055 10345
rect 12081 10319 12082 10345
rect 12054 9842 12082 10319
rect 12166 10345 12194 10374
rect 12166 10319 12167 10345
rect 12193 10319 12194 10345
rect 12166 10313 12194 10319
rect 12838 10178 12866 10486
rect 13006 10457 13034 10710
rect 13174 10705 13202 10710
rect 13006 10431 13007 10457
rect 13033 10431 13034 10457
rect 13006 10425 13034 10431
rect 13174 10458 13202 10463
rect 13230 10458 13258 11103
rect 13566 10850 13594 11886
rect 14518 11578 14546 11942
rect 18830 11970 18858 11975
rect 18830 11923 18858 11942
rect 20006 11802 20034 11999
rect 20006 11769 20034 11774
rect 14630 11634 14658 11639
rect 14630 11587 14658 11606
rect 14294 11577 14546 11578
rect 14294 11551 14519 11577
rect 14545 11551 14546 11577
rect 14294 11550 14546 11551
rect 14294 11521 14322 11550
rect 14518 11545 14546 11550
rect 18830 11578 18858 11583
rect 18830 11531 18858 11550
rect 14294 11495 14295 11521
rect 14321 11495 14322 11521
rect 14294 11489 14322 11495
rect 20006 11466 20034 11471
rect 20006 11419 20034 11438
rect 17598 11382 17730 11387
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17598 11349 17730 11354
rect 20006 11241 20034 11247
rect 20006 11215 20007 11241
rect 20033 11215 20034 11241
rect 18830 11186 18858 11191
rect 18830 11139 18858 11158
rect 20006 11130 20034 11215
rect 20006 11097 20034 11102
rect 13202 10430 13258 10458
rect 13454 10457 13482 10463
rect 13454 10431 13455 10457
rect 13481 10431 13482 10457
rect 12838 10145 12866 10150
rect 12894 10401 12922 10407
rect 12894 10375 12895 10401
rect 12921 10375 12922 10401
rect 12054 9809 12082 9814
rect 12222 9953 12250 9959
rect 12222 9927 12223 9953
rect 12249 9927 12250 9953
rect 11942 9729 12082 9730
rect 11942 9703 11943 9729
rect 11969 9703 12082 9729
rect 11942 9702 12082 9703
rect 11942 9697 11970 9702
rect 11886 9535 11887 9561
rect 11913 9535 11914 9561
rect 11886 9529 11914 9535
rect 11774 9473 11802 9478
rect 12054 9337 12082 9702
rect 12222 9618 12250 9927
rect 12278 9618 12306 9623
rect 12222 9617 12306 9618
rect 12222 9591 12279 9617
rect 12305 9591 12306 9617
rect 12222 9590 12306 9591
rect 12054 9311 12055 9337
rect 12081 9311 12082 9337
rect 11942 9282 11970 9287
rect 11942 9225 11970 9254
rect 11942 9199 11943 9225
rect 11969 9199 11970 9225
rect 11942 9193 11970 9199
rect 11998 8946 12026 8951
rect 12054 8946 12082 9311
rect 12110 9562 12138 9567
rect 12110 9169 12138 9534
rect 12110 9143 12111 9169
rect 12137 9143 12138 9169
rect 12110 9137 12138 9143
rect 11998 8945 12082 8946
rect 11998 8919 11999 8945
rect 12025 8919 12082 8945
rect 11998 8918 12082 8919
rect 11998 8913 12026 8918
rect 11886 8890 11914 8895
rect 11886 8843 11914 8862
rect 11830 8833 11858 8839
rect 11830 8807 11831 8833
rect 11857 8807 11858 8833
rect 11550 8577 11578 8582
rect 11606 8722 11634 8727
rect 10654 7743 10655 7769
rect 10681 7743 10682 7769
rect 10654 7737 10682 7743
rect 10766 7993 10850 7994
rect 10766 7967 10823 7993
rect 10849 7967 10850 7993
rect 10766 7966 10850 7967
rect 10766 7770 10794 7966
rect 10822 7961 10850 7966
rect 10934 8526 11018 8554
rect 10794 7742 10850 7770
rect 10766 7723 10794 7742
rect 10486 7658 10514 7663
rect 10374 7657 10514 7658
rect 10374 7631 10487 7657
rect 10513 7631 10514 7657
rect 10374 7630 10514 7631
rect 10486 7625 10514 7630
rect 10318 7569 10346 7574
rect 10710 7601 10738 7607
rect 10710 7575 10711 7601
rect 10737 7575 10738 7601
rect 9814 7289 9842 7294
rect 9702 7266 9730 7271
rect 9702 7219 9730 7238
rect 10206 7266 10234 7271
rect 9918 7070 10050 7075
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 9918 7037 10050 7042
rect 9534 6930 9562 6935
rect 9478 6902 9534 6930
rect 9198 6897 9226 6902
rect 8302 6818 8330 6823
rect 8190 6817 8330 6818
rect 8190 6791 8303 6817
rect 8329 6791 8330 6817
rect 8190 6790 8330 6791
rect 8302 6762 8330 6790
rect 8302 6734 8442 6762
rect 2238 6678 2370 6683
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2238 6645 2370 6650
rect 2238 5894 2370 5899
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2238 5861 2370 5866
rect 2238 5110 2370 5115
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2238 5077 2370 5082
rect 2238 4326 2370 4331
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2238 4293 2370 4298
rect 8414 4214 8442 6734
rect 8414 4186 8554 4214
rect 2238 3542 2370 3547
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2238 3509 2370 3514
rect 2238 2758 2370 2763
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2238 2725 2370 2730
rect 2238 1974 2370 1979
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2238 1941 2370 1946
rect 8526 1777 8554 4186
rect 9534 2169 9562 6902
rect 10206 6874 10234 7238
rect 10430 7266 10458 7271
rect 10598 7266 10626 7271
rect 10430 7265 10626 7266
rect 10430 7239 10431 7265
rect 10457 7239 10599 7265
rect 10625 7239 10626 7265
rect 10430 7238 10626 7239
rect 10430 7233 10458 7238
rect 10598 7233 10626 7238
rect 10262 7210 10290 7215
rect 10262 7163 10290 7182
rect 10206 6827 10234 6846
rect 10318 7153 10346 7159
rect 10318 7127 10319 7153
rect 10345 7127 10346 7153
rect 9918 6286 10050 6291
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 9918 6253 10050 6258
rect 9758 6033 9786 6039
rect 9758 6007 9759 6033
rect 9785 6007 9786 6033
rect 9758 5978 9786 6007
rect 9758 5945 9786 5950
rect 10318 5978 10346 7127
rect 10542 6930 10570 6935
rect 10710 6930 10738 7575
rect 10822 7265 10850 7742
rect 10822 7239 10823 7265
rect 10849 7239 10850 7265
rect 10822 7233 10850 7239
rect 10934 7265 10962 8526
rect 11606 8497 11634 8694
rect 11606 8471 11607 8497
rect 11633 8471 11634 8497
rect 10990 7657 11018 7663
rect 10990 7631 10991 7657
rect 11017 7631 11018 7657
rect 10990 7574 11018 7631
rect 10990 7546 11186 7574
rect 11158 7377 11186 7546
rect 11158 7351 11159 7377
rect 11185 7351 11186 7377
rect 11158 7345 11186 7351
rect 11606 7322 11634 8471
rect 11830 8386 11858 8807
rect 12222 8833 12250 9590
rect 12278 9585 12306 9590
rect 12670 9562 12698 9567
rect 12670 9515 12698 9534
rect 12894 9058 12922 10375
rect 13118 10402 13146 10407
rect 13118 10355 13146 10374
rect 13174 10401 13202 10430
rect 13174 10375 13175 10401
rect 13201 10375 13202 10401
rect 13174 10369 13202 10375
rect 13342 10401 13370 10407
rect 13342 10375 13343 10401
rect 13369 10375 13370 10401
rect 13342 10178 13370 10375
rect 13454 10402 13482 10431
rect 13454 10369 13482 10374
rect 13510 10402 13538 10407
rect 13566 10402 13594 10822
rect 18830 10794 18858 10799
rect 18830 10747 18858 10766
rect 20006 10794 20034 10799
rect 13510 10401 13594 10402
rect 13510 10375 13511 10401
rect 13537 10375 13594 10401
rect 13510 10374 13594 10375
rect 13622 10738 13650 10743
rect 13510 10369 13538 10374
rect 13622 10345 13650 10710
rect 14238 10738 14266 10743
rect 14238 10691 14266 10710
rect 20006 10737 20034 10766
rect 20006 10711 20007 10737
rect 20033 10711 20034 10737
rect 20006 10705 20034 10711
rect 17598 10598 17730 10603
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17598 10565 17730 10570
rect 13622 10319 13623 10345
rect 13649 10319 13650 10345
rect 13622 10313 13650 10319
rect 13734 10346 13762 10351
rect 13342 10145 13370 10150
rect 13734 9674 13762 10318
rect 18830 10009 18858 10015
rect 18830 9983 18831 10009
rect 18857 9983 18858 10009
rect 17598 9814 17730 9819
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17598 9781 17730 9786
rect 13734 9627 13762 9646
rect 18830 9674 18858 9983
rect 20006 9897 20034 9903
rect 20006 9871 20007 9897
rect 20033 9871 20034 9897
rect 20006 9786 20034 9871
rect 20006 9753 20034 9758
rect 18830 9641 18858 9646
rect 12894 9025 12922 9030
rect 17598 9030 17730 9035
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17598 8997 17730 9002
rect 12222 8807 12223 8833
rect 12249 8807 12250 8833
rect 12054 8778 12082 8783
rect 12054 8731 12082 8750
rect 12222 8722 12250 8807
rect 13678 8889 13706 8895
rect 13678 8863 13679 8889
rect 13705 8863 13706 8889
rect 13678 8834 13706 8863
rect 20006 8889 20034 8895
rect 20006 8863 20007 8889
rect 20033 8863 20034 8889
rect 13902 8834 13930 8839
rect 13678 8833 13930 8834
rect 13678 8807 13903 8833
rect 13929 8807 13930 8833
rect 13678 8806 13930 8807
rect 12614 8778 12642 8783
rect 12614 8731 12642 8750
rect 12222 8689 12250 8694
rect 12782 8666 12810 8671
rect 11830 8353 11858 8358
rect 12222 8610 12250 8615
rect 12222 8161 12250 8582
rect 12782 8441 12810 8638
rect 13902 8666 13930 8806
rect 18830 8833 18858 8839
rect 18830 8807 18831 8833
rect 18857 8807 18858 8833
rect 14014 8722 14042 8727
rect 14014 8675 14042 8694
rect 13902 8633 13930 8638
rect 18830 8666 18858 8807
rect 20006 8778 20034 8863
rect 20006 8745 20034 8750
rect 18830 8633 18858 8638
rect 18942 8722 18970 8727
rect 12782 8415 12783 8441
rect 12809 8415 12810 8441
rect 12782 8409 12810 8415
rect 18942 8441 18970 8694
rect 18942 8415 18943 8441
rect 18969 8415 18970 8441
rect 18942 8409 18970 8415
rect 20006 8442 20034 8447
rect 12670 8386 12698 8391
rect 12670 8339 12698 8358
rect 20006 8385 20034 8414
rect 20006 8359 20007 8385
rect 20033 8359 20034 8385
rect 20006 8353 20034 8359
rect 12222 8135 12223 8161
rect 12249 8135 12250 8161
rect 12222 8129 12250 8135
rect 12614 8330 12642 8335
rect 12390 8106 12418 8111
rect 12558 8106 12586 8111
rect 12390 8105 12586 8106
rect 12390 8079 12391 8105
rect 12417 8079 12559 8105
rect 12585 8079 12586 8105
rect 12390 8078 12586 8079
rect 12390 8073 12418 8078
rect 12558 8073 12586 8078
rect 12614 8050 12642 8302
rect 17598 8246 17730 8251
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17598 8213 17730 8218
rect 12614 8022 12698 8050
rect 12670 7993 12698 8022
rect 12670 7967 12671 7993
rect 12697 7967 12698 7993
rect 12670 7961 12698 7967
rect 12334 7937 12362 7943
rect 12614 7938 12642 7943
rect 12334 7911 12335 7937
rect 12361 7911 12362 7937
rect 12334 7714 12362 7911
rect 12334 7681 12362 7686
rect 12502 7937 12642 7938
rect 12502 7911 12615 7937
rect 12641 7911 12642 7937
rect 12502 7910 12642 7911
rect 12502 7574 12530 7910
rect 12614 7905 12642 7910
rect 12278 7546 12530 7574
rect 12614 7714 12642 7719
rect 11662 7322 11690 7327
rect 12222 7322 12250 7327
rect 12278 7322 12306 7546
rect 10934 7239 10935 7265
rect 10961 7239 10962 7265
rect 10934 7233 10962 7239
rect 11438 7321 11858 7322
rect 11438 7295 11663 7321
rect 11689 7295 11858 7321
rect 11438 7294 11858 7295
rect 11102 7210 11130 7215
rect 11102 7163 11130 7182
rect 10542 6929 10738 6930
rect 10542 6903 10543 6929
rect 10569 6903 10738 6929
rect 10542 6902 10738 6903
rect 10878 7153 10906 7159
rect 10878 7127 10879 7153
rect 10905 7127 10906 7153
rect 10542 6897 10570 6902
rect 10822 6146 10850 6151
rect 10878 6146 10906 7127
rect 11158 7153 11186 7159
rect 11158 7127 11159 7153
rect 11185 7127 11186 7153
rect 11158 6762 11186 7127
rect 11158 6729 11186 6734
rect 11438 6874 11466 7294
rect 11662 7289 11690 7294
rect 11830 7265 11858 7294
rect 12222 7321 12306 7322
rect 12222 7295 12223 7321
rect 12249 7295 12306 7321
rect 12222 7294 12306 7295
rect 12222 7289 12250 7294
rect 11830 7239 11831 7265
rect 11857 7239 11858 7265
rect 11830 6985 11858 7239
rect 11830 6959 11831 6985
rect 11857 6959 11858 6985
rect 11830 6953 11858 6959
rect 11438 6202 11466 6846
rect 11606 6817 11634 6823
rect 11606 6791 11607 6817
rect 11633 6791 11634 6817
rect 11606 6762 11634 6791
rect 11606 6729 11634 6734
rect 12278 6762 12306 6767
rect 10822 6145 10906 6146
rect 10822 6119 10823 6145
rect 10849 6119 10906 6145
rect 10822 6118 10906 6119
rect 11214 6201 11466 6202
rect 11214 6175 11439 6201
rect 11465 6175 11466 6201
rect 11214 6174 11466 6175
rect 10822 6113 10850 6118
rect 11214 6089 11242 6174
rect 11438 6169 11466 6174
rect 11214 6063 11215 6089
rect 11241 6063 11242 6089
rect 11214 6057 11242 6063
rect 10318 5945 10346 5950
rect 10710 5978 10738 5983
rect 9918 5502 10050 5507
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 9918 5469 10050 5474
rect 9918 4718 10050 4723
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 9918 4685 10050 4690
rect 9918 3934 10050 3939
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 9918 3901 10050 3906
rect 9918 3150 10050 3155
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 9918 3117 10050 3122
rect 9918 2366 10050 2371
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 9918 2333 10050 2338
rect 9534 2143 9535 2169
rect 9561 2143 9562 2169
rect 9534 2137 9562 2143
rect 8526 1751 8527 1777
rect 8553 1751 8554 1777
rect 8526 1745 8554 1751
rect 9422 2058 9450 2063
rect 8414 1722 8442 1727
rect 8414 400 8442 1694
rect 9030 1722 9058 1727
rect 9030 1665 9058 1694
rect 9030 1639 9031 1665
rect 9057 1639 9058 1665
rect 9030 1633 9058 1639
rect 9422 400 9450 2030
rect 10038 2058 10066 2063
rect 10038 2011 10066 2030
rect 10710 1777 10738 5950
rect 10710 1751 10711 1777
rect 10737 1751 10738 1777
rect 10710 1745 10738 1751
rect 11438 1834 11466 1839
rect 11214 1666 11242 1671
rect 11102 1665 11242 1666
rect 11102 1639 11215 1665
rect 11241 1639 11242 1665
rect 11102 1638 11242 1639
rect 9918 1582 10050 1587
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 9918 1549 10050 1554
rect 11102 400 11130 1638
rect 11214 1633 11242 1638
rect 11438 400 11466 1806
rect 12278 1777 12306 6734
rect 12614 2169 12642 7686
rect 13286 7714 13314 7719
rect 13286 7321 13314 7686
rect 17598 7462 17730 7467
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17598 7429 17730 7434
rect 13286 7295 13287 7321
rect 13313 7295 13314 7321
rect 13286 7289 13314 7295
rect 17598 6678 17730 6683
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17598 6645 17730 6650
rect 17598 5894 17730 5899
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17598 5861 17730 5866
rect 17598 5110 17730 5115
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17598 5077 17730 5082
rect 17598 4326 17730 4331
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17598 4293 17730 4298
rect 17598 3542 17730 3547
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17598 3509 17730 3514
rect 17598 2758 17730 2763
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17598 2725 17730 2730
rect 12614 2143 12615 2169
rect 12641 2143 12642 2169
rect 12614 2137 12642 2143
rect 12278 1751 12279 1777
rect 12305 1751 12306 1777
rect 12278 1745 12306 1751
rect 12446 2058 12474 2063
rect 12446 400 12474 2030
rect 13118 2058 13146 2063
rect 13118 2011 13146 2030
rect 17598 1974 17730 1979
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17598 1941 17730 1946
rect 12782 1834 12810 1839
rect 12782 1787 12810 1806
rect 8400 0 8456 400
rect 9408 0 9464 400
rect 11088 0 11144 400
rect 11424 0 11480 400
rect 12432 0 12488 400
<< via2 >>
rect 2238 19221 2266 19222
rect 2238 19195 2239 19221
rect 2239 19195 2265 19221
rect 2265 19195 2266 19221
rect 2238 19194 2266 19195
rect 2290 19221 2318 19222
rect 2290 19195 2291 19221
rect 2291 19195 2317 19221
rect 2317 19195 2318 19221
rect 2290 19194 2318 19195
rect 2342 19221 2370 19222
rect 2342 19195 2343 19221
rect 2343 19195 2369 19221
rect 2369 19195 2370 19221
rect 2342 19194 2370 19195
rect 2238 18437 2266 18438
rect 2238 18411 2239 18437
rect 2239 18411 2265 18437
rect 2265 18411 2266 18437
rect 2238 18410 2266 18411
rect 2290 18437 2318 18438
rect 2290 18411 2291 18437
rect 2291 18411 2317 18437
rect 2317 18411 2318 18437
rect 2290 18410 2318 18411
rect 2342 18437 2370 18438
rect 2342 18411 2343 18437
rect 2343 18411 2369 18437
rect 2369 18411 2370 18437
rect 2342 18410 2370 18411
rect 854 18185 882 18186
rect 854 18159 855 18185
rect 855 18159 881 18185
rect 881 18159 882 18185
rect 854 18158 882 18159
rect 2238 17653 2266 17654
rect 2238 17627 2239 17653
rect 2239 17627 2265 17653
rect 2265 17627 2266 17653
rect 2238 17626 2266 17627
rect 2290 17653 2318 17654
rect 2290 17627 2291 17653
rect 2291 17627 2317 17653
rect 2317 17627 2318 17653
rect 2290 17626 2318 17627
rect 2342 17653 2370 17654
rect 2342 17627 2343 17653
rect 2343 17627 2369 17653
rect 2369 17627 2370 17653
rect 2342 17626 2370 17627
rect 2238 16869 2266 16870
rect 2238 16843 2239 16869
rect 2239 16843 2265 16869
rect 2265 16843 2266 16869
rect 2238 16842 2266 16843
rect 2290 16869 2318 16870
rect 2290 16843 2291 16869
rect 2291 16843 2317 16869
rect 2317 16843 2318 16869
rect 2290 16842 2318 16843
rect 2342 16869 2370 16870
rect 2342 16843 2343 16869
rect 2343 16843 2369 16869
rect 2369 16843 2370 16869
rect 2342 16842 2370 16843
rect 2238 16085 2266 16086
rect 2238 16059 2239 16085
rect 2239 16059 2265 16085
rect 2265 16059 2266 16085
rect 2238 16058 2266 16059
rect 2290 16085 2318 16086
rect 2290 16059 2291 16085
rect 2291 16059 2317 16085
rect 2317 16059 2318 16085
rect 2290 16058 2318 16059
rect 2342 16085 2370 16086
rect 2342 16059 2343 16085
rect 2343 16059 2369 16085
rect 2369 16059 2370 16085
rect 2342 16058 2370 16059
rect 2238 15301 2266 15302
rect 2238 15275 2239 15301
rect 2239 15275 2265 15301
rect 2265 15275 2266 15301
rect 2238 15274 2266 15275
rect 2290 15301 2318 15302
rect 2290 15275 2291 15301
rect 2291 15275 2317 15301
rect 2317 15275 2318 15301
rect 2290 15274 2318 15275
rect 2342 15301 2370 15302
rect 2342 15275 2343 15301
rect 2343 15275 2369 15301
rect 2369 15275 2370 15301
rect 2342 15274 2370 15275
rect 2238 14517 2266 14518
rect 2238 14491 2239 14517
rect 2239 14491 2265 14517
rect 2265 14491 2266 14517
rect 2238 14490 2266 14491
rect 2290 14517 2318 14518
rect 2290 14491 2291 14517
rect 2291 14491 2317 14517
rect 2317 14491 2318 14517
rect 2290 14490 2318 14491
rect 2342 14517 2370 14518
rect 2342 14491 2343 14517
rect 2343 14491 2369 14517
rect 2369 14491 2370 14517
rect 2342 14490 2370 14491
rect 9310 14294 9338 14322
rect 2086 13790 2114 13818
rect 966 12249 994 12250
rect 966 12223 967 12249
rect 967 12223 993 12249
rect 993 12223 994 12249
rect 966 12222 994 12223
rect 966 10430 994 10458
rect 1022 10094 1050 10122
rect 2238 13733 2266 13734
rect 2238 13707 2239 13733
rect 2239 13707 2265 13733
rect 2265 13707 2266 13733
rect 2238 13706 2266 13707
rect 2290 13733 2318 13734
rect 2290 13707 2291 13733
rect 2291 13707 2317 13733
rect 2317 13707 2318 13733
rect 2290 13706 2318 13707
rect 2342 13733 2370 13734
rect 2342 13707 2343 13733
rect 2343 13707 2369 13733
rect 2369 13707 2370 13733
rect 2342 13706 2370 13707
rect 8638 13593 8666 13594
rect 8638 13567 8639 13593
rect 8639 13567 8665 13593
rect 8665 13567 8666 13593
rect 8638 13566 8666 13567
rect 2238 12949 2266 12950
rect 2238 12923 2239 12949
rect 2239 12923 2265 12949
rect 2265 12923 2266 12949
rect 2238 12922 2266 12923
rect 2290 12949 2318 12950
rect 2290 12923 2291 12949
rect 2291 12923 2317 12949
rect 2317 12923 2318 12949
rect 2290 12922 2318 12923
rect 2342 12949 2370 12950
rect 2342 12923 2343 12949
rect 2343 12923 2369 12949
rect 2369 12923 2370 12949
rect 2342 12922 2370 12923
rect 2142 12361 2170 12362
rect 2142 12335 2143 12361
rect 2143 12335 2169 12361
rect 2169 12335 2170 12361
rect 2142 12334 2170 12335
rect 5614 12334 5642 12362
rect 7574 13230 7602 13258
rect 9918 18829 9946 18830
rect 9918 18803 9919 18829
rect 9919 18803 9945 18829
rect 9945 18803 9946 18829
rect 9918 18802 9946 18803
rect 9970 18829 9998 18830
rect 9970 18803 9971 18829
rect 9971 18803 9997 18829
rect 9997 18803 9998 18829
rect 9970 18802 9998 18803
rect 10022 18829 10050 18830
rect 10022 18803 10023 18829
rect 10023 18803 10049 18829
rect 10049 18803 10050 18829
rect 10022 18802 10050 18803
rect 11438 19110 11466 19138
rect 12782 19137 12810 19138
rect 12782 19111 12783 19137
rect 12783 19111 12809 19137
rect 12809 19111 12810 19137
rect 12782 19110 12810 19111
rect 10430 18718 10458 18746
rect 11046 18745 11074 18746
rect 11046 18719 11047 18745
rect 11047 18719 11073 18745
rect 11073 18719 11074 18745
rect 11046 18718 11074 18719
rect 10094 18326 10122 18354
rect 10150 18214 10178 18242
rect 9918 18045 9946 18046
rect 9918 18019 9919 18045
rect 9919 18019 9945 18045
rect 9945 18019 9946 18045
rect 9918 18018 9946 18019
rect 9970 18045 9998 18046
rect 9970 18019 9971 18045
rect 9971 18019 9997 18045
rect 9997 18019 9998 18045
rect 9970 18018 9998 18019
rect 10022 18045 10050 18046
rect 10022 18019 10023 18045
rect 10023 18019 10049 18045
rect 10049 18019 10050 18045
rect 10022 18018 10050 18019
rect 9918 17261 9946 17262
rect 9918 17235 9919 17261
rect 9919 17235 9945 17261
rect 9945 17235 9946 17261
rect 9918 17234 9946 17235
rect 9970 17261 9998 17262
rect 9970 17235 9971 17261
rect 9971 17235 9997 17261
rect 9997 17235 9998 17261
rect 9970 17234 9998 17235
rect 10022 17261 10050 17262
rect 10022 17235 10023 17261
rect 10023 17235 10049 17261
rect 10049 17235 10050 17261
rect 10022 17234 10050 17235
rect 9918 16477 9946 16478
rect 9918 16451 9919 16477
rect 9919 16451 9945 16477
rect 9945 16451 9946 16477
rect 9918 16450 9946 16451
rect 9970 16477 9998 16478
rect 9970 16451 9971 16477
rect 9971 16451 9997 16477
rect 9997 16451 9998 16477
rect 9970 16450 9998 16451
rect 10022 16477 10050 16478
rect 10022 16451 10023 16477
rect 10023 16451 10049 16477
rect 10049 16451 10050 16477
rect 10022 16450 10050 16451
rect 9918 15693 9946 15694
rect 9918 15667 9919 15693
rect 9919 15667 9945 15693
rect 9945 15667 9946 15693
rect 9918 15666 9946 15667
rect 9970 15693 9998 15694
rect 9970 15667 9971 15693
rect 9971 15667 9997 15693
rect 9997 15667 9998 15693
rect 9970 15666 9998 15667
rect 10022 15693 10050 15694
rect 10022 15667 10023 15693
rect 10023 15667 10049 15693
rect 10049 15667 10050 15693
rect 10022 15666 10050 15667
rect 9918 14909 9946 14910
rect 9918 14883 9919 14909
rect 9919 14883 9945 14909
rect 9945 14883 9946 14909
rect 9918 14882 9946 14883
rect 9970 14909 9998 14910
rect 9970 14883 9971 14909
rect 9971 14883 9997 14909
rect 9997 14883 9998 14909
rect 9970 14882 9998 14883
rect 10022 14909 10050 14910
rect 10022 14883 10023 14909
rect 10023 14883 10049 14909
rect 10049 14883 10050 14909
rect 10022 14882 10050 14883
rect 10038 14321 10066 14322
rect 10038 14295 10039 14321
rect 10039 14295 10065 14321
rect 10065 14295 10066 14321
rect 10038 14294 10066 14295
rect 9870 14238 9898 14266
rect 10150 14265 10178 14266
rect 10150 14239 10151 14265
rect 10151 14239 10177 14265
rect 10177 14239 10178 14265
rect 10150 14238 10178 14239
rect 9918 14125 9946 14126
rect 9918 14099 9919 14125
rect 9919 14099 9945 14125
rect 9945 14099 9946 14125
rect 9918 14098 9946 14099
rect 9970 14125 9998 14126
rect 9970 14099 9971 14125
rect 9971 14099 9997 14125
rect 9997 14099 9998 14125
rect 9970 14098 9998 14099
rect 10022 14125 10050 14126
rect 10022 14099 10023 14125
rect 10023 14099 10049 14125
rect 10049 14099 10050 14125
rect 10022 14098 10050 14099
rect 9982 14041 10010 14042
rect 9982 14015 9983 14041
rect 9983 14015 10009 14041
rect 10009 14015 10010 14041
rect 9982 14014 10010 14015
rect 9590 13566 9618 13594
rect 8974 13257 9002 13258
rect 8974 13231 8975 13257
rect 8975 13231 9001 13257
rect 9001 13231 9002 13257
rect 8974 13230 9002 13231
rect 9030 13201 9058 13202
rect 9030 13175 9031 13201
rect 9031 13175 9057 13201
rect 9057 13175 9058 13201
rect 9030 13174 9058 13175
rect 6958 12334 6986 12362
rect 2238 12165 2266 12166
rect 2238 12139 2239 12165
rect 2239 12139 2265 12165
rect 2265 12139 2266 12165
rect 2238 12138 2266 12139
rect 2290 12165 2318 12166
rect 2290 12139 2291 12165
rect 2291 12139 2317 12165
rect 2317 12139 2318 12165
rect 2290 12138 2318 12139
rect 2342 12165 2370 12166
rect 2342 12139 2343 12165
rect 2343 12139 2369 12165
rect 2369 12139 2370 12165
rect 2342 12138 2370 12139
rect 6734 11942 6762 11970
rect 6846 11913 6874 11914
rect 6846 11887 6847 11913
rect 6847 11887 6873 11913
rect 6873 11887 6874 11913
rect 6846 11886 6874 11887
rect 7070 12278 7098 12306
rect 7406 12361 7434 12362
rect 7406 12335 7407 12361
rect 7407 12335 7433 12361
rect 7433 12335 7434 12361
rect 7406 12334 7434 12335
rect 7630 12305 7658 12306
rect 7630 12279 7631 12305
rect 7631 12279 7657 12305
rect 7657 12279 7658 12305
rect 7630 12278 7658 12279
rect 7966 12278 7994 12306
rect 7070 11942 7098 11970
rect 2238 11381 2266 11382
rect 2238 11355 2239 11381
rect 2239 11355 2265 11381
rect 2265 11355 2266 11381
rect 2238 11354 2266 11355
rect 2290 11381 2318 11382
rect 2290 11355 2291 11381
rect 2291 11355 2317 11381
rect 2317 11355 2318 11381
rect 2290 11354 2318 11355
rect 2342 11381 2370 11382
rect 2342 11355 2343 11381
rect 2343 11355 2369 11381
rect 2369 11355 2370 11381
rect 2342 11354 2370 11355
rect 6398 10905 6426 10906
rect 6398 10879 6399 10905
rect 6399 10879 6425 10905
rect 6425 10879 6426 10905
rect 6398 10878 6426 10879
rect 4998 10822 5026 10850
rect 2142 10793 2170 10794
rect 2142 10767 2143 10793
rect 2143 10767 2169 10793
rect 2169 10767 2170 10793
rect 2142 10766 2170 10767
rect 2238 10597 2266 10598
rect 2238 10571 2239 10597
rect 2239 10571 2265 10597
rect 2265 10571 2266 10597
rect 2238 10570 2266 10571
rect 2290 10597 2318 10598
rect 2290 10571 2291 10597
rect 2291 10571 2317 10597
rect 2317 10571 2318 10597
rect 2290 10570 2318 10571
rect 2342 10597 2370 10598
rect 2342 10571 2343 10597
rect 2343 10571 2369 10597
rect 2369 10571 2370 10597
rect 2342 10570 2370 10571
rect 6510 10849 6538 10850
rect 6510 10823 6511 10849
rect 6511 10823 6537 10849
rect 6537 10823 6538 10849
rect 6510 10822 6538 10823
rect 6566 10793 6594 10794
rect 6566 10767 6567 10793
rect 6567 10767 6593 10793
rect 6593 10767 6594 10793
rect 6566 10766 6594 10767
rect 6062 10654 6090 10682
rect 2142 10401 2170 10402
rect 2142 10375 2143 10401
rect 2143 10375 2169 10401
rect 2169 10375 2170 10401
rect 2142 10374 2170 10375
rect 6454 10401 6482 10402
rect 6454 10375 6455 10401
rect 6455 10375 6481 10401
rect 6481 10375 6482 10401
rect 6454 10374 6482 10375
rect 7070 11521 7098 11522
rect 7070 11495 7071 11521
rect 7071 11495 7097 11521
rect 7097 11495 7098 11521
rect 7070 11494 7098 11495
rect 6790 10905 6818 10906
rect 6790 10879 6791 10905
rect 6791 10879 6817 10905
rect 6817 10879 6818 10905
rect 6790 10878 6818 10879
rect 6790 10681 6818 10682
rect 6790 10655 6791 10681
rect 6791 10655 6817 10681
rect 6817 10655 6818 10681
rect 6790 10654 6818 10655
rect 6846 10486 6874 10514
rect 6958 10766 6986 10794
rect 8750 12278 8778 12306
rect 8470 11998 8498 12026
rect 7686 11718 7714 11746
rect 8134 11550 8162 11578
rect 7966 11494 7994 11522
rect 8302 11662 8330 11690
rect 8358 11577 8386 11578
rect 8358 11551 8359 11577
rect 8359 11551 8385 11577
rect 8385 11551 8386 11577
rect 8358 11550 8386 11551
rect 8414 11465 8442 11466
rect 8414 11439 8415 11465
rect 8415 11439 8441 11465
rect 8441 11439 8442 11465
rect 8414 11438 8442 11439
rect 9030 11998 9058 12026
rect 8750 11689 8778 11690
rect 8750 11663 8751 11689
rect 8751 11663 8777 11689
rect 8777 11663 8778 11689
rect 8750 11662 8778 11663
rect 7686 11185 7714 11186
rect 7686 11159 7687 11185
rect 7687 11159 7713 11185
rect 7713 11159 7714 11185
rect 7686 11158 7714 11159
rect 8134 11158 8162 11186
rect 7910 11073 7938 11074
rect 7910 11047 7911 11073
rect 7911 11047 7937 11073
rect 7937 11047 7938 11073
rect 7910 11046 7938 11047
rect 8022 10990 8050 11018
rect 8246 11046 8274 11074
rect 7126 10766 7154 10794
rect 8302 10793 8330 10794
rect 8302 10767 8303 10793
rect 8303 10767 8329 10793
rect 8329 10767 8330 10793
rect 8302 10766 8330 10767
rect 6734 10374 6762 10402
rect 2086 9926 2114 9954
rect 5502 10206 5530 10234
rect 6566 10094 6594 10122
rect 2238 9813 2266 9814
rect 2238 9787 2239 9813
rect 2239 9787 2265 9813
rect 2265 9787 2266 9813
rect 2238 9786 2266 9787
rect 2290 9813 2318 9814
rect 2290 9787 2291 9813
rect 2291 9787 2317 9813
rect 2317 9787 2318 9813
rect 2290 9786 2318 9787
rect 2342 9813 2370 9814
rect 2342 9787 2343 9813
rect 2343 9787 2369 9813
rect 2369 9787 2370 9813
rect 2342 9786 2370 9787
rect 6622 9281 6650 9282
rect 6622 9255 6623 9281
rect 6623 9255 6649 9281
rect 6649 9255 6650 9281
rect 6622 9254 6650 9255
rect 5558 9169 5586 9170
rect 5558 9143 5559 9169
rect 5559 9143 5585 9169
rect 5585 9143 5586 9169
rect 5558 9142 5586 9143
rect 2238 9029 2266 9030
rect 2238 9003 2239 9029
rect 2239 9003 2265 9029
rect 2265 9003 2266 9029
rect 2238 9002 2266 9003
rect 2290 9029 2318 9030
rect 2290 9003 2291 9029
rect 2291 9003 2317 9029
rect 2317 9003 2318 9029
rect 2290 9002 2318 9003
rect 2342 9029 2370 9030
rect 2342 9003 2343 9029
rect 2343 9003 2369 9029
rect 2369 9003 2370 9029
rect 2342 9002 2370 9003
rect 6734 8889 6762 8890
rect 6734 8863 6735 8889
rect 6735 8863 6761 8889
rect 6761 8863 6762 8889
rect 6734 8862 6762 8863
rect 2238 8245 2266 8246
rect 2238 8219 2239 8245
rect 2239 8219 2265 8245
rect 2265 8219 2266 8245
rect 2238 8218 2266 8219
rect 2290 8245 2318 8246
rect 2290 8219 2291 8245
rect 2291 8219 2317 8245
rect 2317 8219 2318 8245
rect 2290 8218 2318 8219
rect 2342 8245 2370 8246
rect 2342 8219 2343 8245
rect 2343 8219 2369 8245
rect 2369 8219 2370 8245
rect 2342 8218 2370 8219
rect 2142 8049 2170 8050
rect 2142 8023 2143 8049
rect 2143 8023 2169 8049
rect 2169 8023 2170 8049
rect 2142 8022 2170 8023
rect 5222 8022 5250 8050
rect 966 7742 994 7770
rect 7070 10374 7098 10402
rect 6958 10262 6986 10290
rect 7070 10289 7098 10290
rect 7070 10263 7071 10289
rect 7071 10263 7097 10289
rect 7097 10263 7098 10289
rect 7070 10262 7098 10263
rect 7014 10206 7042 10234
rect 7126 10150 7154 10178
rect 7462 10262 7490 10290
rect 7406 10094 7434 10122
rect 9198 11830 9226 11858
rect 11158 18353 11186 18354
rect 11158 18327 11159 18353
rect 11159 18327 11185 18353
rect 11185 18327 11186 18353
rect 11158 18326 11186 18327
rect 10654 18241 10682 18242
rect 10654 18215 10655 18241
rect 10655 18215 10681 18241
rect 10681 18215 10682 18241
rect 10654 18214 10682 18215
rect 10542 14014 10570 14042
rect 10374 13510 10402 13538
rect 9918 13341 9946 13342
rect 9918 13315 9919 13341
rect 9919 13315 9945 13341
rect 9945 13315 9946 13341
rect 9918 13314 9946 13315
rect 9970 13341 9998 13342
rect 9970 13315 9971 13341
rect 9971 13315 9997 13341
rect 9997 13315 9998 13341
rect 9970 13314 9998 13315
rect 10022 13341 10050 13342
rect 10022 13315 10023 13341
rect 10023 13315 10049 13341
rect 10049 13315 10050 13341
rect 10022 13314 10050 13315
rect 11102 13846 11130 13874
rect 11606 13873 11634 13874
rect 11606 13847 11607 13873
rect 11607 13847 11633 13873
rect 11633 13847 11634 13873
rect 11606 13846 11634 13847
rect 11158 13537 11186 13538
rect 11158 13511 11159 13537
rect 11159 13511 11185 13537
rect 11185 13511 11186 13537
rect 11158 13510 11186 13511
rect 10766 13174 10794 13202
rect 10094 12726 10122 12754
rect 9918 12557 9946 12558
rect 9918 12531 9919 12557
rect 9919 12531 9945 12557
rect 9945 12531 9946 12557
rect 9918 12530 9946 12531
rect 9970 12557 9998 12558
rect 9970 12531 9971 12557
rect 9971 12531 9997 12557
rect 9997 12531 9998 12557
rect 9970 12530 9998 12531
rect 10022 12557 10050 12558
rect 10022 12531 10023 12557
rect 10023 12531 10049 12557
rect 10049 12531 10050 12557
rect 10022 12530 10050 12531
rect 9702 12334 9730 12362
rect 9310 11998 9338 12026
rect 8806 11214 8834 11242
rect 9030 11438 9058 11466
rect 9030 11185 9058 11186
rect 9030 11159 9031 11185
rect 9031 11159 9057 11185
rect 9057 11159 9058 11185
rect 9030 11158 9058 11159
rect 8694 11073 8722 11074
rect 8694 11047 8695 11073
rect 8695 11047 8721 11073
rect 8721 11047 8722 11073
rect 8694 11046 8722 11047
rect 8470 10990 8498 11018
rect 8862 10990 8890 11018
rect 8470 10710 8498 10738
rect 8862 10766 8890 10794
rect 8806 10486 8834 10514
rect 7798 10150 7826 10178
rect 7238 9590 7266 9618
rect 8414 10065 8442 10066
rect 8414 10039 8415 10065
rect 8415 10039 8441 10065
rect 8441 10039 8442 10065
rect 8414 10038 8442 10039
rect 8806 10009 8834 10010
rect 8806 9983 8807 10009
rect 8807 9983 8833 10009
rect 8833 9983 8834 10009
rect 8806 9982 8834 9983
rect 8806 9646 8834 9674
rect 8918 10318 8946 10346
rect 9142 11577 9170 11578
rect 9142 11551 9143 11577
rect 9143 11551 9169 11577
rect 9169 11551 9170 11577
rect 9142 11550 9170 11551
rect 9254 11270 9282 11298
rect 9198 11129 9226 11130
rect 9198 11103 9199 11129
rect 9199 11103 9225 11129
rect 9225 11103 9226 11129
rect 9198 11102 9226 11103
rect 9142 10793 9170 10794
rect 9142 10767 9143 10793
rect 9143 10767 9169 10793
rect 9169 10767 9170 10793
rect 9142 10766 9170 10767
rect 9030 10430 9058 10458
rect 9142 10654 9170 10682
rect 9030 10262 9058 10290
rect 8918 10094 8946 10122
rect 5222 7910 5250 7938
rect 6790 7937 6818 7938
rect 6790 7911 6791 7937
rect 6791 7911 6817 7937
rect 6817 7911 6818 7937
rect 6790 7910 6818 7911
rect 6902 7713 6930 7714
rect 6902 7687 6903 7713
rect 6903 7687 6929 7713
rect 6929 7687 6930 7713
rect 6902 7686 6930 7687
rect 6286 7657 6314 7658
rect 6286 7631 6287 7657
rect 6287 7631 6313 7657
rect 6313 7631 6314 7657
rect 6286 7630 6314 7631
rect 2238 7461 2266 7462
rect 2238 7435 2239 7461
rect 2239 7435 2265 7461
rect 2265 7435 2266 7461
rect 2238 7434 2266 7435
rect 2290 7461 2318 7462
rect 2290 7435 2291 7461
rect 2291 7435 2317 7461
rect 2317 7435 2318 7461
rect 2290 7434 2318 7435
rect 2342 7461 2370 7462
rect 2342 7435 2343 7461
rect 2343 7435 2369 7461
rect 2369 7435 2370 7461
rect 2342 7434 2370 7435
rect 7014 7657 7042 7658
rect 7014 7631 7015 7657
rect 7015 7631 7041 7657
rect 7041 7631 7042 7657
rect 7014 7630 7042 7631
rect 7462 9142 7490 9170
rect 7630 9142 7658 9170
rect 7574 8862 7602 8890
rect 7966 9505 7994 9506
rect 7966 9479 7967 9505
rect 7967 9479 7993 9505
rect 7993 9479 7994 9505
rect 7966 9478 7994 9479
rect 8078 9505 8106 9506
rect 8078 9479 8079 9505
rect 8079 9479 8105 9505
rect 8105 9479 8106 9505
rect 8078 9478 8106 9479
rect 8078 9254 8106 9282
rect 8190 9254 8218 9282
rect 9030 10094 9058 10122
rect 9086 10065 9114 10066
rect 9086 10039 9087 10065
rect 9087 10039 9113 10065
rect 9113 10039 9114 10065
rect 9086 10038 9114 10039
rect 8974 9478 9002 9506
rect 8246 9225 8274 9226
rect 8246 9199 8247 9225
rect 8247 9199 8273 9225
rect 8273 9199 8274 9225
rect 8246 9198 8274 9199
rect 8526 9198 8554 9226
rect 8134 9142 8162 9170
rect 8694 9225 8722 9226
rect 8694 9199 8695 9225
rect 8695 9199 8721 9225
rect 8721 9199 8722 9225
rect 8694 9198 8722 9199
rect 8862 9086 8890 9114
rect 9086 9142 9114 9170
rect 8526 8862 8554 8890
rect 8694 8806 8722 8834
rect 9366 11185 9394 11186
rect 9366 11159 9367 11185
rect 9367 11159 9393 11185
rect 9393 11159 9394 11185
rect 9366 11158 9394 11159
rect 10766 13089 10794 13090
rect 10766 13063 10767 13089
rect 10767 13063 10793 13089
rect 10793 13063 10794 13089
rect 10766 13062 10794 13063
rect 10654 12753 10682 12754
rect 10654 12727 10655 12753
rect 10655 12727 10681 12753
rect 10681 12727 10682 12753
rect 10654 12726 10682 12727
rect 10822 12473 10850 12474
rect 10822 12447 10823 12473
rect 10823 12447 10849 12473
rect 10849 12447 10850 12473
rect 10822 12446 10850 12447
rect 10486 12334 10514 12362
rect 10766 12361 10794 12362
rect 10766 12335 10767 12361
rect 10767 12335 10793 12361
rect 10793 12335 10794 12361
rect 10766 12334 10794 12335
rect 9926 12278 9954 12306
rect 10822 12249 10850 12250
rect 10822 12223 10823 12249
rect 10823 12223 10849 12249
rect 10849 12223 10850 12249
rect 10822 12222 10850 12223
rect 11830 13062 11858 13090
rect 12054 13089 12082 13090
rect 12054 13063 12055 13089
rect 12055 13063 12081 13089
rect 12081 13063 12082 13089
rect 12054 13062 12082 13063
rect 12054 12782 12082 12810
rect 17598 19221 17626 19222
rect 17598 19195 17599 19221
rect 17599 19195 17625 19221
rect 17625 19195 17626 19221
rect 17598 19194 17626 19195
rect 17650 19221 17678 19222
rect 17650 19195 17651 19221
rect 17651 19195 17677 19221
rect 17677 19195 17678 19221
rect 17650 19194 17678 19195
rect 17702 19221 17730 19222
rect 17702 19195 17703 19221
rect 17703 19195 17729 19221
rect 17729 19195 17730 19221
rect 17702 19194 17730 19195
rect 13454 18718 13482 18746
rect 14070 18745 14098 18746
rect 14070 18719 14071 18745
rect 14071 18719 14097 18745
rect 14097 18719 14098 18745
rect 14070 18718 14098 18719
rect 17598 18437 17626 18438
rect 17598 18411 17599 18437
rect 17599 18411 17625 18437
rect 17625 18411 17626 18437
rect 17598 18410 17626 18411
rect 17650 18437 17678 18438
rect 17650 18411 17651 18437
rect 17651 18411 17677 18437
rect 17677 18411 17678 18437
rect 17650 18410 17678 18411
rect 17702 18437 17730 18438
rect 17702 18411 17703 18437
rect 17703 18411 17729 18437
rect 17729 18411 17730 18437
rect 17702 18410 17730 18411
rect 17598 17653 17626 17654
rect 17598 17627 17599 17653
rect 17599 17627 17625 17653
rect 17625 17627 17626 17653
rect 17598 17626 17626 17627
rect 17650 17653 17678 17654
rect 17650 17627 17651 17653
rect 17651 17627 17677 17653
rect 17677 17627 17678 17653
rect 17650 17626 17678 17627
rect 17702 17653 17730 17654
rect 17702 17627 17703 17653
rect 17703 17627 17729 17653
rect 17729 17627 17730 17653
rect 17702 17626 17730 17627
rect 17598 16869 17626 16870
rect 17598 16843 17599 16869
rect 17599 16843 17625 16869
rect 17625 16843 17626 16869
rect 17598 16842 17626 16843
rect 17650 16869 17678 16870
rect 17650 16843 17651 16869
rect 17651 16843 17677 16869
rect 17677 16843 17678 16869
rect 17650 16842 17678 16843
rect 17702 16869 17730 16870
rect 17702 16843 17703 16869
rect 17703 16843 17729 16869
rect 17729 16843 17730 16869
rect 17702 16842 17730 16843
rect 17598 16085 17626 16086
rect 17598 16059 17599 16085
rect 17599 16059 17625 16085
rect 17625 16059 17626 16085
rect 17598 16058 17626 16059
rect 17650 16085 17678 16086
rect 17650 16059 17651 16085
rect 17651 16059 17677 16085
rect 17677 16059 17678 16085
rect 17650 16058 17678 16059
rect 17702 16085 17730 16086
rect 17702 16059 17703 16085
rect 17703 16059 17729 16085
rect 17729 16059 17730 16085
rect 17702 16058 17730 16059
rect 12950 14041 12978 14042
rect 12950 14015 12951 14041
rect 12951 14015 12977 14041
rect 12977 14015 12978 14041
rect 12950 14014 12978 14015
rect 17598 15301 17626 15302
rect 17598 15275 17599 15301
rect 17599 15275 17625 15301
rect 17625 15275 17626 15301
rect 17598 15274 17626 15275
rect 17650 15301 17678 15302
rect 17650 15275 17651 15301
rect 17651 15275 17677 15301
rect 17677 15275 17678 15301
rect 17650 15274 17678 15275
rect 17702 15301 17730 15302
rect 17702 15275 17703 15301
rect 17703 15275 17729 15301
rect 17729 15275 17730 15301
rect 17702 15274 17730 15275
rect 17598 14517 17626 14518
rect 17598 14491 17599 14517
rect 17599 14491 17625 14517
rect 17625 14491 17626 14517
rect 17598 14490 17626 14491
rect 17650 14517 17678 14518
rect 17650 14491 17651 14517
rect 17651 14491 17677 14517
rect 17677 14491 17678 14517
rect 17650 14490 17678 14491
rect 17702 14517 17730 14518
rect 17702 14491 17703 14517
rect 17703 14491 17729 14517
rect 17729 14491 17730 14517
rect 17702 14490 17730 14491
rect 13454 14014 13482 14042
rect 12278 13846 12306 13874
rect 12334 13790 12362 13818
rect 9926 11830 9954 11858
rect 9918 11773 9946 11774
rect 9918 11747 9919 11773
rect 9919 11747 9945 11773
rect 9945 11747 9946 11773
rect 9918 11746 9946 11747
rect 9970 11773 9998 11774
rect 9970 11747 9971 11773
rect 9971 11747 9997 11773
rect 9997 11747 9998 11773
rect 9970 11746 9998 11747
rect 10022 11773 10050 11774
rect 10022 11747 10023 11773
rect 10023 11747 10049 11773
rect 10049 11747 10050 11773
rect 10022 11746 10050 11747
rect 9534 11270 9562 11298
rect 9646 11662 9674 11690
rect 9478 11046 9506 11074
rect 9534 10990 9562 11018
rect 9478 10766 9506 10794
rect 9310 10318 9338 10346
rect 9366 10430 9394 10458
rect 9702 11073 9730 11074
rect 9702 11047 9703 11073
rect 9703 11047 9729 11073
rect 9729 11047 9730 11073
rect 9702 11046 9730 11047
rect 9590 10766 9618 10794
rect 9646 10878 9674 10906
rect 9702 10654 9730 10682
rect 9534 10513 9562 10514
rect 9534 10487 9535 10513
rect 9535 10487 9561 10513
rect 9561 10487 9562 10513
rect 9534 10486 9562 10487
rect 9646 10486 9674 10514
rect 9366 10094 9394 10122
rect 9310 10009 9338 10010
rect 9310 9983 9311 10009
rect 9311 9983 9337 10009
rect 9337 9983 9338 10009
rect 9310 9982 9338 9983
rect 9198 8918 9226 8946
rect 9366 9561 9394 9562
rect 9366 9535 9367 9561
rect 9367 9535 9393 9561
rect 9393 9535 9394 9561
rect 9366 9534 9394 9535
rect 9422 10262 9450 10290
rect 9590 10150 9618 10178
rect 9702 10094 9730 10122
rect 10318 11185 10346 11186
rect 10318 11159 10319 11185
rect 10319 11159 10345 11185
rect 10345 11159 10346 11185
rect 10318 11158 10346 11159
rect 10094 11102 10122 11130
rect 9918 10989 9946 10990
rect 9918 10963 9919 10989
rect 9919 10963 9945 10989
rect 9945 10963 9946 10989
rect 9918 10962 9946 10963
rect 9970 10989 9998 10990
rect 9970 10963 9971 10989
rect 9971 10963 9997 10989
rect 9997 10963 9998 10989
rect 9970 10962 9998 10963
rect 10022 10989 10050 10990
rect 10022 10963 10023 10989
rect 10023 10963 10049 10989
rect 10049 10963 10050 10989
rect 10022 10962 10050 10963
rect 9870 10878 9898 10906
rect 10654 11129 10682 11130
rect 10654 11103 10655 11129
rect 10655 11103 10681 11129
rect 10681 11103 10682 11129
rect 10654 11102 10682 11103
rect 10710 11046 10738 11074
rect 10318 10849 10346 10850
rect 10318 10823 10319 10849
rect 10319 10823 10345 10849
rect 10345 10823 10346 10849
rect 10318 10822 10346 10823
rect 10710 10822 10738 10850
rect 9870 10766 9898 10794
rect 9814 10486 9842 10514
rect 10038 10654 10066 10682
rect 10206 10766 10234 10794
rect 10430 10374 10458 10402
rect 10710 10318 10738 10346
rect 9926 10262 9954 10290
rect 10374 10289 10402 10290
rect 10374 10263 10375 10289
rect 10375 10263 10401 10289
rect 10401 10263 10402 10289
rect 10374 10262 10402 10263
rect 10542 10262 10570 10290
rect 9814 10206 9842 10234
rect 9918 10205 9946 10206
rect 9918 10179 9919 10205
rect 9919 10179 9945 10205
rect 9945 10179 9946 10205
rect 9918 10178 9946 10179
rect 9970 10205 9998 10206
rect 9970 10179 9971 10205
rect 9971 10179 9997 10205
rect 9997 10179 9998 10205
rect 9970 10178 9998 10179
rect 10022 10205 10050 10206
rect 10022 10179 10023 10205
rect 10023 10179 10049 10205
rect 10049 10179 10050 10205
rect 10022 10178 10050 10179
rect 10038 10094 10066 10122
rect 9814 9926 9842 9954
rect 9590 9561 9618 9562
rect 9590 9535 9591 9561
rect 9591 9535 9617 9561
rect 9617 9535 9618 9561
rect 9590 9534 9618 9535
rect 9254 8806 9282 8834
rect 9030 8721 9058 8722
rect 9030 8695 9031 8721
rect 9031 8695 9057 8721
rect 9057 8695 9058 8721
rect 9030 8694 9058 8695
rect 7630 7574 7658 7602
rect 6902 7238 6930 7266
rect 7182 7238 7210 7266
rect 8078 7265 8106 7266
rect 8078 7239 8079 7265
rect 8079 7239 8105 7265
rect 8105 7239 8106 7265
rect 8078 7238 8106 7239
rect 8302 7657 8330 7658
rect 8302 7631 8303 7657
rect 8303 7631 8329 7657
rect 8329 7631 8330 7657
rect 8302 7630 8330 7631
rect 9310 7966 9338 7994
rect 9254 7630 9282 7658
rect 8302 7238 8330 7266
rect 8750 7238 8778 7266
rect 8414 7209 8442 7210
rect 8414 7183 8415 7209
rect 8415 7183 8441 7209
rect 8441 7183 8442 7209
rect 8414 7182 8442 7183
rect 9086 7182 9114 7210
rect 9142 6929 9170 6930
rect 9142 6903 9143 6929
rect 9143 6903 9169 6929
rect 9169 6903 9170 6929
rect 9142 6902 9170 6903
rect 9422 9169 9450 9170
rect 9422 9143 9423 9169
rect 9423 9143 9449 9169
rect 9449 9143 9450 9169
rect 9422 9142 9450 9143
rect 9422 8918 9450 8946
rect 9646 9310 9674 9338
rect 9758 9478 9786 9506
rect 9534 8974 9562 9002
rect 9646 9198 9674 9226
rect 9534 8862 9562 8890
rect 9590 8833 9618 8834
rect 9590 8807 9591 8833
rect 9591 8807 9617 8833
rect 9617 8807 9618 8833
rect 9590 8806 9618 8807
rect 9646 8694 9674 8722
rect 9926 9561 9954 9562
rect 9926 9535 9927 9561
rect 9927 9535 9953 9561
rect 9953 9535 9954 9561
rect 9926 9534 9954 9535
rect 10318 9953 10346 9954
rect 10318 9927 10319 9953
rect 10319 9927 10345 9953
rect 10345 9927 10346 9953
rect 10318 9926 10346 9927
rect 10374 9814 10402 9842
rect 9918 9421 9946 9422
rect 9918 9395 9919 9421
rect 9919 9395 9945 9421
rect 9945 9395 9946 9421
rect 9918 9394 9946 9395
rect 9970 9421 9998 9422
rect 9970 9395 9971 9421
rect 9971 9395 9997 9421
rect 9997 9395 9998 9421
rect 9970 9394 9998 9395
rect 10022 9421 10050 9422
rect 10022 9395 10023 9421
rect 10023 9395 10049 9421
rect 10049 9395 10050 9421
rect 10022 9394 10050 9395
rect 9870 9310 9898 9338
rect 10206 9310 10234 9338
rect 10318 9534 10346 9562
rect 10150 9225 10178 9226
rect 10150 9199 10151 9225
rect 10151 9199 10177 9225
rect 10177 9199 10178 9225
rect 10150 9198 10178 9199
rect 10262 9225 10290 9226
rect 10262 9199 10263 9225
rect 10263 9199 10289 9225
rect 10289 9199 10290 9225
rect 10262 9198 10290 9199
rect 9982 9113 10010 9114
rect 9982 9087 9983 9113
rect 9983 9087 10009 9113
rect 10009 9087 10010 9113
rect 9982 9086 10010 9087
rect 9926 9030 9954 9058
rect 9870 8918 9898 8946
rect 10374 9254 10402 9282
rect 9918 8637 9946 8638
rect 9918 8611 9919 8637
rect 9919 8611 9945 8637
rect 9945 8611 9946 8637
rect 9918 8610 9946 8611
rect 9970 8637 9998 8638
rect 9970 8611 9971 8637
rect 9971 8611 9997 8637
rect 9997 8611 9998 8637
rect 9970 8610 9998 8611
rect 10022 8637 10050 8638
rect 10022 8611 10023 8637
rect 10023 8611 10049 8637
rect 10049 8611 10050 8637
rect 10022 8610 10050 8611
rect 10710 10206 10738 10234
rect 10598 9310 10626 9338
rect 10542 9169 10570 9170
rect 10542 9143 10543 9169
rect 10543 9143 10569 9169
rect 10569 9143 10570 9169
rect 10542 9142 10570 9143
rect 10654 8974 10682 9002
rect 10710 8889 10738 8890
rect 10710 8863 10711 8889
rect 10711 8863 10737 8889
rect 10737 8863 10738 8889
rect 10710 8862 10738 8863
rect 10934 11718 10962 11746
rect 10878 11046 10906 11074
rect 10934 10878 10962 10906
rect 10822 10849 10850 10850
rect 10822 10823 10823 10849
rect 10823 10823 10849 10849
rect 10849 10823 10850 10849
rect 10822 10822 10850 10823
rect 10934 10401 10962 10402
rect 10934 10375 10935 10401
rect 10935 10375 10961 10401
rect 10961 10375 10962 10401
rect 10934 10374 10962 10375
rect 9758 7993 9786 7994
rect 9758 7967 9759 7993
rect 9759 7967 9785 7993
rect 9785 7967 9786 7993
rect 9758 7966 9786 7967
rect 10430 8302 10458 8330
rect 9926 8049 9954 8050
rect 9926 8023 9927 8049
rect 9927 8023 9953 8049
rect 9953 8023 9954 8049
rect 9926 8022 9954 8023
rect 10654 8694 10682 8722
rect 9918 7853 9946 7854
rect 9918 7827 9919 7853
rect 9919 7827 9945 7853
rect 9945 7827 9946 7853
rect 9918 7826 9946 7827
rect 9970 7853 9998 7854
rect 9970 7827 9971 7853
rect 9971 7827 9997 7853
rect 9997 7827 9998 7853
rect 9970 7826 9998 7827
rect 10022 7853 10050 7854
rect 10022 7827 10023 7853
rect 10023 7827 10049 7853
rect 10049 7827 10050 7853
rect 10022 7826 10050 7827
rect 9814 7630 9842 7658
rect 10430 7769 10458 7770
rect 10430 7743 10431 7769
rect 10431 7743 10457 7769
rect 10457 7743 10458 7769
rect 10430 7742 10458 7743
rect 10710 8049 10738 8050
rect 10710 8023 10711 8049
rect 10711 8023 10737 8049
rect 10737 8023 10738 8049
rect 10710 8022 10738 8023
rect 10878 8833 10906 8834
rect 10878 8807 10879 8833
rect 10879 8807 10905 8833
rect 10905 8807 10906 8833
rect 10878 8806 10906 8807
rect 12110 12446 12138 12474
rect 11102 12222 11130 12250
rect 12950 13817 12978 13818
rect 12950 13791 12951 13817
rect 12951 13791 12977 13817
rect 12977 13791 12978 13817
rect 12950 13790 12978 13791
rect 17598 13733 17626 13734
rect 17598 13707 17599 13733
rect 17599 13707 17625 13733
rect 17625 13707 17626 13733
rect 17598 13706 17626 13707
rect 17650 13733 17678 13734
rect 17650 13707 17651 13733
rect 17651 13707 17677 13733
rect 17677 13707 17678 13733
rect 17650 13706 17678 13707
rect 17702 13733 17730 13734
rect 17702 13707 17703 13733
rect 17703 13707 17729 13733
rect 17729 13707 17730 13733
rect 17702 13706 17730 13707
rect 13062 13510 13090 13538
rect 12334 12809 12362 12810
rect 12334 12783 12335 12809
rect 12335 12783 12361 12809
rect 12361 12783 12362 12809
rect 12334 12782 12362 12783
rect 12614 12782 12642 12810
rect 13230 13062 13258 13090
rect 12222 11662 12250 11690
rect 12222 11382 12250 11410
rect 12278 11718 12306 11746
rect 11046 10822 11074 10850
rect 11102 11158 11130 11186
rect 10990 10094 11018 10122
rect 12782 11382 12810 11410
rect 11494 11046 11522 11074
rect 11382 10878 11410 10906
rect 11270 10793 11298 10794
rect 11270 10767 11271 10793
rect 11271 10767 11297 10793
rect 11297 10767 11298 10793
rect 11270 10766 11298 10767
rect 11550 10849 11578 10850
rect 11550 10823 11551 10849
rect 11551 10823 11577 10849
rect 11577 10823 11578 10849
rect 11550 10822 11578 10823
rect 11942 10542 11970 10570
rect 14070 13089 14098 13090
rect 14070 13063 14071 13089
rect 14071 13063 14097 13089
rect 14097 13063 14098 13089
rect 14070 13062 14098 13063
rect 20006 13118 20034 13146
rect 18830 13062 18858 13090
rect 17598 12949 17626 12950
rect 17598 12923 17599 12949
rect 17599 12923 17625 12949
rect 17625 12923 17626 12949
rect 17598 12922 17626 12923
rect 17650 12949 17678 12950
rect 17650 12923 17651 12949
rect 17651 12923 17677 12949
rect 17677 12923 17678 12949
rect 17650 12922 17678 12923
rect 17702 12949 17730 12950
rect 17702 12923 17703 12949
rect 17703 12923 17729 12949
rect 17729 12923 17730 12949
rect 17702 12922 17730 12923
rect 17598 12165 17626 12166
rect 17598 12139 17599 12165
rect 17599 12139 17625 12165
rect 17625 12139 17626 12165
rect 17598 12138 17626 12139
rect 17650 12165 17678 12166
rect 17650 12139 17651 12165
rect 17651 12139 17677 12165
rect 17677 12139 17678 12165
rect 17650 12138 17678 12139
rect 17702 12165 17730 12166
rect 17702 12139 17703 12165
rect 17703 12139 17729 12165
rect 17729 12139 17730 12165
rect 17702 12138 17730 12139
rect 13454 11942 13482 11970
rect 14518 11942 14546 11970
rect 12222 10457 12250 10458
rect 12222 10431 12223 10457
rect 12223 10431 12249 10457
rect 12249 10431 12250 10457
rect 12222 10430 12250 10431
rect 11886 10374 11914 10402
rect 11662 10345 11690 10346
rect 11662 10319 11663 10345
rect 11663 10319 11689 10345
rect 11689 10319 11690 10345
rect 11662 10318 11690 10319
rect 11270 10206 11298 10234
rect 11102 9646 11130 9674
rect 11158 10150 11186 10178
rect 11046 9534 11074 9562
rect 10878 8694 10906 8722
rect 10990 8918 11018 8946
rect 11158 9225 11186 9226
rect 11158 9199 11159 9225
rect 11159 9199 11185 9225
rect 11185 9199 11186 9225
rect 11158 9198 11186 9199
rect 11326 10094 11354 10122
rect 11494 10289 11522 10290
rect 11494 10263 11495 10289
rect 11495 10263 11521 10289
rect 11521 10263 11522 10289
rect 11494 10262 11522 10263
rect 11718 10094 11746 10122
rect 11606 9814 11634 9842
rect 11382 9254 11410 9282
rect 11550 9646 11578 9674
rect 11326 8974 11354 9002
rect 12166 10374 12194 10402
rect 18830 11969 18858 11970
rect 18830 11943 18831 11969
rect 18831 11943 18857 11969
rect 18857 11943 18858 11969
rect 18830 11942 18858 11943
rect 20006 11774 20034 11802
rect 14630 11633 14658 11634
rect 14630 11607 14631 11633
rect 14631 11607 14657 11633
rect 14657 11607 14658 11633
rect 14630 11606 14658 11607
rect 18830 11577 18858 11578
rect 18830 11551 18831 11577
rect 18831 11551 18857 11577
rect 18857 11551 18858 11577
rect 18830 11550 18858 11551
rect 20006 11465 20034 11466
rect 20006 11439 20007 11465
rect 20007 11439 20033 11465
rect 20033 11439 20034 11465
rect 20006 11438 20034 11439
rect 17598 11381 17626 11382
rect 17598 11355 17599 11381
rect 17599 11355 17625 11381
rect 17625 11355 17626 11381
rect 17598 11354 17626 11355
rect 17650 11381 17678 11382
rect 17650 11355 17651 11381
rect 17651 11355 17677 11381
rect 17677 11355 17678 11381
rect 17650 11354 17678 11355
rect 17702 11381 17730 11382
rect 17702 11355 17703 11381
rect 17703 11355 17729 11381
rect 17729 11355 17730 11381
rect 17702 11354 17730 11355
rect 18830 11185 18858 11186
rect 18830 11159 18831 11185
rect 18831 11159 18857 11185
rect 18857 11159 18858 11185
rect 18830 11158 18858 11159
rect 20006 11102 20034 11130
rect 13566 10822 13594 10850
rect 13174 10430 13202 10458
rect 12838 10150 12866 10178
rect 12054 9814 12082 9842
rect 11774 9478 11802 9506
rect 11942 9254 11970 9282
rect 12110 9534 12138 9562
rect 11886 8889 11914 8890
rect 11886 8863 11887 8889
rect 11887 8863 11913 8889
rect 11913 8863 11914 8889
rect 11886 8862 11914 8863
rect 11550 8582 11578 8610
rect 11606 8721 11634 8722
rect 11606 8695 11607 8721
rect 11607 8695 11633 8721
rect 11633 8695 11634 8721
rect 11606 8694 11634 8695
rect 10766 7769 10794 7770
rect 10766 7743 10767 7769
rect 10767 7743 10793 7769
rect 10793 7743 10794 7769
rect 10766 7742 10794 7743
rect 10318 7574 10346 7602
rect 9814 7294 9842 7322
rect 9702 7265 9730 7266
rect 9702 7239 9703 7265
rect 9703 7239 9729 7265
rect 9729 7239 9730 7265
rect 9702 7238 9730 7239
rect 10206 7238 10234 7266
rect 9918 7069 9946 7070
rect 9918 7043 9919 7069
rect 9919 7043 9945 7069
rect 9945 7043 9946 7069
rect 9918 7042 9946 7043
rect 9970 7069 9998 7070
rect 9970 7043 9971 7069
rect 9971 7043 9997 7069
rect 9997 7043 9998 7069
rect 9970 7042 9998 7043
rect 10022 7069 10050 7070
rect 10022 7043 10023 7069
rect 10023 7043 10049 7069
rect 10049 7043 10050 7069
rect 10022 7042 10050 7043
rect 9534 6902 9562 6930
rect 2238 6677 2266 6678
rect 2238 6651 2239 6677
rect 2239 6651 2265 6677
rect 2265 6651 2266 6677
rect 2238 6650 2266 6651
rect 2290 6677 2318 6678
rect 2290 6651 2291 6677
rect 2291 6651 2317 6677
rect 2317 6651 2318 6677
rect 2290 6650 2318 6651
rect 2342 6677 2370 6678
rect 2342 6651 2343 6677
rect 2343 6651 2369 6677
rect 2369 6651 2370 6677
rect 2342 6650 2370 6651
rect 2238 5893 2266 5894
rect 2238 5867 2239 5893
rect 2239 5867 2265 5893
rect 2265 5867 2266 5893
rect 2238 5866 2266 5867
rect 2290 5893 2318 5894
rect 2290 5867 2291 5893
rect 2291 5867 2317 5893
rect 2317 5867 2318 5893
rect 2290 5866 2318 5867
rect 2342 5893 2370 5894
rect 2342 5867 2343 5893
rect 2343 5867 2369 5893
rect 2369 5867 2370 5893
rect 2342 5866 2370 5867
rect 2238 5109 2266 5110
rect 2238 5083 2239 5109
rect 2239 5083 2265 5109
rect 2265 5083 2266 5109
rect 2238 5082 2266 5083
rect 2290 5109 2318 5110
rect 2290 5083 2291 5109
rect 2291 5083 2317 5109
rect 2317 5083 2318 5109
rect 2290 5082 2318 5083
rect 2342 5109 2370 5110
rect 2342 5083 2343 5109
rect 2343 5083 2369 5109
rect 2369 5083 2370 5109
rect 2342 5082 2370 5083
rect 2238 4325 2266 4326
rect 2238 4299 2239 4325
rect 2239 4299 2265 4325
rect 2265 4299 2266 4325
rect 2238 4298 2266 4299
rect 2290 4325 2318 4326
rect 2290 4299 2291 4325
rect 2291 4299 2317 4325
rect 2317 4299 2318 4325
rect 2290 4298 2318 4299
rect 2342 4325 2370 4326
rect 2342 4299 2343 4325
rect 2343 4299 2369 4325
rect 2369 4299 2370 4325
rect 2342 4298 2370 4299
rect 2238 3541 2266 3542
rect 2238 3515 2239 3541
rect 2239 3515 2265 3541
rect 2265 3515 2266 3541
rect 2238 3514 2266 3515
rect 2290 3541 2318 3542
rect 2290 3515 2291 3541
rect 2291 3515 2317 3541
rect 2317 3515 2318 3541
rect 2290 3514 2318 3515
rect 2342 3541 2370 3542
rect 2342 3515 2343 3541
rect 2343 3515 2369 3541
rect 2369 3515 2370 3541
rect 2342 3514 2370 3515
rect 2238 2757 2266 2758
rect 2238 2731 2239 2757
rect 2239 2731 2265 2757
rect 2265 2731 2266 2757
rect 2238 2730 2266 2731
rect 2290 2757 2318 2758
rect 2290 2731 2291 2757
rect 2291 2731 2317 2757
rect 2317 2731 2318 2757
rect 2290 2730 2318 2731
rect 2342 2757 2370 2758
rect 2342 2731 2343 2757
rect 2343 2731 2369 2757
rect 2369 2731 2370 2757
rect 2342 2730 2370 2731
rect 2238 1973 2266 1974
rect 2238 1947 2239 1973
rect 2239 1947 2265 1973
rect 2265 1947 2266 1973
rect 2238 1946 2266 1947
rect 2290 1973 2318 1974
rect 2290 1947 2291 1973
rect 2291 1947 2317 1973
rect 2317 1947 2318 1973
rect 2290 1946 2318 1947
rect 2342 1973 2370 1974
rect 2342 1947 2343 1973
rect 2343 1947 2369 1973
rect 2369 1947 2370 1973
rect 2342 1946 2370 1947
rect 10262 7209 10290 7210
rect 10262 7183 10263 7209
rect 10263 7183 10289 7209
rect 10289 7183 10290 7209
rect 10262 7182 10290 7183
rect 10206 6873 10234 6874
rect 10206 6847 10207 6873
rect 10207 6847 10233 6873
rect 10233 6847 10234 6873
rect 10206 6846 10234 6847
rect 9918 6285 9946 6286
rect 9918 6259 9919 6285
rect 9919 6259 9945 6285
rect 9945 6259 9946 6285
rect 9918 6258 9946 6259
rect 9970 6285 9998 6286
rect 9970 6259 9971 6285
rect 9971 6259 9997 6285
rect 9997 6259 9998 6285
rect 9970 6258 9998 6259
rect 10022 6285 10050 6286
rect 10022 6259 10023 6285
rect 10023 6259 10049 6285
rect 10049 6259 10050 6285
rect 10022 6258 10050 6259
rect 9758 5950 9786 5978
rect 12670 9561 12698 9562
rect 12670 9535 12671 9561
rect 12671 9535 12697 9561
rect 12697 9535 12698 9561
rect 12670 9534 12698 9535
rect 13118 10401 13146 10402
rect 13118 10375 13119 10401
rect 13119 10375 13145 10401
rect 13145 10375 13146 10401
rect 13118 10374 13146 10375
rect 13454 10374 13482 10402
rect 18830 10793 18858 10794
rect 18830 10767 18831 10793
rect 18831 10767 18857 10793
rect 18857 10767 18858 10793
rect 18830 10766 18858 10767
rect 20006 10766 20034 10794
rect 13622 10710 13650 10738
rect 14238 10737 14266 10738
rect 14238 10711 14239 10737
rect 14239 10711 14265 10737
rect 14265 10711 14266 10737
rect 14238 10710 14266 10711
rect 17598 10597 17626 10598
rect 17598 10571 17599 10597
rect 17599 10571 17625 10597
rect 17625 10571 17626 10597
rect 17598 10570 17626 10571
rect 17650 10597 17678 10598
rect 17650 10571 17651 10597
rect 17651 10571 17677 10597
rect 17677 10571 17678 10597
rect 17650 10570 17678 10571
rect 17702 10597 17730 10598
rect 17702 10571 17703 10597
rect 17703 10571 17729 10597
rect 17729 10571 17730 10597
rect 17702 10570 17730 10571
rect 13734 10318 13762 10346
rect 13342 10150 13370 10178
rect 17598 9813 17626 9814
rect 17598 9787 17599 9813
rect 17599 9787 17625 9813
rect 17625 9787 17626 9813
rect 17598 9786 17626 9787
rect 17650 9813 17678 9814
rect 17650 9787 17651 9813
rect 17651 9787 17677 9813
rect 17677 9787 17678 9813
rect 17650 9786 17678 9787
rect 17702 9813 17730 9814
rect 17702 9787 17703 9813
rect 17703 9787 17729 9813
rect 17729 9787 17730 9813
rect 17702 9786 17730 9787
rect 13734 9673 13762 9674
rect 13734 9647 13735 9673
rect 13735 9647 13761 9673
rect 13761 9647 13762 9673
rect 13734 9646 13762 9647
rect 20006 9758 20034 9786
rect 18830 9646 18858 9674
rect 12894 9030 12922 9058
rect 17598 9029 17626 9030
rect 17598 9003 17599 9029
rect 17599 9003 17625 9029
rect 17625 9003 17626 9029
rect 17598 9002 17626 9003
rect 17650 9029 17678 9030
rect 17650 9003 17651 9029
rect 17651 9003 17677 9029
rect 17677 9003 17678 9029
rect 17650 9002 17678 9003
rect 17702 9029 17730 9030
rect 17702 9003 17703 9029
rect 17703 9003 17729 9029
rect 17729 9003 17730 9029
rect 17702 9002 17730 9003
rect 12054 8777 12082 8778
rect 12054 8751 12055 8777
rect 12055 8751 12081 8777
rect 12081 8751 12082 8777
rect 12054 8750 12082 8751
rect 12614 8777 12642 8778
rect 12614 8751 12615 8777
rect 12615 8751 12641 8777
rect 12641 8751 12642 8777
rect 12614 8750 12642 8751
rect 12222 8694 12250 8722
rect 12782 8638 12810 8666
rect 11830 8358 11858 8386
rect 12222 8582 12250 8610
rect 14014 8721 14042 8722
rect 14014 8695 14015 8721
rect 14015 8695 14041 8721
rect 14041 8695 14042 8721
rect 14014 8694 14042 8695
rect 13902 8638 13930 8666
rect 20006 8750 20034 8778
rect 18830 8638 18858 8666
rect 18942 8694 18970 8722
rect 20006 8414 20034 8442
rect 12670 8385 12698 8386
rect 12670 8359 12671 8385
rect 12671 8359 12697 8385
rect 12697 8359 12698 8385
rect 12670 8358 12698 8359
rect 12614 8329 12642 8330
rect 12614 8303 12615 8329
rect 12615 8303 12641 8329
rect 12641 8303 12642 8329
rect 12614 8302 12642 8303
rect 17598 8245 17626 8246
rect 17598 8219 17599 8245
rect 17599 8219 17625 8245
rect 17625 8219 17626 8245
rect 17598 8218 17626 8219
rect 17650 8245 17678 8246
rect 17650 8219 17651 8245
rect 17651 8219 17677 8245
rect 17677 8219 17678 8245
rect 17650 8218 17678 8219
rect 17702 8245 17730 8246
rect 17702 8219 17703 8245
rect 17703 8219 17729 8245
rect 17729 8219 17730 8245
rect 17702 8218 17730 8219
rect 12334 7686 12362 7714
rect 12614 7686 12642 7714
rect 11102 7209 11130 7210
rect 11102 7183 11103 7209
rect 11103 7183 11129 7209
rect 11129 7183 11130 7209
rect 11102 7182 11130 7183
rect 11158 6734 11186 6762
rect 11438 6846 11466 6874
rect 11606 6734 11634 6762
rect 12278 6734 12306 6762
rect 10318 5950 10346 5978
rect 10710 5950 10738 5978
rect 9918 5501 9946 5502
rect 9918 5475 9919 5501
rect 9919 5475 9945 5501
rect 9945 5475 9946 5501
rect 9918 5474 9946 5475
rect 9970 5501 9998 5502
rect 9970 5475 9971 5501
rect 9971 5475 9997 5501
rect 9997 5475 9998 5501
rect 9970 5474 9998 5475
rect 10022 5501 10050 5502
rect 10022 5475 10023 5501
rect 10023 5475 10049 5501
rect 10049 5475 10050 5501
rect 10022 5474 10050 5475
rect 9918 4717 9946 4718
rect 9918 4691 9919 4717
rect 9919 4691 9945 4717
rect 9945 4691 9946 4717
rect 9918 4690 9946 4691
rect 9970 4717 9998 4718
rect 9970 4691 9971 4717
rect 9971 4691 9997 4717
rect 9997 4691 9998 4717
rect 9970 4690 9998 4691
rect 10022 4717 10050 4718
rect 10022 4691 10023 4717
rect 10023 4691 10049 4717
rect 10049 4691 10050 4717
rect 10022 4690 10050 4691
rect 9918 3933 9946 3934
rect 9918 3907 9919 3933
rect 9919 3907 9945 3933
rect 9945 3907 9946 3933
rect 9918 3906 9946 3907
rect 9970 3933 9998 3934
rect 9970 3907 9971 3933
rect 9971 3907 9997 3933
rect 9997 3907 9998 3933
rect 9970 3906 9998 3907
rect 10022 3933 10050 3934
rect 10022 3907 10023 3933
rect 10023 3907 10049 3933
rect 10049 3907 10050 3933
rect 10022 3906 10050 3907
rect 9918 3149 9946 3150
rect 9918 3123 9919 3149
rect 9919 3123 9945 3149
rect 9945 3123 9946 3149
rect 9918 3122 9946 3123
rect 9970 3149 9998 3150
rect 9970 3123 9971 3149
rect 9971 3123 9997 3149
rect 9997 3123 9998 3149
rect 9970 3122 9998 3123
rect 10022 3149 10050 3150
rect 10022 3123 10023 3149
rect 10023 3123 10049 3149
rect 10049 3123 10050 3149
rect 10022 3122 10050 3123
rect 9918 2365 9946 2366
rect 9918 2339 9919 2365
rect 9919 2339 9945 2365
rect 9945 2339 9946 2365
rect 9918 2338 9946 2339
rect 9970 2365 9998 2366
rect 9970 2339 9971 2365
rect 9971 2339 9997 2365
rect 9997 2339 9998 2365
rect 9970 2338 9998 2339
rect 10022 2365 10050 2366
rect 10022 2339 10023 2365
rect 10023 2339 10049 2365
rect 10049 2339 10050 2365
rect 10022 2338 10050 2339
rect 9422 2030 9450 2058
rect 8414 1694 8442 1722
rect 9030 1694 9058 1722
rect 10038 2057 10066 2058
rect 10038 2031 10039 2057
rect 10039 2031 10065 2057
rect 10065 2031 10066 2057
rect 10038 2030 10066 2031
rect 11438 1806 11466 1834
rect 9918 1581 9946 1582
rect 9918 1555 9919 1581
rect 9919 1555 9945 1581
rect 9945 1555 9946 1581
rect 9918 1554 9946 1555
rect 9970 1581 9998 1582
rect 9970 1555 9971 1581
rect 9971 1555 9997 1581
rect 9997 1555 9998 1581
rect 9970 1554 9998 1555
rect 10022 1581 10050 1582
rect 10022 1555 10023 1581
rect 10023 1555 10049 1581
rect 10049 1555 10050 1581
rect 10022 1554 10050 1555
rect 13286 7686 13314 7714
rect 17598 7461 17626 7462
rect 17598 7435 17599 7461
rect 17599 7435 17625 7461
rect 17625 7435 17626 7461
rect 17598 7434 17626 7435
rect 17650 7461 17678 7462
rect 17650 7435 17651 7461
rect 17651 7435 17677 7461
rect 17677 7435 17678 7461
rect 17650 7434 17678 7435
rect 17702 7461 17730 7462
rect 17702 7435 17703 7461
rect 17703 7435 17729 7461
rect 17729 7435 17730 7461
rect 17702 7434 17730 7435
rect 17598 6677 17626 6678
rect 17598 6651 17599 6677
rect 17599 6651 17625 6677
rect 17625 6651 17626 6677
rect 17598 6650 17626 6651
rect 17650 6677 17678 6678
rect 17650 6651 17651 6677
rect 17651 6651 17677 6677
rect 17677 6651 17678 6677
rect 17650 6650 17678 6651
rect 17702 6677 17730 6678
rect 17702 6651 17703 6677
rect 17703 6651 17729 6677
rect 17729 6651 17730 6677
rect 17702 6650 17730 6651
rect 17598 5893 17626 5894
rect 17598 5867 17599 5893
rect 17599 5867 17625 5893
rect 17625 5867 17626 5893
rect 17598 5866 17626 5867
rect 17650 5893 17678 5894
rect 17650 5867 17651 5893
rect 17651 5867 17677 5893
rect 17677 5867 17678 5893
rect 17650 5866 17678 5867
rect 17702 5893 17730 5894
rect 17702 5867 17703 5893
rect 17703 5867 17729 5893
rect 17729 5867 17730 5893
rect 17702 5866 17730 5867
rect 17598 5109 17626 5110
rect 17598 5083 17599 5109
rect 17599 5083 17625 5109
rect 17625 5083 17626 5109
rect 17598 5082 17626 5083
rect 17650 5109 17678 5110
rect 17650 5083 17651 5109
rect 17651 5083 17677 5109
rect 17677 5083 17678 5109
rect 17650 5082 17678 5083
rect 17702 5109 17730 5110
rect 17702 5083 17703 5109
rect 17703 5083 17729 5109
rect 17729 5083 17730 5109
rect 17702 5082 17730 5083
rect 17598 4325 17626 4326
rect 17598 4299 17599 4325
rect 17599 4299 17625 4325
rect 17625 4299 17626 4325
rect 17598 4298 17626 4299
rect 17650 4325 17678 4326
rect 17650 4299 17651 4325
rect 17651 4299 17677 4325
rect 17677 4299 17678 4325
rect 17650 4298 17678 4299
rect 17702 4325 17730 4326
rect 17702 4299 17703 4325
rect 17703 4299 17729 4325
rect 17729 4299 17730 4325
rect 17702 4298 17730 4299
rect 17598 3541 17626 3542
rect 17598 3515 17599 3541
rect 17599 3515 17625 3541
rect 17625 3515 17626 3541
rect 17598 3514 17626 3515
rect 17650 3541 17678 3542
rect 17650 3515 17651 3541
rect 17651 3515 17677 3541
rect 17677 3515 17678 3541
rect 17650 3514 17678 3515
rect 17702 3541 17730 3542
rect 17702 3515 17703 3541
rect 17703 3515 17729 3541
rect 17729 3515 17730 3541
rect 17702 3514 17730 3515
rect 17598 2757 17626 2758
rect 17598 2731 17599 2757
rect 17599 2731 17625 2757
rect 17625 2731 17626 2757
rect 17598 2730 17626 2731
rect 17650 2757 17678 2758
rect 17650 2731 17651 2757
rect 17651 2731 17677 2757
rect 17677 2731 17678 2757
rect 17650 2730 17678 2731
rect 17702 2757 17730 2758
rect 17702 2731 17703 2757
rect 17703 2731 17729 2757
rect 17729 2731 17730 2757
rect 17702 2730 17730 2731
rect 12446 2030 12474 2058
rect 13118 2057 13146 2058
rect 13118 2031 13119 2057
rect 13119 2031 13145 2057
rect 13145 2031 13146 2057
rect 13118 2030 13146 2031
rect 17598 1973 17626 1974
rect 17598 1947 17599 1973
rect 17599 1947 17625 1973
rect 17625 1947 17626 1973
rect 17598 1946 17626 1947
rect 17650 1973 17678 1974
rect 17650 1947 17651 1973
rect 17651 1947 17677 1973
rect 17677 1947 17678 1973
rect 17650 1946 17678 1947
rect 17702 1973 17730 1974
rect 17702 1947 17703 1973
rect 17703 1947 17729 1973
rect 17729 1947 17730 1973
rect 17702 1946 17730 1947
rect 12782 1833 12810 1834
rect 12782 1807 12783 1833
rect 12783 1807 12809 1833
rect 12809 1807 12810 1833
rect 12782 1806 12810 1807
<< metal3 >>
rect 2233 19194 2238 19222
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2370 19194 2375 19222
rect 17593 19194 17598 19222
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17730 19194 17735 19222
rect 11433 19110 11438 19138
rect 11466 19110 12782 19138
rect 12810 19110 12815 19138
rect 9913 18802 9918 18830
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 10050 18802 10055 18830
rect 10425 18718 10430 18746
rect 10458 18718 11046 18746
rect 11074 18718 11079 18746
rect 13449 18718 13454 18746
rect 13482 18718 14070 18746
rect 14098 18718 14103 18746
rect 2233 18410 2238 18438
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2370 18410 2375 18438
rect 17593 18410 17598 18438
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17730 18410 17735 18438
rect 10089 18326 10094 18354
rect 10122 18326 11158 18354
rect 11186 18326 11191 18354
rect 10145 18214 10150 18242
rect 10178 18214 10654 18242
rect 10682 18214 10687 18242
rect 0 18186 400 18200
rect 0 18158 854 18186
rect 882 18158 887 18186
rect 0 18144 400 18158
rect 9913 18018 9918 18046
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 10050 18018 10055 18046
rect 2233 17626 2238 17654
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2370 17626 2375 17654
rect 17593 17626 17598 17654
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17730 17626 17735 17654
rect 9913 17234 9918 17262
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 10050 17234 10055 17262
rect 2233 16842 2238 16870
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2370 16842 2375 16870
rect 17593 16842 17598 16870
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17730 16842 17735 16870
rect 9913 16450 9918 16478
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 10050 16450 10055 16478
rect 2233 16058 2238 16086
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2370 16058 2375 16086
rect 17593 16058 17598 16086
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17730 16058 17735 16086
rect 9913 15666 9918 15694
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 10050 15666 10055 15694
rect 2233 15274 2238 15302
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2370 15274 2375 15302
rect 17593 15274 17598 15302
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17730 15274 17735 15302
rect 9913 14882 9918 14910
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 10050 14882 10055 14910
rect 2233 14490 2238 14518
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2370 14490 2375 14518
rect 17593 14490 17598 14518
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17730 14490 17735 14518
rect 9305 14294 9310 14322
rect 9338 14294 10038 14322
rect 10066 14294 10071 14322
rect 9865 14238 9870 14266
rect 9898 14238 10150 14266
rect 10178 14238 10183 14266
rect 9913 14098 9918 14126
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 10050 14098 10055 14126
rect 9977 14014 9982 14042
rect 10010 14014 10542 14042
rect 10570 14014 10575 14042
rect 12945 14014 12950 14042
rect 12978 14014 13454 14042
rect 13482 14014 13487 14042
rect 11097 13846 11102 13874
rect 11130 13846 11606 13874
rect 11634 13846 12278 13874
rect 12306 13846 12311 13874
rect 0 13818 400 13832
rect 0 13790 2086 13818
rect 2114 13790 2119 13818
rect 12329 13790 12334 13818
rect 12362 13790 12950 13818
rect 12978 13790 12983 13818
rect 0 13776 400 13790
rect 2233 13706 2238 13734
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2370 13706 2375 13734
rect 17593 13706 17598 13734
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17730 13706 17735 13734
rect 8633 13566 8638 13594
rect 8666 13566 9590 13594
rect 9618 13566 9623 13594
rect 10369 13510 10374 13538
rect 10402 13510 11158 13538
rect 11186 13510 13062 13538
rect 13090 13510 13095 13538
rect 9913 13314 9918 13342
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 10050 13314 10055 13342
rect 7569 13230 7574 13258
rect 7602 13230 8974 13258
rect 9002 13230 9007 13258
rect 9025 13174 9030 13202
rect 9058 13174 10766 13202
rect 10794 13174 10799 13202
rect 20600 13146 21000 13160
rect 20001 13118 20006 13146
rect 20034 13118 21000 13146
rect 20600 13104 21000 13118
rect 10761 13062 10766 13090
rect 10794 13062 11830 13090
rect 11858 13062 12054 13090
rect 12082 13062 12087 13090
rect 13225 13062 13230 13090
rect 13258 13062 14070 13090
rect 14098 13062 18830 13090
rect 18858 13062 18863 13090
rect 2233 12922 2238 12950
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2370 12922 2375 12950
rect 17593 12922 17598 12950
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17730 12922 17735 12950
rect 12049 12782 12054 12810
rect 12082 12782 12334 12810
rect 12362 12782 12614 12810
rect 12642 12782 12647 12810
rect 10089 12726 10094 12754
rect 10122 12726 10654 12754
rect 10682 12726 10687 12754
rect 9913 12530 9918 12558
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 10050 12530 10055 12558
rect 10817 12446 10822 12474
rect 10850 12446 12110 12474
rect 12138 12446 12143 12474
rect 2137 12334 2142 12362
rect 2170 12334 5614 12362
rect 5642 12334 6958 12362
rect 6986 12334 6991 12362
rect 7401 12334 7406 12362
rect 7434 12334 9702 12362
rect 9730 12334 10486 12362
rect 10514 12334 10766 12362
rect 10794 12334 10799 12362
rect 7065 12278 7070 12306
rect 7098 12278 7630 12306
rect 7658 12278 7966 12306
rect 7994 12278 8750 12306
rect 8778 12278 9926 12306
rect 9954 12278 9959 12306
rect 961 12222 966 12250
rect 994 12222 999 12250
rect 10817 12222 10822 12250
rect 10850 12222 11102 12250
rect 11130 12222 11135 12250
rect 0 12138 400 12152
rect 966 12138 994 12222
rect 2233 12138 2238 12166
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2370 12138 2375 12166
rect 17593 12138 17598 12166
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17730 12138 17735 12166
rect 0 12110 994 12138
rect 0 12096 400 12110
rect 8465 11998 8470 12026
rect 8498 11998 9030 12026
rect 9058 11998 9310 12026
rect 9338 11998 9343 12026
rect 6729 11942 6734 11970
rect 6762 11942 7070 11970
rect 7098 11942 7103 11970
rect 13449 11942 13454 11970
rect 13482 11942 14518 11970
rect 14546 11942 18830 11970
rect 18858 11942 18863 11970
rect 6841 11886 6846 11914
rect 6874 11886 6879 11914
rect 6846 11746 6874 11886
rect 9193 11830 9198 11858
rect 9226 11830 9282 11858
rect 9921 11830 9926 11858
rect 9954 11830 10122 11858
rect 6846 11718 7686 11746
rect 7714 11718 7719 11746
rect 9254 11690 9282 11830
rect 9913 11746 9918 11774
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 10050 11746 10055 11774
rect 10094 11746 10122 11830
rect 20600 11802 21000 11816
rect 20001 11774 20006 11802
rect 20034 11774 21000 11802
rect 20600 11760 21000 11774
rect 10094 11718 10934 11746
rect 10962 11718 12278 11746
rect 12306 11718 12311 11746
rect 8297 11662 8302 11690
rect 8330 11662 8750 11690
rect 8778 11662 8783 11690
rect 9254 11662 9646 11690
rect 9674 11662 12222 11690
rect 12250 11662 12255 11690
rect 14625 11606 14630 11634
rect 14658 11606 15974 11634
rect 15946 11578 15974 11606
rect 8129 11550 8134 11578
rect 8162 11550 8358 11578
rect 8386 11550 9142 11578
rect 9170 11550 9175 11578
rect 15946 11550 18830 11578
rect 18858 11550 18863 11578
rect 7065 11494 7070 11522
rect 7098 11494 7966 11522
rect 7994 11494 7999 11522
rect 20600 11466 21000 11480
rect 8409 11438 8414 11466
rect 8442 11438 9030 11466
rect 9058 11438 9063 11466
rect 20001 11438 20006 11466
rect 20034 11438 21000 11466
rect 20600 11424 21000 11438
rect 12217 11382 12222 11410
rect 12250 11382 12782 11410
rect 12810 11382 12815 11410
rect 2233 11354 2238 11382
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2370 11354 2375 11382
rect 17593 11354 17598 11382
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17730 11354 17735 11382
rect 9249 11270 9254 11298
rect 9282 11270 9534 11298
rect 9562 11270 9567 11298
rect 8801 11214 8806 11242
rect 8834 11214 10346 11242
rect 10318 11186 10346 11214
rect 7681 11158 7686 11186
rect 7714 11158 8134 11186
rect 8162 11158 8167 11186
rect 9025 11158 9030 11186
rect 9058 11158 9366 11186
rect 9394 11158 9399 11186
rect 10313 11158 10318 11186
rect 10346 11158 11102 11186
rect 11130 11158 11135 11186
rect 15946 11158 18830 11186
rect 18858 11158 18863 11186
rect 9193 11102 9198 11130
rect 9226 11102 10094 11130
rect 10122 11102 10654 11130
rect 10682 11102 10687 11130
rect 15946 11074 15974 11158
rect 20600 11130 21000 11144
rect 20001 11102 20006 11130
rect 20034 11102 21000 11130
rect 20600 11088 21000 11102
rect 7905 11046 7910 11074
rect 7938 11046 8246 11074
rect 8274 11046 8694 11074
rect 8722 11046 8727 11074
rect 9473 11046 9478 11074
rect 9506 11046 9702 11074
rect 9730 11046 10710 11074
rect 10738 11046 10743 11074
rect 10873 11046 10878 11074
rect 10906 11046 11494 11074
rect 11522 11046 15974 11074
rect 8017 10990 8022 11018
rect 8050 10990 8470 11018
rect 8498 10990 8503 11018
rect 8857 10990 8862 11018
rect 8890 10990 9534 11018
rect 9562 10990 9567 11018
rect 9913 10962 9918 10990
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 10050 10962 10055 10990
rect 6393 10878 6398 10906
rect 6426 10878 6790 10906
rect 6818 10878 6823 10906
rect 9641 10878 9646 10906
rect 9674 10878 9870 10906
rect 9898 10878 10934 10906
rect 10962 10878 11382 10906
rect 11410 10878 11415 10906
rect 4186 10822 4998 10850
rect 5026 10822 6510 10850
rect 6538 10822 6543 10850
rect 10313 10822 10318 10850
rect 10346 10822 10710 10850
rect 10738 10822 10743 10850
rect 10817 10822 10822 10850
rect 10850 10822 11046 10850
rect 11074 10822 11550 10850
rect 11578 10822 13566 10850
rect 13594 10822 13599 10850
rect 4186 10794 4214 10822
rect 20600 10794 21000 10808
rect 2137 10766 2142 10794
rect 2170 10766 4214 10794
rect 6561 10766 6566 10794
rect 6594 10766 6958 10794
rect 6986 10766 7126 10794
rect 7154 10766 7159 10794
rect 8297 10766 8302 10794
rect 8330 10766 8862 10794
rect 8890 10766 8895 10794
rect 9137 10766 9142 10794
rect 9170 10766 9478 10794
rect 9506 10766 9511 10794
rect 9585 10766 9590 10794
rect 9618 10766 9870 10794
rect 9898 10766 9903 10794
rect 10201 10766 10206 10794
rect 10234 10766 11270 10794
rect 11298 10766 11303 10794
rect 15946 10766 18830 10794
rect 18858 10766 18863 10794
rect 20001 10766 20006 10794
rect 20034 10766 21000 10794
rect 10206 10738 10234 10766
rect 15946 10738 15974 10766
rect 20600 10752 21000 10766
rect 8465 10710 8470 10738
rect 8498 10710 10234 10738
rect 13617 10710 13622 10738
rect 13650 10710 14238 10738
rect 14266 10710 15974 10738
rect 6057 10654 6062 10682
rect 6090 10654 6790 10682
rect 6818 10654 6823 10682
rect 9137 10654 9142 10682
rect 9170 10654 9702 10682
rect 9730 10654 10038 10682
rect 10066 10654 10071 10682
rect 2233 10570 2238 10598
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2370 10570 2375 10598
rect 17593 10570 17598 10598
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17730 10570 17735 10598
rect 9534 10542 11942 10570
rect 11970 10542 11975 10570
rect 9534 10514 9562 10542
rect 6841 10486 6846 10514
rect 6874 10486 8806 10514
rect 8834 10486 8839 10514
rect 9529 10486 9534 10514
rect 9562 10486 9567 10514
rect 9641 10486 9646 10514
rect 9674 10486 9814 10514
rect 9842 10486 9847 10514
rect 0 10458 400 10472
rect 0 10430 966 10458
rect 994 10430 999 10458
rect 9025 10430 9030 10458
rect 9058 10430 9366 10458
rect 9394 10430 9399 10458
rect 12217 10430 12222 10458
rect 12250 10430 13174 10458
rect 13202 10430 13207 10458
rect 0 10416 400 10430
rect 2137 10374 2142 10402
rect 2170 10374 4214 10402
rect 6449 10374 6454 10402
rect 6482 10374 6734 10402
rect 6762 10374 7070 10402
rect 7098 10374 7103 10402
rect 10425 10374 10430 10402
rect 10458 10374 10934 10402
rect 10962 10374 11886 10402
rect 11914 10374 12166 10402
rect 12194 10374 12199 10402
rect 13113 10374 13118 10402
rect 13146 10374 13454 10402
rect 13482 10374 13487 10402
rect 4186 10234 4214 10374
rect 6958 10290 6986 10374
rect 8913 10318 8918 10346
rect 8946 10318 9310 10346
rect 9338 10318 10710 10346
rect 10738 10318 10743 10346
rect 11657 10318 11662 10346
rect 11690 10318 13734 10346
rect 13762 10318 13767 10346
rect 6953 10262 6958 10290
rect 6986 10262 6991 10290
rect 7065 10262 7070 10290
rect 7098 10262 7462 10290
rect 7490 10262 7495 10290
rect 9025 10262 9030 10290
rect 9058 10262 9114 10290
rect 9417 10262 9422 10290
rect 9450 10262 9926 10290
rect 9954 10262 9959 10290
rect 10369 10262 10374 10290
rect 10402 10262 10542 10290
rect 10570 10262 11494 10290
rect 11522 10262 11527 10290
rect 9086 10234 9114 10262
rect 4186 10206 5502 10234
rect 5530 10206 7014 10234
rect 7042 10206 7047 10234
rect 9086 10206 9814 10234
rect 9842 10206 9847 10234
rect 10705 10206 10710 10234
rect 10738 10206 11270 10234
rect 11298 10206 11303 10234
rect 9913 10178 9918 10206
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 10050 10178 10055 10206
rect 7121 10150 7126 10178
rect 7154 10150 7798 10178
rect 7826 10150 7831 10178
rect 9254 10150 9590 10178
rect 9618 10150 9623 10178
rect 11153 10150 11158 10178
rect 11186 10150 12838 10178
rect 12866 10150 13342 10178
rect 13370 10150 13375 10178
rect 0 10122 400 10136
rect 9254 10122 9282 10150
rect 0 10094 1022 10122
rect 1050 10094 1055 10122
rect 6561 10094 6566 10122
rect 6594 10094 7406 10122
rect 7434 10094 7439 10122
rect 8913 10094 8918 10122
rect 8946 10094 9030 10122
rect 9058 10094 9282 10122
rect 9361 10094 9366 10122
rect 9394 10094 9702 10122
rect 9730 10094 9735 10122
rect 10033 10094 10038 10122
rect 10066 10094 10990 10122
rect 11018 10094 11023 10122
rect 11321 10094 11326 10122
rect 11354 10094 11718 10122
rect 11746 10094 11751 10122
rect 0 10080 400 10094
rect 8409 10038 8414 10066
rect 8442 10038 9086 10066
rect 9114 10038 9119 10066
rect 7546 9982 8806 10010
rect 8834 9982 9310 10010
rect 9338 9982 9343 10010
rect 7546 9954 7574 9982
rect 2081 9926 2086 9954
rect 2114 9926 7574 9954
rect 9809 9926 9814 9954
rect 9842 9926 10318 9954
rect 10346 9926 10351 9954
rect 10369 9814 10374 9842
rect 10402 9814 11606 9842
rect 11634 9814 12054 9842
rect 12082 9814 12087 9842
rect 2233 9786 2238 9814
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2370 9786 2375 9814
rect 17593 9786 17598 9814
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17730 9786 17735 9814
rect 20600 9786 21000 9800
rect 20001 9758 20006 9786
rect 20034 9758 21000 9786
rect 20600 9744 21000 9758
rect 8801 9646 8806 9674
rect 8834 9646 11102 9674
rect 11130 9646 11550 9674
rect 11578 9646 11583 9674
rect 13729 9646 13734 9674
rect 13762 9646 18830 9674
rect 18858 9646 18863 9674
rect 7233 9590 7238 9618
rect 7266 9590 7574 9618
rect 7546 9338 7574 9590
rect 7966 9590 10346 9618
rect 7966 9506 7994 9590
rect 10318 9562 10346 9590
rect 8078 9534 9366 9562
rect 9394 9534 9399 9562
rect 9585 9534 9590 9562
rect 9618 9534 9926 9562
rect 9954 9534 9959 9562
rect 10313 9534 10318 9562
rect 10346 9534 11046 9562
rect 11074 9534 11079 9562
rect 12105 9534 12110 9562
rect 12138 9534 12670 9562
rect 12698 9534 12703 9562
rect 8078 9506 8106 9534
rect 7961 9478 7966 9506
rect 7994 9478 7999 9506
rect 8073 9478 8078 9506
rect 8106 9478 8111 9506
rect 8969 9478 8974 9506
rect 9002 9478 9758 9506
rect 9786 9478 11774 9506
rect 11802 9478 11807 9506
rect 9913 9394 9918 9422
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 10050 9394 10055 9422
rect 7546 9310 8218 9338
rect 9641 9310 9646 9338
rect 9674 9310 9870 9338
rect 9898 9310 10206 9338
rect 10234 9310 10598 9338
rect 10626 9310 10631 9338
rect 8190 9282 8218 9310
rect 6617 9254 6622 9282
rect 6650 9254 8078 9282
rect 8106 9254 8111 9282
rect 8185 9254 8190 9282
rect 8218 9254 10374 9282
rect 10402 9254 10407 9282
rect 11377 9254 11382 9282
rect 11410 9254 11942 9282
rect 11970 9254 11975 9282
rect 8241 9198 8246 9226
rect 8274 9198 8526 9226
rect 8554 9198 8694 9226
rect 8722 9198 8727 9226
rect 9641 9198 9646 9226
rect 9674 9198 10150 9226
rect 10178 9198 10183 9226
rect 10257 9198 10262 9226
rect 10290 9198 11158 9226
rect 11186 9198 11191 9226
rect 5553 9142 5558 9170
rect 5586 9142 7462 9170
rect 7490 9142 7495 9170
rect 7625 9142 7630 9170
rect 7658 9142 8134 9170
rect 8162 9142 9086 9170
rect 9114 9142 9119 9170
rect 9417 9142 9422 9170
rect 9450 9142 10542 9170
rect 10570 9142 10575 9170
rect 8857 9086 8862 9114
rect 8890 9086 9982 9114
rect 10010 9086 10015 9114
rect 9921 9030 9926 9058
rect 9954 9030 12894 9058
rect 12922 9030 12927 9058
rect 2233 9002 2238 9030
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2370 9002 2375 9030
rect 17593 9002 17598 9030
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17730 9002 17735 9030
rect 9529 8974 9534 9002
rect 9562 8974 10654 9002
rect 10682 8974 11326 9002
rect 11354 8974 11359 9002
rect 9193 8918 9198 8946
rect 9226 8918 9422 8946
rect 9450 8918 9870 8946
rect 9898 8918 10990 8946
rect 11018 8918 11023 8946
rect 6729 8862 6734 8890
rect 6762 8862 7574 8890
rect 7602 8862 8526 8890
rect 8554 8862 8559 8890
rect 9529 8862 9534 8890
rect 9562 8862 10122 8890
rect 10705 8862 10710 8890
rect 10738 8862 11886 8890
rect 11914 8862 11919 8890
rect 10094 8834 10122 8862
rect 8689 8806 8694 8834
rect 8722 8806 9254 8834
rect 9282 8806 9590 8834
rect 9618 8806 9623 8834
rect 10094 8806 10878 8834
rect 10906 8806 10911 8834
rect 20600 8778 21000 8792
rect 12049 8750 12054 8778
rect 12082 8750 12614 8778
rect 12642 8750 12647 8778
rect 20001 8750 20006 8778
rect 20034 8750 21000 8778
rect 20600 8736 21000 8750
rect 9025 8694 9030 8722
rect 9058 8694 9646 8722
rect 9674 8694 9679 8722
rect 10649 8694 10654 8722
rect 10682 8694 10878 8722
rect 10906 8694 10911 8722
rect 11601 8694 11606 8722
rect 11634 8694 12222 8722
rect 12250 8694 12255 8722
rect 14009 8694 14014 8722
rect 14042 8694 18942 8722
rect 18970 8694 18975 8722
rect 12777 8638 12782 8666
rect 12810 8638 13902 8666
rect 13930 8638 18830 8666
rect 18858 8638 18863 8666
rect 9913 8610 9918 8638
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 10050 8610 10055 8638
rect 11545 8582 11550 8610
rect 11578 8582 12222 8610
rect 12250 8582 12255 8610
rect 20600 8442 21000 8456
rect 20001 8414 20006 8442
rect 20034 8414 21000 8442
rect 20600 8400 21000 8414
rect 11825 8358 11830 8386
rect 11858 8358 12670 8386
rect 12698 8358 12703 8386
rect 10425 8302 10430 8330
rect 10458 8302 12614 8330
rect 12642 8302 12647 8330
rect 2233 8218 2238 8246
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2370 8218 2375 8246
rect 17593 8218 17598 8246
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17730 8218 17735 8246
rect 2137 8022 2142 8050
rect 2170 8022 5222 8050
rect 5250 8022 5255 8050
rect 9921 8022 9926 8050
rect 9954 8022 10710 8050
rect 10738 8022 10743 8050
rect 9305 7966 9310 7994
rect 9338 7966 9758 7994
rect 9786 7966 9791 7994
rect 5217 7910 5222 7938
rect 5250 7910 6790 7938
rect 6818 7910 6823 7938
rect 9913 7826 9918 7854
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 10050 7826 10055 7854
rect 0 7770 400 7784
rect 0 7742 966 7770
rect 994 7742 999 7770
rect 10425 7742 10430 7770
rect 10458 7742 10766 7770
rect 10794 7742 10799 7770
rect 0 7728 400 7742
rect 6897 7686 6902 7714
rect 6930 7686 7574 7714
rect 12329 7686 12334 7714
rect 12362 7686 12614 7714
rect 12642 7686 13286 7714
rect 13314 7686 13319 7714
rect 6281 7630 6286 7658
rect 6314 7630 7014 7658
rect 7042 7630 7047 7658
rect 7546 7602 7574 7686
rect 8297 7630 8302 7658
rect 8330 7630 9254 7658
rect 9282 7630 9814 7658
rect 9842 7630 9847 7658
rect 7546 7574 7630 7602
rect 7658 7574 10318 7602
rect 10346 7574 10351 7602
rect 2233 7434 2238 7462
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2370 7434 2375 7462
rect 17593 7434 17598 7462
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17730 7434 17735 7462
rect 9809 7294 9814 7322
rect 9842 7294 10346 7322
rect 6897 7238 6902 7266
rect 6930 7238 7182 7266
rect 7210 7238 8078 7266
rect 8106 7238 8302 7266
rect 8330 7238 8750 7266
rect 8778 7238 9702 7266
rect 9730 7238 10206 7266
rect 10234 7238 10239 7266
rect 10318 7210 10346 7294
rect 8409 7182 8414 7210
rect 8442 7182 9086 7210
rect 9114 7182 9119 7210
rect 10257 7182 10262 7210
rect 10290 7182 11102 7210
rect 11130 7182 11135 7210
rect 9913 7042 9918 7070
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 10050 7042 10055 7070
rect 9137 6902 9142 6930
rect 9170 6902 9534 6930
rect 9562 6902 9567 6930
rect 10201 6846 10206 6874
rect 10234 6846 11438 6874
rect 11466 6846 11471 6874
rect 11153 6734 11158 6762
rect 11186 6734 11606 6762
rect 11634 6734 12278 6762
rect 12306 6734 12311 6762
rect 2233 6650 2238 6678
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2370 6650 2375 6678
rect 17593 6650 17598 6678
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17730 6650 17735 6678
rect 9913 6258 9918 6286
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 10050 6258 10055 6286
rect 9753 5950 9758 5978
rect 9786 5950 10318 5978
rect 10346 5950 10710 5978
rect 10738 5950 10743 5978
rect 2233 5866 2238 5894
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2370 5866 2375 5894
rect 17593 5866 17598 5894
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17730 5866 17735 5894
rect 9913 5474 9918 5502
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 10050 5474 10055 5502
rect 2233 5082 2238 5110
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2370 5082 2375 5110
rect 17593 5082 17598 5110
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17730 5082 17735 5110
rect 9913 4690 9918 4718
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 10050 4690 10055 4718
rect 2233 4298 2238 4326
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2370 4298 2375 4326
rect 17593 4298 17598 4326
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17730 4298 17735 4326
rect 9913 3906 9918 3934
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 10050 3906 10055 3934
rect 2233 3514 2238 3542
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2370 3514 2375 3542
rect 17593 3514 17598 3542
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17730 3514 17735 3542
rect 9913 3122 9918 3150
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 10050 3122 10055 3150
rect 2233 2730 2238 2758
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2370 2730 2375 2758
rect 17593 2730 17598 2758
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17730 2730 17735 2758
rect 9913 2338 9918 2366
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 10050 2338 10055 2366
rect 9417 2030 9422 2058
rect 9450 2030 10038 2058
rect 10066 2030 10071 2058
rect 12441 2030 12446 2058
rect 12474 2030 13118 2058
rect 13146 2030 13151 2058
rect 2233 1946 2238 1974
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2370 1946 2375 1974
rect 17593 1946 17598 1974
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17730 1946 17735 1974
rect 11433 1806 11438 1834
rect 11466 1806 12782 1834
rect 12810 1806 12815 1834
rect 8409 1694 8414 1722
rect 8442 1694 9030 1722
rect 9058 1694 9063 1722
rect 9913 1554 9918 1582
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 10050 1554 10055 1582
<< via3 >>
rect 2238 19194 2266 19222
rect 2290 19194 2318 19222
rect 2342 19194 2370 19222
rect 17598 19194 17626 19222
rect 17650 19194 17678 19222
rect 17702 19194 17730 19222
rect 9918 18802 9946 18830
rect 9970 18802 9998 18830
rect 10022 18802 10050 18830
rect 2238 18410 2266 18438
rect 2290 18410 2318 18438
rect 2342 18410 2370 18438
rect 17598 18410 17626 18438
rect 17650 18410 17678 18438
rect 17702 18410 17730 18438
rect 9918 18018 9946 18046
rect 9970 18018 9998 18046
rect 10022 18018 10050 18046
rect 2238 17626 2266 17654
rect 2290 17626 2318 17654
rect 2342 17626 2370 17654
rect 17598 17626 17626 17654
rect 17650 17626 17678 17654
rect 17702 17626 17730 17654
rect 9918 17234 9946 17262
rect 9970 17234 9998 17262
rect 10022 17234 10050 17262
rect 2238 16842 2266 16870
rect 2290 16842 2318 16870
rect 2342 16842 2370 16870
rect 17598 16842 17626 16870
rect 17650 16842 17678 16870
rect 17702 16842 17730 16870
rect 9918 16450 9946 16478
rect 9970 16450 9998 16478
rect 10022 16450 10050 16478
rect 2238 16058 2266 16086
rect 2290 16058 2318 16086
rect 2342 16058 2370 16086
rect 17598 16058 17626 16086
rect 17650 16058 17678 16086
rect 17702 16058 17730 16086
rect 9918 15666 9946 15694
rect 9970 15666 9998 15694
rect 10022 15666 10050 15694
rect 2238 15274 2266 15302
rect 2290 15274 2318 15302
rect 2342 15274 2370 15302
rect 17598 15274 17626 15302
rect 17650 15274 17678 15302
rect 17702 15274 17730 15302
rect 9918 14882 9946 14910
rect 9970 14882 9998 14910
rect 10022 14882 10050 14910
rect 2238 14490 2266 14518
rect 2290 14490 2318 14518
rect 2342 14490 2370 14518
rect 17598 14490 17626 14518
rect 17650 14490 17678 14518
rect 17702 14490 17730 14518
rect 9918 14098 9946 14126
rect 9970 14098 9998 14126
rect 10022 14098 10050 14126
rect 2238 13706 2266 13734
rect 2290 13706 2318 13734
rect 2342 13706 2370 13734
rect 17598 13706 17626 13734
rect 17650 13706 17678 13734
rect 17702 13706 17730 13734
rect 9918 13314 9946 13342
rect 9970 13314 9998 13342
rect 10022 13314 10050 13342
rect 2238 12922 2266 12950
rect 2290 12922 2318 12950
rect 2342 12922 2370 12950
rect 17598 12922 17626 12950
rect 17650 12922 17678 12950
rect 17702 12922 17730 12950
rect 9918 12530 9946 12558
rect 9970 12530 9998 12558
rect 10022 12530 10050 12558
rect 2238 12138 2266 12166
rect 2290 12138 2318 12166
rect 2342 12138 2370 12166
rect 17598 12138 17626 12166
rect 17650 12138 17678 12166
rect 17702 12138 17730 12166
rect 9918 11746 9946 11774
rect 9970 11746 9998 11774
rect 10022 11746 10050 11774
rect 2238 11354 2266 11382
rect 2290 11354 2318 11382
rect 2342 11354 2370 11382
rect 17598 11354 17626 11382
rect 17650 11354 17678 11382
rect 17702 11354 17730 11382
rect 9918 10962 9946 10990
rect 9970 10962 9998 10990
rect 10022 10962 10050 10990
rect 2238 10570 2266 10598
rect 2290 10570 2318 10598
rect 2342 10570 2370 10598
rect 17598 10570 17626 10598
rect 17650 10570 17678 10598
rect 17702 10570 17730 10598
rect 9918 10178 9946 10206
rect 9970 10178 9998 10206
rect 10022 10178 10050 10206
rect 2238 9786 2266 9814
rect 2290 9786 2318 9814
rect 2342 9786 2370 9814
rect 17598 9786 17626 9814
rect 17650 9786 17678 9814
rect 17702 9786 17730 9814
rect 9918 9394 9946 9422
rect 9970 9394 9998 9422
rect 10022 9394 10050 9422
rect 2238 9002 2266 9030
rect 2290 9002 2318 9030
rect 2342 9002 2370 9030
rect 17598 9002 17626 9030
rect 17650 9002 17678 9030
rect 17702 9002 17730 9030
rect 9918 8610 9946 8638
rect 9970 8610 9998 8638
rect 10022 8610 10050 8638
rect 2238 8218 2266 8246
rect 2290 8218 2318 8246
rect 2342 8218 2370 8246
rect 17598 8218 17626 8246
rect 17650 8218 17678 8246
rect 17702 8218 17730 8246
rect 9918 7826 9946 7854
rect 9970 7826 9998 7854
rect 10022 7826 10050 7854
rect 2238 7434 2266 7462
rect 2290 7434 2318 7462
rect 2342 7434 2370 7462
rect 17598 7434 17626 7462
rect 17650 7434 17678 7462
rect 17702 7434 17730 7462
rect 9918 7042 9946 7070
rect 9970 7042 9998 7070
rect 10022 7042 10050 7070
rect 2238 6650 2266 6678
rect 2290 6650 2318 6678
rect 2342 6650 2370 6678
rect 17598 6650 17626 6678
rect 17650 6650 17678 6678
rect 17702 6650 17730 6678
rect 9918 6258 9946 6286
rect 9970 6258 9998 6286
rect 10022 6258 10050 6286
rect 2238 5866 2266 5894
rect 2290 5866 2318 5894
rect 2342 5866 2370 5894
rect 17598 5866 17626 5894
rect 17650 5866 17678 5894
rect 17702 5866 17730 5894
rect 9918 5474 9946 5502
rect 9970 5474 9998 5502
rect 10022 5474 10050 5502
rect 2238 5082 2266 5110
rect 2290 5082 2318 5110
rect 2342 5082 2370 5110
rect 17598 5082 17626 5110
rect 17650 5082 17678 5110
rect 17702 5082 17730 5110
rect 9918 4690 9946 4718
rect 9970 4690 9998 4718
rect 10022 4690 10050 4718
rect 2238 4298 2266 4326
rect 2290 4298 2318 4326
rect 2342 4298 2370 4326
rect 17598 4298 17626 4326
rect 17650 4298 17678 4326
rect 17702 4298 17730 4326
rect 9918 3906 9946 3934
rect 9970 3906 9998 3934
rect 10022 3906 10050 3934
rect 2238 3514 2266 3542
rect 2290 3514 2318 3542
rect 2342 3514 2370 3542
rect 17598 3514 17626 3542
rect 17650 3514 17678 3542
rect 17702 3514 17730 3542
rect 9918 3122 9946 3150
rect 9970 3122 9998 3150
rect 10022 3122 10050 3150
rect 2238 2730 2266 2758
rect 2290 2730 2318 2758
rect 2342 2730 2370 2758
rect 17598 2730 17626 2758
rect 17650 2730 17678 2758
rect 17702 2730 17730 2758
rect 9918 2338 9946 2366
rect 9970 2338 9998 2366
rect 10022 2338 10050 2366
rect 2238 1946 2266 1974
rect 2290 1946 2318 1974
rect 2342 1946 2370 1974
rect 17598 1946 17626 1974
rect 17650 1946 17678 1974
rect 17702 1946 17730 1974
rect 9918 1554 9946 1582
rect 9970 1554 9998 1582
rect 10022 1554 10050 1582
<< metal4 >>
rect 2224 19222 2384 19238
rect 2224 19194 2238 19222
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2370 19194 2384 19222
rect 2224 18438 2384 19194
rect 2224 18410 2238 18438
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2370 18410 2384 18438
rect 2224 17654 2384 18410
rect 2224 17626 2238 17654
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2370 17626 2384 17654
rect 2224 16870 2384 17626
rect 2224 16842 2238 16870
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2370 16842 2384 16870
rect 2224 16086 2384 16842
rect 2224 16058 2238 16086
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2370 16058 2384 16086
rect 2224 15302 2384 16058
rect 2224 15274 2238 15302
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2370 15274 2384 15302
rect 2224 14518 2384 15274
rect 2224 14490 2238 14518
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2370 14490 2384 14518
rect 2224 13734 2384 14490
rect 2224 13706 2238 13734
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2370 13706 2384 13734
rect 2224 12950 2384 13706
rect 2224 12922 2238 12950
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2370 12922 2384 12950
rect 2224 12166 2384 12922
rect 2224 12138 2238 12166
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2370 12138 2384 12166
rect 2224 11382 2384 12138
rect 2224 11354 2238 11382
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2370 11354 2384 11382
rect 2224 10598 2384 11354
rect 2224 10570 2238 10598
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2370 10570 2384 10598
rect 2224 9814 2384 10570
rect 2224 9786 2238 9814
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2370 9786 2384 9814
rect 2224 9030 2384 9786
rect 2224 9002 2238 9030
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2370 9002 2384 9030
rect 2224 8246 2384 9002
rect 2224 8218 2238 8246
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2370 8218 2384 8246
rect 2224 7462 2384 8218
rect 2224 7434 2238 7462
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2370 7434 2384 7462
rect 2224 6678 2384 7434
rect 2224 6650 2238 6678
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2370 6650 2384 6678
rect 2224 5894 2384 6650
rect 2224 5866 2238 5894
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2370 5866 2384 5894
rect 2224 5110 2384 5866
rect 2224 5082 2238 5110
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2370 5082 2384 5110
rect 2224 4326 2384 5082
rect 2224 4298 2238 4326
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2370 4298 2384 4326
rect 2224 3542 2384 4298
rect 2224 3514 2238 3542
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2370 3514 2384 3542
rect 2224 2758 2384 3514
rect 2224 2730 2238 2758
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2370 2730 2384 2758
rect 2224 1974 2384 2730
rect 2224 1946 2238 1974
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2370 1946 2384 1974
rect 2224 1538 2384 1946
rect 9904 18830 10064 19238
rect 9904 18802 9918 18830
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 10050 18802 10064 18830
rect 9904 18046 10064 18802
rect 9904 18018 9918 18046
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 10050 18018 10064 18046
rect 9904 17262 10064 18018
rect 9904 17234 9918 17262
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 10050 17234 10064 17262
rect 9904 16478 10064 17234
rect 9904 16450 9918 16478
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 10050 16450 10064 16478
rect 9904 15694 10064 16450
rect 9904 15666 9918 15694
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 10050 15666 10064 15694
rect 9904 14910 10064 15666
rect 9904 14882 9918 14910
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 10050 14882 10064 14910
rect 9904 14126 10064 14882
rect 9904 14098 9918 14126
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 10050 14098 10064 14126
rect 9904 13342 10064 14098
rect 9904 13314 9918 13342
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 10050 13314 10064 13342
rect 9904 12558 10064 13314
rect 9904 12530 9918 12558
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 10050 12530 10064 12558
rect 9904 11774 10064 12530
rect 9904 11746 9918 11774
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 10050 11746 10064 11774
rect 9904 10990 10064 11746
rect 9904 10962 9918 10990
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 10050 10962 10064 10990
rect 9904 10206 10064 10962
rect 9904 10178 9918 10206
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 10050 10178 10064 10206
rect 9904 9422 10064 10178
rect 9904 9394 9918 9422
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 10050 9394 10064 9422
rect 9904 8638 10064 9394
rect 9904 8610 9918 8638
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 10050 8610 10064 8638
rect 9904 7854 10064 8610
rect 9904 7826 9918 7854
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 10050 7826 10064 7854
rect 9904 7070 10064 7826
rect 9904 7042 9918 7070
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 10050 7042 10064 7070
rect 9904 6286 10064 7042
rect 9904 6258 9918 6286
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 10050 6258 10064 6286
rect 9904 5502 10064 6258
rect 9904 5474 9918 5502
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 10050 5474 10064 5502
rect 9904 4718 10064 5474
rect 9904 4690 9918 4718
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 10050 4690 10064 4718
rect 9904 3934 10064 4690
rect 9904 3906 9918 3934
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 10050 3906 10064 3934
rect 9904 3150 10064 3906
rect 9904 3122 9918 3150
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 10050 3122 10064 3150
rect 9904 2366 10064 3122
rect 9904 2338 9918 2366
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 10050 2338 10064 2366
rect 9904 1582 10064 2338
rect 9904 1554 9918 1582
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 10050 1554 10064 1582
rect 9904 1538 10064 1554
rect 17584 19222 17744 19238
rect 17584 19194 17598 19222
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17730 19194 17744 19222
rect 17584 18438 17744 19194
rect 17584 18410 17598 18438
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17730 18410 17744 18438
rect 17584 17654 17744 18410
rect 17584 17626 17598 17654
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17730 17626 17744 17654
rect 17584 16870 17744 17626
rect 17584 16842 17598 16870
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17730 16842 17744 16870
rect 17584 16086 17744 16842
rect 17584 16058 17598 16086
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17730 16058 17744 16086
rect 17584 15302 17744 16058
rect 17584 15274 17598 15302
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17730 15274 17744 15302
rect 17584 14518 17744 15274
rect 17584 14490 17598 14518
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17730 14490 17744 14518
rect 17584 13734 17744 14490
rect 17584 13706 17598 13734
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17730 13706 17744 13734
rect 17584 12950 17744 13706
rect 17584 12922 17598 12950
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17730 12922 17744 12950
rect 17584 12166 17744 12922
rect 17584 12138 17598 12166
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17730 12138 17744 12166
rect 17584 11382 17744 12138
rect 17584 11354 17598 11382
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17730 11354 17744 11382
rect 17584 10598 17744 11354
rect 17584 10570 17598 10598
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17730 10570 17744 10598
rect 17584 9814 17744 10570
rect 17584 9786 17598 9814
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17730 9786 17744 9814
rect 17584 9030 17744 9786
rect 17584 9002 17598 9030
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17730 9002 17744 9030
rect 17584 8246 17744 9002
rect 17584 8218 17598 8246
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17730 8218 17744 8246
rect 17584 7462 17744 8218
rect 17584 7434 17598 7462
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17730 7434 17744 7462
rect 17584 6678 17744 7434
rect 17584 6650 17598 6678
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17730 6650 17744 6678
rect 17584 5894 17744 6650
rect 17584 5866 17598 5894
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17730 5866 17744 5894
rect 17584 5110 17744 5866
rect 17584 5082 17598 5110
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17730 5082 17744 5110
rect 17584 4326 17744 5082
rect 17584 4298 17598 4326
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17730 4298 17744 4326
rect 17584 3542 17744 4298
rect 17584 3514 17598 3542
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17730 3514 17744 3542
rect 17584 2758 17744 3514
rect 17584 2730 17598 2758
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17730 2730 17744 2758
rect 17584 1974 17744 2730
rect 17584 1946 17598 1974
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17730 1946 17744 1974
rect 17584 1538 17744 1946
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _097_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 7392 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _098_
timestamp 1698175906
transform 1 0 8792 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _099_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8456 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _100_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9072 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _101_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9688 0 1 7840
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _102_
timestamp 1698175906
transform 1 0 10584 0 1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _103_
timestamp 1698175906
transform 1 0 9072 0 -1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _104_
timestamp 1698175906
transform -1 0 10808 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _105_
timestamp 1698175906
transform 1 0 10192 0 -1 10976
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _106_
timestamp 1698175906
transform 1 0 8288 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _107_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 9296 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _108_
timestamp 1698175906
transform 1 0 9576 0 -1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _109_
timestamp 1698175906
transform 1 0 11032 0 1 7056
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _110_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10584 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _111_
timestamp 1698175906
transform 1 0 9464 0 1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _112_
timestamp 1698175906
transform -1 0 7504 0 -1 12544
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _113_
timestamp 1698175906
transform -1 0 7224 0 1 11760
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _114_
timestamp 1698175906
transform 1 0 9296 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _115_
timestamp 1698175906
transform -1 0 8960 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _116_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9968 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _117_
timestamp 1698175906
transform 1 0 9520 0 1 8624
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _118_
timestamp 1698175906
transform -1 0 9072 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _119_
timestamp 1698175906
transform -1 0 8400 0 -1 10976
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _120_
timestamp 1698175906
transform -1 0 6944 0 1 11760
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _121_
timestamp 1698175906
transform -1 0 10192 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _122_
timestamp 1698175906
transform -1 0 9744 0 1 9408
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _123_
timestamp 1698175906
transform -1 0 11480 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _124_
timestamp 1698175906
transform -1 0 9296 0 -1 7056
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _125_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8960 0 -1 7840
box -43 -43 659 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _126_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 8232 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _127_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 7056 0 -1 8624
box -43 -43 715 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _128_
timestamp 1698175906
transform 1 0 7728 0 -1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _129_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9072 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _130_
timestamp 1698175906
transform -1 0 10472 0 1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _131_
timestamp 1698175906
transform -1 0 9240 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _132_
timestamp 1698175906
transform -1 0 8512 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _133_
timestamp 1698175906
transform 1 0 8344 0 1 10976
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _134_
timestamp 1698175906
transform 1 0 8624 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _135_
timestamp 1698175906
transform -1 0 8120 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _136_
timestamp 1698175906
transform 1 0 10192 0 1 7056
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _137_
timestamp 1698175906
transform -1 0 11032 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _138_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 8344 0 -1 9408
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _139_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9744 0 1 9408
box -43 -43 771 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _140_
timestamp 1698175906
transform -1 0 10640 0 -1 13328
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _141_
timestamp 1698175906
transform -1 0 11256 0 1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _142_
timestamp 1698175906
transform -1 0 10920 0 1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _143_
timestamp 1698175906
transform -1 0 10304 0 1 14112
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _144_
timestamp 1698175906
transform -1 0 9408 0 -1 14112
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _145_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9072 0 1 9408
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _146_
timestamp 1698175906
transform -1 0 10136 0 1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _147_
timestamp 1698175906
transform -1 0 13104 0 -1 14112
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _148_
timestamp 1698175906
transform -1 0 12432 0 -1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _149_
timestamp 1698175906
transform 1 0 10584 0 -1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _150_
timestamp 1698175906
transform 1 0 9632 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _151_
timestamp 1698175906
transform 1 0 10696 0 -1 12544
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _152_
timestamp 1698175906
transform -1 0 11200 0 1 11760
box -43 -43 659 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _153_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 7336 0 1 10192
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _154_
timestamp 1698175906
transform -1 0 7560 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _155_
timestamp 1698175906
transform 1 0 11200 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _156_
timestamp 1698175906
transform 1 0 10976 0 1 9408
box -43 -43 771 435
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _157_
timestamp 1698175906
transform 1 0 12712 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _158_
timestamp 1698175906
transform -1 0 13608 0 1 11760
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _159_
timestamp 1698175906
transform 1 0 11984 0 1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _160_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 13608 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _161_
timestamp 1698175906
transform 1 0 13328 0 1 10192
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _162_
timestamp 1698175906
transform 1 0 8624 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _163_
timestamp 1698175906
transform -1 0 10360 0 -1 9408
box -43 -43 659 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _164_
timestamp 1698175906
transform 1 0 7728 0 1 9408
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _165_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9800 0 1 8624
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _166_
timestamp 1698175906
transform 1 0 12880 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _167_
timestamp 1698175906
transform -1 0 6664 0 -1 10976
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _168_
timestamp 1698175906
transform -1 0 9296 0 1 10192
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _169_
timestamp 1698175906
transform -1 0 6944 0 -1 10976
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _170_
timestamp 1698175906
transform 1 0 13104 0 1 12544
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _171_
timestamp 1698175906
transform -1 0 13104 0 1 12544
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _172_
timestamp 1698175906
transform -1 0 9744 0 -1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _173_
timestamp 1698175906
transform 1 0 9408 0 1 10192
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _174_
timestamp 1698175906
transform 1 0 11200 0 -1 10976
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _175_
timestamp 1698175906
transform 1 0 11704 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _176_
timestamp 1698175906
transform 1 0 11760 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _177_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 11200 0 -1 9408
box -43 -43 883 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _178_
timestamp 1698175906
transform 1 0 12152 0 1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _179_
timestamp 1698175906
transform 1 0 12488 0 1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _180_
timestamp 1698175906
transform 1 0 10584 0 1 8624
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _181_
timestamp 1698175906
transform 1 0 12544 0 -1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _182_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 11704 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _183_
timestamp 1698175906
transform 1 0 11424 0 1 10192
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _184_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10808 0 1 10192
box -43 -43 659 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _185_
timestamp 1698175906
transform 1 0 11872 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _186_
timestamp 1698175906
transform 1 0 8736 0 -1 10976
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _187_
timestamp 1698175906
transform -1 0 9744 0 -1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _188_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 9464 0 -1 13328
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _189_
timestamp 1698175906
transform -1 0 10584 0 -1 7840
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _190_
timestamp 1698175906
transform 1 0 6664 0 1 7840
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _191_
timestamp 1698175906
transform 1 0 6776 0 -1 7840
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _192_
timestamp 1698175906
transform -1 0 8400 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _193_
timestamp 1698175906
transform -1 0 7784 0 1 7056
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _194_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10080 0 -1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _195_
timestamp 1698175906
transform -1 0 7168 0 -1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _196_
timestamp 1698175906
transform 1 0 7952 0 1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _197_
timestamp 1698175906
transform -1 0 7112 0 -1 9408
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _198_
timestamp 1698175906
transform -1 0 8288 0 1 8624
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _199_
timestamp 1698175906
transform 1 0 7840 0 1 11760
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _200_
timestamp 1698175906
transform 1 0 6608 0 -1 11760
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _201_
timestamp 1698175906
transform -1 0 11312 0 -1 6272
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _202_
timestamp 1698175906
transform 1 0 10080 0 -1 14112
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _203_
timestamp 1698175906
transform 1 0 8736 0 1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _204_
timestamp 1698175906
transform 1 0 11928 0 1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _205_
timestamp 1698175906
transform 1 0 10584 0 1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _206_
timestamp 1698175906
transform -1 0 7056 0 -1 10192
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _207_
timestamp 1698175906
transform 1 0 12768 0 -1 11760
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _208_
timestamp 1698175906
transform 1 0 12712 0 -1 10976
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _209_
timestamp 1698175906
transform -1 0 6552 0 1 10192
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _210_
timestamp 1698175906
transform 1 0 12544 0 -1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _211_
timestamp 1698175906
transform -1 0 12432 0 1 10976
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _212_
timestamp 1698175906
transform 1 0 11760 0 1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _213_
timestamp 1698175906
transform 1 0 12152 0 1 8624
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _214_
timestamp 1698175906
transform 1 0 12208 0 1 9408
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _215_
timestamp 1698175906
transform 1 0 7112 0 1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _216_
timestamp 1698175906
transform -1 0 6776 0 -1 7840
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _217_
timestamp 1698175906
transform 1 0 6776 0 -1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _221_
timestamp 1698175906
transform 1 0 14392 0 -1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _222_
timestamp 1698175906
transform 1 0 13776 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _223_
timestamp 1698175906
transform 1 0 9744 0 -1 14112
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__194__CLK dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 11816 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__195__CLK
timestamp 1698175906
transform 1 0 7616 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__196__CLK
timestamp 1698175906
transform 1 0 9688 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__197__CLK
timestamp 1698175906
transform 1 0 7224 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__198__CLK
timestamp 1698175906
transform 1 0 8288 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__199__CLK
timestamp 1698175906
transform 1 0 9912 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__200__CLK
timestamp 1698175906
transform 1 0 8232 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__201__CLK
timestamp 1698175906
transform 1 0 11424 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__202__CLK
timestamp 1698175906
transform -1 0 11928 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__203__CLK
timestamp 1698175906
transform 1 0 10752 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__204__CLK
timestamp 1698175906
transform 1 0 11816 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__205__CLK
timestamp 1698175906
transform 1 0 12320 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__206__CLK
timestamp 1698175906
transform 1 0 7168 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__207__CLK
timestamp 1698175906
transform 1 0 12656 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__208__CLK
timestamp 1698175906
transform 1 0 12320 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__209__CLK
timestamp 1698175906
transform 1 0 7056 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__210__CLK
timestamp 1698175906
transform 1 0 12040 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__211__CLK
timestamp 1698175906
transform 1 0 12544 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__212__CLK
timestamp 1698175906
transform 1 0 11648 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__213__CLK
timestamp 1698175906
transform 1 0 11592 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__214__CLK
timestamp 1698175906
transform -1 0 12264 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__215__CLK
timestamp 1698175906
transform 1 0 8736 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__216__CLK
timestamp 1698175906
transform 1 0 7168 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__217__CLK
timestamp 1698175906
transform 1 0 8736 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1698175906
transform 1 0 8792 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9240 0 -1 10192
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1698175906
transform 1 0 9296 0 -1 8624
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1698175906
transform 1 0 9464 0 -1 11760
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 784 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698175906
transform 1 0 2688 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698175906
transform 1 0 4592 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698175906
transform 1 0 6496 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_138 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8400 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_165 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9912 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_169
timestamp 1698175906
transform 1 0 10136 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_172
timestamp 1698175906
transform 1 0 10304 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_176 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10528 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_232
timestamp 1698175906
transform 1 0 13664 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_236
timestamp 1698175906
transform 1 0 13888 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_240
timestamp 1698175906
transform 1 0 14112 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_274
timestamp 1698175906
transform 1 0 16016 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_308
timestamp 1698175906
transform 1 0 17920 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_342
timestamp 1698175906
transform 1 0 19824 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_346
timestamp 1698175906
transform 1 0 20048 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_348
timestamp 1698175906
transform 1 0 20160 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 784 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698175906
transform 1 0 4368 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698175906
transform 1 0 4704 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698175906
transform 1 0 8288 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_142 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8624 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_150
timestamp 1698175906
transform 1 0 9072 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_154
timestamp 1698175906
transform 1 0 9296 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_156
timestamp 1698175906
transform 1 0 9408 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_183 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10920 0 -1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_199
timestamp 1698175906
transform 1 0 11816 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_207
timestamp 1698175906
transform 1 0 12264 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_209
timestamp 1698175906
transform 1 0 12376 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_238
timestamp 1698175906
transform 1 0 14000 0 -1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_270
timestamp 1698175906
transform 1 0 15792 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_278
timestamp 1698175906
transform 1 0 16240 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_282
timestamp 1698175906
transform 1 0 16464 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_346
timestamp 1698175906
transform 1 0 20048 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_348
timestamp 1698175906
transform 1 0 20160 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698175906
transform 1 0 784 0 1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698175906
transform 1 0 2576 0 1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698175906
transform 1 0 2744 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698175906
transform 1 0 6328 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_107
timestamp 1698175906
transform 1 0 6664 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_171
timestamp 1698175906
transform 1 0 10248 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_177
timestamp 1698175906
transform 1 0 10584 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_241
timestamp 1698175906
transform 1 0 14168 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698175906
transform 1 0 14504 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698175906
transform 1 0 18088 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_317
timestamp 1698175906
transform 1 0 18424 0 1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698175906
transform 1 0 784 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698175906
transform 1 0 4368 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698175906
transform 1 0 4704 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698175906
transform 1 0 8288 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_142
timestamp 1698175906
transform 1 0 8624 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_206
timestamp 1698175906
transform 1 0 12208 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_212
timestamp 1698175906
transform 1 0 12544 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_276
timestamp 1698175906
transform 1 0 16128 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_282
timestamp 1698175906
transform 1 0 16464 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_346
timestamp 1698175906
transform 1 0 20048 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_348
timestamp 1698175906
transform 1 0 20160 0 -1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698175906
transform 1 0 784 0 1 3136
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698175906
transform 1 0 2576 0 1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698175906
transform 1 0 2744 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698175906
transform 1 0 6328 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_107
timestamp 1698175906
transform 1 0 6664 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698175906
transform 1 0 10248 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_177
timestamp 1698175906
transform 1 0 10584 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_241
timestamp 1698175906
transform 1 0 14168 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698175906
transform 1 0 14504 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698175906
transform 1 0 18088 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_317
timestamp 1698175906
transform 1 0 18424 0 1 3136
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698175906
transform 1 0 784 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698175906
transform 1 0 4368 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698175906
transform 1 0 4704 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698175906
transform 1 0 8288 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_142
timestamp 1698175906
transform 1 0 8624 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_206
timestamp 1698175906
transform 1 0 12208 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_212
timestamp 1698175906
transform 1 0 12544 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698175906
transform 1 0 16128 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_282
timestamp 1698175906
transform 1 0 16464 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_346
timestamp 1698175906
transform 1 0 20048 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_348
timestamp 1698175906
transform 1 0 20160 0 -1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698175906
transform 1 0 784 0 1 3920
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698175906
transform 1 0 2576 0 1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698175906
transform 1 0 2744 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698175906
transform 1 0 6328 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_107
timestamp 1698175906
transform 1 0 6664 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_171
timestamp 1698175906
transform 1 0 10248 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_177
timestamp 1698175906
transform 1 0 10584 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_241
timestamp 1698175906
transform 1 0 14168 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_247
timestamp 1698175906
transform 1 0 14504 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_311
timestamp 1698175906
transform 1 0 18088 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_317
timestamp 1698175906
transform 1 0 18424 0 1 3920
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698175906
transform 1 0 784 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698175906
transform 1 0 4368 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_72
timestamp 1698175906
transform 1 0 4704 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698175906
transform 1 0 8288 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_142
timestamp 1698175906
transform 1 0 8624 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_206
timestamp 1698175906
transform 1 0 12208 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_212
timestamp 1698175906
transform 1 0 12544 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_276
timestamp 1698175906
transform 1 0 16128 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_282
timestamp 1698175906
transform 1 0 16464 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_346
timestamp 1698175906
transform 1 0 20048 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_348
timestamp 1698175906
transform 1 0 20160 0 -1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698175906
transform 1 0 784 0 1 4704
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698175906
transform 1 0 2576 0 1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_37
timestamp 1698175906
transform 1 0 2744 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_101
timestamp 1698175906
transform 1 0 6328 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_107
timestamp 1698175906
transform 1 0 6664 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_171
timestamp 1698175906
transform 1 0 10248 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_177
timestamp 1698175906
transform 1 0 10584 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_241
timestamp 1698175906
transform 1 0 14168 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_247
timestamp 1698175906
transform 1 0 14504 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_311
timestamp 1698175906
transform 1 0 18088 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_317
timestamp 1698175906
transform 1 0 18424 0 1 4704
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698175906
transform 1 0 784 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698175906
transform 1 0 4368 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_72
timestamp 1698175906
transform 1 0 4704 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_136
timestamp 1698175906
transform 1 0 8288 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_142
timestamp 1698175906
transform 1 0 8624 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_206
timestamp 1698175906
transform 1 0 12208 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_212
timestamp 1698175906
transform 1 0 12544 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_276
timestamp 1698175906
transform 1 0 16128 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_282
timestamp 1698175906
transform 1 0 16464 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_346
timestamp 1698175906
transform 1 0 20048 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_348
timestamp 1698175906
transform 1 0 20160 0 -1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698175906
transform 1 0 784 0 1 5488
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698175906
transform 1 0 2576 0 1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_37
timestamp 1698175906
transform 1 0 2744 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698175906
transform 1 0 6328 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_107
timestamp 1698175906
transform 1 0 6664 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_171
timestamp 1698175906
transform 1 0 10248 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_177
timestamp 1698175906
transform 1 0 10584 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_241
timestamp 1698175906
transform 1 0 14168 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_247
timestamp 1698175906
transform 1 0 14504 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_311
timestamp 1698175906
transform 1 0 18088 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_317
timestamp 1698175906
transform 1 0 18424 0 1 5488
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2
timestamp 1698175906
transform 1 0 784 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698175906
transform 1 0 4368 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_72
timestamp 1698175906
transform 1 0 4704 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698175906
transform 1 0 8288 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_142
timestamp 1698175906
transform 1 0 8624 0 -1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_158
timestamp 1698175906
transform 1 0 9520 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_160
timestamp 1698175906
transform 1 0 9632 0 -1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_190
timestamp 1698175906
transform 1 0 11312 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_194
timestamp 1698175906
transform 1 0 11536 0 -1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_212
timestamp 1698175906
transform 1 0 12544 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_276
timestamp 1698175906
transform 1 0 16128 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_282
timestamp 1698175906
transform 1 0 16464 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_346
timestamp 1698175906
transform 1 0 20048 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_348
timestamp 1698175906
transform 1 0 20160 0 -1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698175906
transform 1 0 784 0 1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698175906
transform 1 0 2576 0 1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_37
timestamp 1698175906
transform 1 0 2744 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698175906
transform 1 0 6328 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_107
timestamp 1698175906
transform 1 0 6664 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_171
timestamp 1698175906
transform 1 0 10248 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_177
timestamp 1698175906
transform 1 0 10584 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_241
timestamp 1698175906
transform 1 0 14168 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_247
timestamp 1698175906
transform 1 0 14504 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_311
timestamp 1698175906
transform 1 0 18088 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_317
timestamp 1698175906
transform 1 0 18424 0 1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_2
timestamp 1698175906
transform 1 0 784 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_66
timestamp 1698175906
transform 1 0 4368 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_72
timestamp 1698175906
transform 1 0 4704 0 -1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_104
timestamp 1698175906
transform 1 0 6496 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_108
timestamp 1698175906
transform 1 0 6720 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_138
timestamp 1698175906
transform 1 0 8400 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_142
timestamp 1698175906
transform 1 0 8624 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_146
timestamp 1698175906
transform 1 0 8848 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_148
timestamp 1698175906
transform 1 0 8960 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_154
timestamp 1698175906
transform 1 0 9296 0 -1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_162
timestamp 1698175906
transform 1 0 9744 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_166
timestamp 1698175906
transform 1 0 9968 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_197
timestamp 1698175906
transform 1 0 11704 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_201
timestamp 1698175906
transform 1 0 11928 0 -1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_209
timestamp 1698175906
transform 1 0 12376 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_212
timestamp 1698175906
transform 1 0 12544 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_276
timestamp 1698175906
transform 1 0 16128 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_282
timestamp 1698175906
transform 1 0 16464 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_346
timestamp 1698175906
transform 1 0 20048 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_348
timestamp 1698175906
transform 1 0 20160 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698175906
transform 1 0 784 0 1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698175906
transform 1 0 2576 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_37
timestamp 1698175906
transform 1 0 2744 0 1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_101
timestamp 1698175906
transform 1 0 6328 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_107
timestamp 1698175906
transform 1 0 6664 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_115
timestamp 1698175906
transform 1 0 7112 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_119
timestamp 1698175906
transform 1 0 7336 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_121
timestamp 1698175906
transform 1 0 7448 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_127
timestamp 1698175906
transform 1 0 7784 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_129
timestamp 1698175906
transform 1 0 7896 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_159
timestamp 1698175906
transform 1 0 9576 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_163
timestamp 1698175906
transform 1 0 9800 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_167
timestamp 1698175906
transform 1 0 10024 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_169
timestamp 1698175906
transform 1 0 10136 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_190
timestamp 1698175906
transform 1 0 11312 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_194
timestamp 1698175906
transform 1 0 11536 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_227
timestamp 1698175906
transform 1 0 13384 0 1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_243
timestamp 1698175906
transform 1 0 14280 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_247
timestamp 1698175906
transform 1 0 14504 0 1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_311
timestamp 1698175906
transform 1 0 18088 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_317
timestamp 1698175906
transform 1 0 18424 0 1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_2
timestamp 1698175906
transform 1 0 784 0 -1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_66
timestamp 1698175906
transform 1 0 4368 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_72
timestamp 1698175906
transform 1 0 4704 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_114
timestamp 1698175906
transform 1 0 7056 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_118
timestamp 1698175906
transform 1 0 7280 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_126
timestamp 1698175906
transform 1 0 7728 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_138
timestamp 1698175906
transform 1 0 8400 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_142
timestamp 1698175906
transform 1 0 8624 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_146
timestamp 1698175906
transform 1 0 8848 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_165
timestamp 1698175906
transform 1 0 9912 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_169
timestamp 1698175906
transform 1 0 10136 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_171
timestamp 1698175906
transform 1 0 10248 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_185
timestamp 1698175906
transform 1 0 11032 0 -1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_201
timestamp 1698175906
transform 1 0 11928 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_209
timestamp 1698175906
transform 1 0 12376 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_212
timestamp 1698175906
transform 1 0 12544 0 -1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_276
timestamp 1698175906
transform 1 0 16128 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_282
timestamp 1698175906
transform 1 0 16464 0 -1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_346
timestamp 1698175906
transform 1 0 20048 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_348
timestamp 1698175906
transform 1 0 20160 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_28
timestamp 1698175906
transform 1 0 2240 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_32
timestamp 1698175906
transform 1 0 2464 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698175906
transform 1 0 2576 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_37
timestamp 1698175906
transform 1 0 2744 0 1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_101
timestamp 1698175906
transform 1 0 6328 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_112
timestamp 1698175906
transform 1 0 6944 0 1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_144
timestamp 1698175906
transform 1 0 8736 0 1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_160
timestamp 1698175906
transform 1 0 9632 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_166
timestamp 1698175906
transform 1 0 9968 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_174
timestamp 1698175906
transform 1 0 10416 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_183
timestamp 1698175906
transform 1 0 10920 0 1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_199
timestamp 1698175906
transform 1 0 11816 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_203
timestamp 1698175906
transform 1 0 12040 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_217
timestamp 1698175906
transform 1 0 12824 0 1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_233
timestamp 1698175906
transform 1 0 13720 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_241
timestamp 1698175906
transform 1 0 14168 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_247
timestamp 1698175906
transform 1 0 14504 0 1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_311
timestamp 1698175906
transform 1 0 18088 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_317
timestamp 1698175906
transform 1 0 18424 0 1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_2
timestamp 1698175906
transform 1 0 784 0 -1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_66
timestamp 1698175906
transform 1 0 4368 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_72
timestamp 1698175906
transform 1 0 4704 0 -1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_104
timestamp 1698175906
transform 1 0 6496 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_112
timestamp 1698175906
transform 1 0 6944 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_132
timestamp 1698175906
transform 1 0 8064 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_138
timestamp 1698175906
transform 1 0 8400 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_142
timestamp 1698175906
transform 1 0 8624 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_204
timestamp 1698175906
transform 1 0 12096 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_208
timestamp 1698175906
transform 1 0 12320 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_218
timestamp 1698175906
transform 1 0 12880 0 -1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_250
timestamp 1698175906
transform 1 0 14672 0 -1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_266
timestamp 1698175906
transform 1 0 15568 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_274
timestamp 1698175906
transform 1 0 16016 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_278
timestamp 1698175906
transform 1 0 16240 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_282
timestamp 1698175906
transform 1 0 16464 0 -1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_314
timestamp 1698175906
transform 1 0 18256 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_322
timestamp 1698175906
transform 1 0 18704 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_2
timestamp 1698175906
transform 1 0 784 0 1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698175906
transform 1 0 2576 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_37
timestamp 1698175906
transform 1 0 2744 0 1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_101
timestamp 1698175906
transform 1 0 6328 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_136
timestamp 1698175906
transform 1 0 8288 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_138
timestamp 1698175906
transform 1 0 8400 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_151
timestamp 1698175906
transform 1 0 9128 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_155
timestamp 1698175906
transform 1 0 9352 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_157
timestamp 1698175906
transform 1 0 9464 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_173
timestamp 1698175906
transform 1 0 10360 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_193
timestamp 1698175906
transform 1 0 11480 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_240
timestamp 1698175906
transform 1 0 14112 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_244
timestamp 1698175906
transform 1 0 14336 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_247
timestamp 1698175906
transform 1 0 14504 0 1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_311
timestamp 1698175906
transform 1 0 18088 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_317
timestamp 1698175906
transform 1 0 18424 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_321
timestamp 1698175906
transform 1 0 18648 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_2
timestamp 1698175906
transform 1 0 784 0 -1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_66
timestamp 1698175906
transform 1 0 4368 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_72
timestamp 1698175906
transform 1 0 4704 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_80
timestamp 1698175906
transform 1 0 5152 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_84
timestamp 1698175906
transform 1 0 5376 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_115
timestamp 1698175906
transform 1 0 7112 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_119
timestamp 1698175906
transform 1 0 7336 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_126
timestamp 1698175906
transform 1 0 7728 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_137
timestamp 1698175906
transform 1 0 8344 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_139
timestamp 1698175906
transform 1 0 8456 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_148
timestamp 1698175906
transform 1 0 8960 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_158
timestamp 1698175906
transform 1 0 9520 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_196
timestamp 1698175906
transform 1 0 11648 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_206
timestamp 1698175906
transform 1 0 12208 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_212
timestamp 1698175906
transform 1 0 12544 0 -1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_276
timestamp 1698175906
transform 1 0 16128 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_282
timestamp 1698175906
transform 1 0 16464 0 -1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_346
timestamp 1698175906
transform 1 0 20048 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_348
timestamp 1698175906
transform 1 0 20160 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_2
timestamp 1698175906
transform 1 0 784 0 1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698175906
transform 1 0 2576 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_37
timestamp 1698175906
transform 1 0 2744 0 1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_101
timestamp 1698175906
transform 1 0 6328 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_107
timestamp 1698175906
transform 1 0 6664 0 1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_123
timestamp 1698175906
transform 1 0 7560 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_125
timestamp 1698175906
transform 1 0 7672 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_135
timestamp 1698175906
transform 1 0 8232 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_143
timestamp 1698175906
transform 1 0 8680 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_177
timestamp 1698175906
transform 1 0 10584 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_181
timestamp 1698175906
transform 1 0 10808 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_183
timestamp 1698175906
transform 1 0 10920 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_203
timestamp 1698175906
transform 1 0 12040 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_205
timestamp 1698175906
transform 1 0 12152 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_235
timestamp 1698175906
transform 1 0 13832 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_243
timestamp 1698175906
transform 1 0 14280 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_247
timestamp 1698175906
transform 1 0 14504 0 1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_311
timestamp 1698175906
transform 1 0 18088 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_317
timestamp 1698175906
transform 1 0 18424 0 1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_2
timestamp 1698175906
transform 1 0 784 0 -1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_66
timestamp 1698175906
transform 1 0 4368 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_72
timestamp 1698175906
transform 1 0 4704 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_80
timestamp 1698175906
transform 1 0 5152 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_84
timestamp 1698175906
transform 1 0 5376 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_114
timestamp 1698175906
transform 1 0 7056 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_118
timestamp 1698175906
transform 1 0 7280 0 -1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_142
timestamp 1698175906
transform 1 0 8624 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_144
timestamp 1698175906
transform 1 0 8736 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_203
timestamp 1698175906
transform 1 0 12040 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_207
timestamp 1698175906
transform 1 0 12264 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_209
timestamp 1698175906
transform 1 0 12376 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_212
timestamp 1698175906
transform 1 0 12544 0 -1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_276
timestamp 1698175906
transform 1 0 16128 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_282
timestamp 1698175906
transform 1 0 16464 0 -1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_314
timestamp 1698175906
transform 1 0 18256 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_322
timestamp 1698175906
transform 1 0 18704 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_28
timestamp 1698175906
transform 1 0 2240 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_32
timestamp 1698175906
transform 1 0 2464 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698175906
transform 1 0 2576 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_37
timestamp 1698175906
transform 1 0 2744 0 1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_69
timestamp 1698175906
transform 1 0 4536 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_73
timestamp 1698175906
transform 1 0 4760 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_75
timestamp 1698175906
transform 1 0 4872 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_107
timestamp 1698175906
transform 1 0 6664 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_109
timestamp 1698175906
transform 1 0 6776 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_123
timestamp 1698175906
transform 1 0 7560 0 1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_139
timestamp 1698175906
transform 1 0 8456 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_143
timestamp 1698175906
transform 1 0 8680 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_154
timestamp 1698175906
transform 1 0 9296 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_177
timestamp 1698175906
transform 1 0 10584 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_208
timestamp 1698175906
transform 1 0 12320 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_216
timestamp 1698175906
transform 1 0 12768 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_233
timestamp 1698175906
transform 1 0 13720 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_241
timestamp 1698175906
transform 1 0 14168 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_247
timestamp 1698175906
transform 1 0 14504 0 1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_311
timestamp 1698175906
transform 1 0 18088 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_317
timestamp 1698175906
transform 1 0 18424 0 1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_28
timestamp 1698175906
transform 1 0 2240 0 -1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_60
timestamp 1698175906
transform 1 0 4032 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_68
timestamp 1698175906
transform 1 0 4480 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_72
timestamp 1698175906
transform 1 0 4704 0 -1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_88
timestamp 1698175906
transform 1 0 5600 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_96
timestamp 1698175906
transform 1 0 6048 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_100
timestamp 1698175906
transform 1 0 6272 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_112
timestamp 1698175906
transform 1 0 6944 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_116
timestamp 1698175906
transform 1 0 7168 0 -1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_132
timestamp 1698175906
transform 1 0 8064 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_138
timestamp 1698175906
transform 1 0 8400 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_142
timestamp 1698175906
transform 1 0 8624 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_153
timestamp 1698175906
transform 1 0 9240 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_155
timestamp 1698175906
transform 1 0 9352 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_175
timestamp 1698175906
transform 1 0 10472 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_183
timestamp 1698175906
transform 1 0 10920 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_187
timestamp 1698175906
transform 1 0 11144 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_206
timestamp 1698175906
transform 1 0 12208 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_212
timestamp 1698175906
transform 1 0 12544 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_214
timestamp 1698175906
transform 1 0 12656 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_244
timestamp 1698175906
transform 1 0 14336 0 -1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_276
timestamp 1698175906
transform 1 0 16128 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_282
timestamp 1698175906
transform 1 0 16464 0 -1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_314
timestamp 1698175906
transform 1 0 18256 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_322
timestamp 1698175906
transform 1 0 18704 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_2
timestamp 1698175906
transform 1 0 784 0 1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698175906
transform 1 0 2576 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_37
timestamp 1698175906
transform 1 0 2744 0 1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_101
timestamp 1698175906
transform 1 0 6328 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_107
timestamp 1698175906
transform 1 0 6664 0 1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_123
timestamp 1698175906
transform 1 0 7560 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_133
timestamp 1698175906
transform 1 0 8120 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_174
timestamp 1698175906
transform 1 0 10416 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_210
timestamp 1698175906
transform 1 0 12432 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_214
timestamp 1698175906
transform 1 0 12656 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_231
timestamp 1698175906
transform 1 0 13608 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_239
timestamp 1698175906
transform 1 0 14056 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_243
timestamp 1698175906
transform 1 0 14280 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_247
timestamp 1698175906
transform 1 0 14504 0 1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_311
timestamp 1698175906
transform 1 0 18088 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_317
timestamp 1698175906
transform 1 0 18424 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_321
timestamp 1698175906
transform 1 0 18648 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_2
timestamp 1698175906
transform 1 0 784 0 -1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_66
timestamp 1698175906
transform 1 0 4368 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_72
timestamp 1698175906
transform 1 0 4704 0 -1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_104
timestamp 1698175906
transform 1 0 6496 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_135
timestamp 1698175906
transform 1 0 8232 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_156
timestamp 1698175906
transform 1 0 9408 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_207
timestamp 1698175906
transform 1 0 12264 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_209
timestamp 1698175906
transform 1 0 12376 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_212
timestamp 1698175906
transform 1 0 12544 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_251
timestamp 1698175906
transform 1 0 14728 0 -1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_267
timestamp 1698175906
transform 1 0 15624 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_275
timestamp 1698175906
transform 1 0 16072 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_279
timestamp 1698175906
transform 1 0 16296 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_282
timestamp 1698175906
transform 1 0 16464 0 -1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_314
timestamp 1698175906
transform 1 0 18256 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_322
timestamp 1698175906
transform 1 0 18704 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_2
timestamp 1698175906
transform 1 0 784 0 1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698175906
transform 1 0 2576 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_37
timestamp 1698175906
transform 1 0 2744 0 1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_101
timestamp 1698175906
transform 1 0 6328 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_117
timestamp 1698175906
transform 1 0 7224 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_125
timestamp 1698175906
transform 1 0 7672 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_127
timestamp 1698175906
transform 1 0 7784 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_163
timestamp 1698175906
transform 1 0 9800 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_167
timestamp 1698175906
transform 1 0 10024 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_188
timestamp 1698175906
transform 1 0 11200 0 1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_220
timestamp 1698175906
transform 1 0 12992 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_224
timestamp 1698175906
transform 1 0 13216 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_231
timestamp 1698175906
transform 1 0 13608 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_239
timestamp 1698175906
transform 1 0 14056 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_243
timestamp 1698175906
transform 1 0 14280 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_247
timestamp 1698175906
transform 1 0 14504 0 1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_311
timestamp 1698175906
transform 1 0 18088 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_317
timestamp 1698175906
transform 1 0 18424 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_321
timestamp 1698175906
transform 1 0 18648 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_28
timestamp 1698175906
transform 1 0 2240 0 -1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_60
timestamp 1698175906
transform 1 0 4032 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_68
timestamp 1698175906
transform 1 0 4480 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_72
timestamp 1698175906
transform 1 0 4704 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_80
timestamp 1698175906
transform 1 0 5152 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_84
timestamp 1698175906
transform 1 0 5376 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_86
timestamp 1698175906
transform 1 0 5488 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_122
timestamp 1698175906
transform 1 0 7504 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_126
timestamp 1698175906
transform 1 0 7728 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_134
timestamp 1698175906
transform 1 0 8176 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_138
timestamp 1698175906
transform 1 0 8400 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_142
timestamp 1698175906
transform 1 0 8624 0 -1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_174
timestamp 1698175906
transform 1 0 10416 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_178
timestamp 1698175906
transform 1 0 10640 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_184
timestamp 1698175906
transform 1 0 10976 0 -1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_200
timestamp 1698175906
transform 1 0 11872 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_208
timestamp 1698175906
transform 1 0 12320 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_212
timestamp 1698175906
transform 1 0 12544 0 -1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_276
timestamp 1698175906
transform 1 0 16128 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_282
timestamp 1698175906
transform 1 0 16464 0 -1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_346
timestamp 1698175906
transform 1 0 20048 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_348
timestamp 1698175906
transform 1 0 20160 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_2
timestamp 1698175906
transform 1 0 784 0 1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698175906
transform 1 0 2576 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_37
timestamp 1698175906
transform 1 0 2744 0 1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_101
timestamp 1698175906
transform 1 0 6328 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_107
timestamp 1698175906
transform 1 0 6664 0 1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_171
timestamp 1698175906
transform 1 0 10248 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_206
timestamp 1698175906
transform 1 0 12208 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_210
timestamp 1698175906
transform 1 0 12432 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_214
timestamp 1698175906
transform 1 0 12656 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_216
timestamp 1698175906
transform 1 0 12768 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_227
timestamp 1698175906
transform 1 0 13384 0 1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_243
timestamp 1698175906
transform 1 0 14280 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_247
timestamp 1698175906
transform 1 0 14504 0 1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_311
timestamp 1698175906
transform 1 0 18088 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_317
timestamp 1698175906
transform 1 0 18424 0 1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_2
timestamp 1698175906
transform 1 0 784 0 -1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_66
timestamp 1698175906
transform 1 0 4368 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_72
timestamp 1698175906
transform 1 0 4704 0 -1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_136
timestamp 1698175906
transform 1 0 8288 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_142
timestamp 1698175906
transform 1 0 8624 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_146
timestamp 1698175906
transform 1 0 8848 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_162
timestamp 1698175906
transform 1 0 9744 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_170
timestamp 1698175906
transform 1 0 10192 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_178
timestamp 1698175906
transform 1 0 10640 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_182
timestamp 1698175906
transform 1 0 10864 0 -1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_198
timestamp 1698175906
transform 1 0 11760 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_202
timestamp 1698175906
transform 1 0 11984 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_241
timestamp 1698175906
transform 1 0 14168 0 -1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_273
timestamp 1698175906
transform 1 0 15960 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_277
timestamp 1698175906
transform 1 0 16184 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_279
timestamp 1698175906
transform 1 0 16296 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_282
timestamp 1698175906
transform 1 0 16464 0 -1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_346
timestamp 1698175906
transform 1 0 20048 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_348
timestamp 1698175906
transform 1 0 20160 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_2
timestamp 1698175906
transform 1 0 784 0 1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698175906
transform 1 0 2576 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_37
timestamp 1698175906
transform 1 0 2744 0 1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_101
timestamp 1698175906
transform 1 0 6328 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_107
timestamp 1698175906
transform 1 0 6664 0 1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_173
timestamp 1698175906
transform 1 0 10360 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_177
timestamp 1698175906
transform 1 0 10584 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_183
timestamp 1698175906
transform 1 0 10920 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_189
timestamp 1698175906
transform 1 0 11256 0 1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_197
timestamp 1698175906
transform 1 0 11704 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_230
timestamp 1698175906
transform 1 0 13552 0 1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_238
timestamp 1698175906
transform 1 0 14000 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_242
timestamp 1698175906
transform 1 0 14224 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_244
timestamp 1698175906
transform 1 0 14336 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_247
timestamp 1698175906
transform 1 0 14504 0 1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_311
timestamp 1698175906
transform 1 0 18088 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_317
timestamp 1698175906
transform 1 0 18424 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_321
timestamp 1698175906
transform 1 0 18648 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_2
timestamp 1698175906
transform 1 0 784 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_66
timestamp 1698175906
transform 1 0 4368 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_72
timestamp 1698175906
transform 1 0 4704 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_136
timestamp 1698175906
transform 1 0 8288 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_142
timestamp 1698175906
transform 1 0 8624 0 -1 14112
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_150
timestamp 1698175906
transform 1 0 9072 0 -1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_156
timestamp 1698175906
transform 1 0 9408 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_160
timestamp 1698175906
transform 1 0 9632 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_197
timestamp 1698175906
transform 1 0 11704 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_201
timestamp 1698175906
transform 1 0 11928 0 -1 14112
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_209
timestamp 1698175906
transform 1 0 12376 0 -1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_212
timestamp 1698175906
transform 1 0 12544 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_216
timestamp 1698175906
transform 1 0 12768 0 -1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_222
timestamp 1698175906
transform 1 0 13104 0 -1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_254
timestamp 1698175906
transform 1 0 14896 0 -1 14112
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_270
timestamp 1698175906
transform 1 0 15792 0 -1 14112
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_278
timestamp 1698175906
transform 1 0 16240 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_282
timestamp 1698175906
transform 1 0 16464 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_346
timestamp 1698175906
transform 1 0 20048 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_348
timestamp 1698175906
transform 1 0 20160 0 -1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_2
timestamp 1698175906
transform 1 0 784 0 1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698175906
transform 1 0 2576 0 1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_37
timestamp 1698175906
transform 1 0 2744 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_101
timestamp 1698175906
transform 1 0 6328 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_107
timestamp 1698175906
transform 1 0 6664 0 1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_139
timestamp 1698175906
transform 1 0 8456 0 1 14112
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_155
timestamp 1698175906
transform 1 0 9352 0 1 14112
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_163
timestamp 1698175906
transform 1 0 9800 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_172
timestamp 1698175906
transform 1 0 10304 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_174
timestamp 1698175906
transform 1 0 10416 0 1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_177
timestamp 1698175906
transform 1 0 10584 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_241
timestamp 1698175906
transform 1 0 14168 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_247
timestamp 1698175906
transform 1 0 14504 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_311
timestamp 1698175906
transform 1 0 18088 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_317
timestamp 1698175906
transform 1 0 18424 0 1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_2
timestamp 1698175906
transform 1 0 784 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_66
timestamp 1698175906
transform 1 0 4368 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_72
timestamp 1698175906
transform 1 0 4704 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_136
timestamp 1698175906
transform 1 0 8288 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_142
timestamp 1698175906
transform 1 0 8624 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_206
timestamp 1698175906
transform 1 0 12208 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_212
timestamp 1698175906
transform 1 0 12544 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_276
timestamp 1698175906
transform 1 0 16128 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_282
timestamp 1698175906
transform 1 0 16464 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_346
timestamp 1698175906
transform 1 0 20048 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_348
timestamp 1698175906
transform 1 0 20160 0 -1 14896
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698175906
transform 1 0 784 0 1 14896
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698175906
transform 1 0 2576 0 1 14896
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_37
timestamp 1698175906
transform 1 0 2744 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_101
timestamp 1698175906
transform 1 0 6328 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_107
timestamp 1698175906
transform 1 0 6664 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_171
timestamp 1698175906
transform 1 0 10248 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_177
timestamp 1698175906
transform 1 0 10584 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_241
timestamp 1698175906
transform 1 0 14168 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_247
timestamp 1698175906
transform 1 0 14504 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_311
timestamp 1698175906
transform 1 0 18088 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_317
timestamp 1698175906
transform 1 0 18424 0 1 14896
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2
timestamp 1698175906
transform 1 0 784 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_66
timestamp 1698175906
transform 1 0 4368 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_72
timestamp 1698175906
transform 1 0 4704 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_136
timestamp 1698175906
transform 1 0 8288 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_142
timestamp 1698175906
transform 1 0 8624 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_206
timestamp 1698175906
transform 1 0 12208 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_212
timestamp 1698175906
transform 1 0 12544 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_276
timestamp 1698175906
transform 1 0 16128 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_282
timestamp 1698175906
transform 1 0 16464 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_346
timestamp 1698175906
transform 1 0 20048 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_348
timestamp 1698175906
transform 1 0 20160 0 -1 15680
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_2
timestamp 1698175906
transform 1 0 784 0 1 15680
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698175906
transform 1 0 2576 0 1 15680
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_37
timestamp 1698175906
transform 1 0 2744 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_101
timestamp 1698175906
transform 1 0 6328 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_107
timestamp 1698175906
transform 1 0 6664 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_171
timestamp 1698175906
transform 1 0 10248 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_177
timestamp 1698175906
transform 1 0 10584 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_241
timestamp 1698175906
transform 1 0 14168 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_247
timestamp 1698175906
transform 1 0 14504 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_311
timestamp 1698175906
transform 1 0 18088 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_317
timestamp 1698175906
transform 1 0 18424 0 1 15680
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2
timestamp 1698175906
transform 1 0 784 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_66
timestamp 1698175906
transform 1 0 4368 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_72
timestamp 1698175906
transform 1 0 4704 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_136
timestamp 1698175906
transform 1 0 8288 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_142
timestamp 1698175906
transform 1 0 8624 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_206
timestamp 1698175906
transform 1 0 12208 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_212
timestamp 1698175906
transform 1 0 12544 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_276
timestamp 1698175906
transform 1 0 16128 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_282
timestamp 1698175906
transform 1 0 16464 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_346
timestamp 1698175906
transform 1 0 20048 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_348
timestamp 1698175906
transform 1 0 20160 0 -1 16464
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698175906
transform 1 0 784 0 1 16464
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698175906
transform 1 0 2576 0 1 16464
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_37
timestamp 1698175906
transform 1 0 2744 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_101
timestamp 1698175906
transform 1 0 6328 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_107
timestamp 1698175906
transform 1 0 6664 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_171
timestamp 1698175906
transform 1 0 10248 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_177
timestamp 1698175906
transform 1 0 10584 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_241
timestamp 1698175906
transform 1 0 14168 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_247
timestamp 1698175906
transform 1 0 14504 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_311
timestamp 1698175906
transform 1 0 18088 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_317
timestamp 1698175906
transform 1 0 18424 0 1 16464
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_2
timestamp 1698175906
transform 1 0 784 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_66
timestamp 1698175906
transform 1 0 4368 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_72
timestamp 1698175906
transform 1 0 4704 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_136
timestamp 1698175906
transform 1 0 8288 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_142
timestamp 1698175906
transform 1 0 8624 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_206
timestamp 1698175906
transform 1 0 12208 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_212
timestamp 1698175906
transform 1 0 12544 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_276
timestamp 1698175906
transform 1 0 16128 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_282
timestamp 1698175906
transform 1 0 16464 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_346
timestamp 1698175906
transform 1 0 20048 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_348
timestamp 1698175906
transform 1 0 20160 0 -1 17248
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698175906
transform 1 0 784 0 1 17248
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698175906
transform 1 0 2576 0 1 17248
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_37
timestamp 1698175906
transform 1 0 2744 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_101
timestamp 1698175906
transform 1 0 6328 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_107
timestamp 1698175906
transform 1 0 6664 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_171
timestamp 1698175906
transform 1 0 10248 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_177
timestamp 1698175906
transform 1 0 10584 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_241
timestamp 1698175906
transform 1 0 14168 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_247
timestamp 1698175906
transform 1 0 14504 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_311
timestamp 1698175906
transform 1 0 18088 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_317
timestamp 1698175906
transform 1 0 18424 0 1 17248
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2
timestamp 1698175906
transform 1 0 784 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1698175906
transform 1 0 4368 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_72
timestamp 1698175906
transform 1 0 4704 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_136
timestamp 1698175906
transform 1 0 8288 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_142
timestamp 1698175906
transform 1 0 8624 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_206
timestamp 1698175906
transform 1 0 12208 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_212
timestamp 1698175906
transform 1 0 12544 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_276
timestamp 1698175906
transform 1 0 16128 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_282
timestamp 1698175906
transform 1 0 16464 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_346
timestamp 1698175906
transform 1 0 20048 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_348
timestamp 1698175906
transform 1 0 20160 0 -1 18032
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_6
timestamp 1698175906
transform 1 0 1008 0 1 18032
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_22
timestamp 1698175906
transform 1 0 1904 0 1 18032
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_30
timestamp 1698175906
transform 1 0 2352 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698175906
transform 1 0 2576 0 1 18032
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_37
timestamp 1698175906
transform 1 0 2744 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_101
timestamp 1698175906
transform 1 0 6328 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_107
timestamp 1698175906
transform 1 0 6664 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_171
timestamp 1698175906
transform 1 0 10248 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_203
timestamp 1698175906
transform 1 0 12040 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_235
timestamp 1698175906
transform 1 0 13832 0 1 18032
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_243
timestamp 1698175906
transform 1 0 14280 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_247
timestamp 1698175906
transform 1 0 14504 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_311
timestamp 1698175906
transform 1 0 18088 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_317
timestamp 1698175906
transform 1 0 18424 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_2
timestamp 1698175906
transform 1 0 784 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_66
timestamp 1698175906
transform 1 0 4368 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_72
timestamp 1698175906
transform 1 0 4704 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_136
timestamp 1698175906
transform 1 0 8288 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_142
timestamp 1698175906
transform 1 0 8624 0 -1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_174
timestamp 1698175906
transform 1 0 10416 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_201
timestamp 1698175906
transform 1 0 11928 0 -1 18816
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_209
timestamp 1698175906
transform 1 0 12376 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_212
timestamp 1698175906
transform 1 0 12544 0 -1 18816
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_228
timestamp 1698175906
transform 1 0 13440 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_255
timestamp 1698175906
transform 1 0 14952 0 -1 18816
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_271
timestamp 1698175906
transform 1 0 15848 0 -1 18816
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_279
timestamp 1698175906
transform 1 0 16296 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_282
timestamp 1698175906
transform 1 0 16464 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_346
timestamp 1698175906
transform 1 0 20048 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_348
timestamp 1698175906
transform 1 0 20160 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_2
timestamp 1698175906
transform 1 0 784 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_36
timestamp 1698175906
transform 1 0 2688 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_70
timestamp 1698175906
transform 1 0 4592 0 1 18816
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_86
timestamp 1698175906
transform 1 0 5488 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_90
timestamp 1698175906
transform 1 0 5712 0 1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_95
timestamp 1698175906
transform 1 0 5992 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_99
timestamp 1698175906
transform 1 0 6216 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_101
timestamp 1698175906
transform 1 0 6328 0 1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_104
timestamp 1698175906
transform 1 0 6496 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_138
timestamp 1698175906
transform 1 0 8400 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_142
timestamp 1698175906
transform 1 0 8624 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_172
timestamp 1698175906
transform 1 0 10304 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_176
timestamp 1698175906
transform 1 0 10528 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_232
timestamp 1698175906
transform 1 0 13664 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_236
timestamp 1698175906
transform 1 0 13888 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_240
timestamp 1698175906
transform 1 0 14112 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_274
timestamp 1698175906
transform 1 0 16016 0 1 18816
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_290
timestamp 1698175906
transform 1 0 16912 0 1 18816
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_298
timestamp 1698175906
transform 1 0 17360 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_300
timestamp 1698175906
transform 1 0 17472 0 1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_305
timestamp 1698175906
transform 1 0 17752 0 1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_308
timestamp 1698175906
transform 1 0 17920 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_342
timestamp 1698175906
transform 1 0 19824 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_346
timestamp 1698175906
transform 1 0 20048 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_348
timestamp 1698175906
transform 1 0 20160 0 1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita51_24 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 5992 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita51_25
timestamp 1698175906
transform -1 0 1008 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita51_26
timestamp 1698175906
transform -1 0 17752 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18760 0 -1 10192
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output2
timestamp 1698175906
transform -1 0 10192 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output3
timestamp 1698175906
transform -1 0 2240 0 1 7840
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output4
timestamp 1698175906
transform 1 0 8456 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output5
timestamp 1698175906
transform 1 0 18760 0 -1 11760
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output6
timestamp 1698175906
transform 1 0 10584 0 1 18032
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output7
timestamp 1698175906
transform 1 0 18760 0 1 11760
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output8
timestamp 1698175906
transform 1 0 18760 0 -1 10976
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output9
timestamp 1698175906
transform -1 0 2240 0 -1 10976
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output10
timestamp 1698175906
transform 1 0 18760 0 -1 8624
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output11
timestamp 1698175906
transform 1 0 18760 0 1 8624
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output12
timestamp 1698175906
transform -1 0 2240 0 1 10192
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output13
timestamp 1698175906
transform 1 0 18760 0 1 10976
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output14
timestamp 1698175906
transform 1 0 12544 0 -1 2352
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output15
timestamp 1698175906
transform -1 0 12096 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output16
timestamp 1698175906
transform 1 0 13496 0 -1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output17
timestamp 1698175906
transform 1 0 10472 0 -1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output18
timestamp 1698175906
transform 1 0 12208 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output19
timestamp 1698175906
transform 1 0 10640 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output20
timestamp 1698175906
transform 1 0 9464 0 -1 2352
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output21
timestamp 1698175906
transform -1 0 2240 0 -1 12544
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output22
timestamp 1698175906
transform 1 0 18760 0 1 13328
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output23
timestamp 1698175906
transform 1 0 12208 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_45 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 672 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698175906
transform -1 0 20328 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_46
timestamp 1698175906
transform 1 0 672 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698175906
transform -1 0 20328 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_47
timestamp 1698175906
transform 1 0 672 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698175906
transform -1 0 20328 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_48
timestamp 1698175906
transform 1 0 672 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698175906
transform -1 0 20328 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_49
timestamp 1698175906
transform 1 0 672 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698175906
transform -1 0 20328 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_50
timestamp 1698175906
transform 1 0 672 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698175906
transform -1 0 20328 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_51
timestamp 1698175906
transform 1 0 672 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698175906
transform -1 0 20328 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_52
timestamp 1698175906
transform 1 0 672 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698175906
transform -1 0 20328 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_53
timestamp 1698175906
transform 1 0 672 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698175906
transform -1 0 20328 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_54
timestamp 1698175906
transform 1 0 672 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698175906
transform -1 0 20328 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_55
timestamp 1698175906
transform 1 0 672 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698175906
transform -1 0 20328 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_56
timestamp 1698175906
transform 1 0 672 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698175906
transform -1 0 20328 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_57
timestamp 1698175906
transform 1 0 672 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698175906
transform -1 0 20328 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_58
timestamp 1698175906
transform 1 0 672 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698175906
transform -1 0 20328 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_59
timestamp 1698175906
transform 1 0 672 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698175906
transform -1 0 20328 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_60
timestamp 1698175906
transform 1 0 672 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698175906
transform -1 0 20328 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_61
timestamp 1698175906
transform 1 0 672 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698175906
transform -1 0 20328 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_62
timestamp 1698175906
transform 1 0 672 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698175906
transform -1 0 20328 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_63
timestamp 1698175906
transform 1 0 672 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698175906
transform -1 0 20328 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_64
timestamp 1698175906
transform 1 0 672 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698175906
transform -1 0 20328 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_65
timestamp 1698175906
transform 1 0 672 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698175906
transform -1 0 20328 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_66
timestamp 1698175906
transform 1 0 672 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698175906
transform -1 0 20328 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_67
timestamp 1698175906
transform 1 0 672 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698175906
transform -1 0 20328 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_68
timestamp 1698175906
transform 1 0 672 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698175906
transform -1 0 20328 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_69
timestamp 1698175906
transform 1 0 672 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698175906
transform -1 0 20328 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_70
timestamp 1698175906
transform 1 0 672 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698175906
transform -1 0 20328 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_71
timestamp 1698175906
transform 1 0 672 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698175906
transform -1 0 20328 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_72
timestamp 1698175906
transform 1 0 672 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698175906
transform -1 0 20328 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_73
timestamp 1698175906
transform 1 0 672 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698175906
transform -1 0 20328 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_74
timestamp 1698175906
transform 1 0 672 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698175906
transform -1 0 20328 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_75
timestamp 1698175906
transform 1 0 672 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698175906
transform -1 0 20328 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_76
timestamp 1698175906
transform 1 0 672 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698175906
transform -1 0 20328 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_77
timestamp 1698175906
transform 1 0 672 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698175906
transform -1 0 20328 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_78
timestamp 1698175906
transform 1 0 672 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698175906
transform -1 0 20328 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_79
timestamp 1698175906
transform 1 0 672 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698175906
transform -1 0 20328 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_80
timestamp 1698175906
transform 1 0 672 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698175906
transform -1 0 20328 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_81
timestamp 1698175906
transform 1 0 672 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698175906
transform -1 0 20328 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_82
timestamp 1698175906
transform 1 0 672 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698175906
transform -1 0 20328 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_83
timestamp 1698175906
transform 1 0 672 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698175906
transform -1 0 20328 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_84
timestamp 1698175906
transform 1 0 672 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698175906
transform -1 0 20328 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_85
timestamp 1698175906
transform 1 0 672 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698175906
transform -1 0 20328 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_86
timestamp 1698175906
transform 1 0 672 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698175906
transform -1 0 20328 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_87
timestamp 1698175906
transform 1 0 672 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698175906
transform -1 0 20328 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_88
timestamp 1698175906
transform 1 0 672 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698175906
transform -1 0 20328 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_89
timestamp 1698175906
transform 1 0 672 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698175906
transform -1 0 20328 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_90 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 2576 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_91
timestamp 1698175906
transform 1 0 4480 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_92
timestamp 1698175906
transform 1 0 6384 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_93
timestamp 1698175906
transform 1 0 8288 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_94
timestamp 1698175906
transform 1 0 10192 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_95
timestamp 1698175906
transform 1 0 12096 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_96
timestamp 1698175906
transform 1 0 14000 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_97
timestamp 1698175906
transform 1 0 15904 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_98
timestamp 1698175906
transform 1 0 17808 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_99
timestamp 1698175906
transform 1 0 19712 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_100
timestamp 1698175906
transform 1 0 4592 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_101
timestamp 1698175906
transform 1 0 8512 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_102
timestamp 1698175906
transform 1 0 12432 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_103
timestamp 1698175906
transform 1 0 16352 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_104
timestamp 1698175906
transform 1 0 2632 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_105
timestamp 1698175906
transform 1 0 6552 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_106
timestamp 1698175906
transform 1 0 10472 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_107
timestamp 1698175906
transform 1 0 14392 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_108
timestamp 1698175906
transform 1 0 18312 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_109
timestamp 1698175906
transform 1 0 4592 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_110
timestamp 1698175906
transform 1 0 8512 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_111
timestamp 1698175906
transform 1 0 12432 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_112
timestamp 1698175906
transform 1 0 16352 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_113
timestamp 1698175906
transform 1 0 2632 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_114
timestamp 1698175906
transform 1 0 6552 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_115
timestamp 1698175906
transform 1 0 10472 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_116
timestamp 1698175906
transform 1 0 14392 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_117
timestamp 1698175906
transform 1 0 18312 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_118
timestamp 1698175906
transform 1 0 4592 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_119
timestamp 1698175906
transform 1 0 8512 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_120
timestamp 1698175906
transform 1 0 12432 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_121
timestamp 1698175906
transform 1 0 16352 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_122
timestamp 1698175906
transform 1 0 2632 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_123
timestamp 1698175906
transform 1 0 6552 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_124
timestamp 1698175906
transform 1 0 10472 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_125
timestamp 1698175906
transform 1 0 14392 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_126
timestamp 1698175906
transform 1 0 18312 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_127
timestamp 1698175906
transform 1 0 4592 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_128
timestamp 1698175906
transform 1 0 8512 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_129
timestamp 1698175906
transform 1 0 12432 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_130
timestamp 1698175906
transform 1 0 16352 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_131
timestamp 1698175906
transform 1 0 2632 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_132
timestamp 1698175906
transform 1 0 6552 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_133
timestamp 1698175906
transform 1 0 10472 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_134
timestamp 1698175906
transform 1 0 14392 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_135
timestamp 1698175906
transform 1 0 18312 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_136
timestamp 1698175906
transform 1 0 4592 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_137
timestamp 1698175906
transform 1 0 8512 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_138
timestamp 1698175906
transform 1 0 12432 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_139
timestamp 1698175906
transform 1 0 16352 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_140
timestamp 1698175906
transform 1 0 2632 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_141
timestamp 1698175906
transform 1 0 6552 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_142
timestamp 1698175906
transform 1 0 10472 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_143
timestamp 1698175906
transform 1 0 14392 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_144
timestamp 1698175906
transform 1 0 18312 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_145
timestamp 1698175906
transform 1 0 4592 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_146
timestamp 1698175906
transform 1 0 8512 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_147
timestamp 1698175906
transform 1 0 12432 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_148
timestamp 1698175906
transform 1 0 16352 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_149
timestamp 1698175906
transform 1 0 2632 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_150
timestamp 1698175906
transform 1 0 6552 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_151
timestamp 1698175906
transform 1 0 10472 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_152
timestamp 1698175906
transform 1 0 14392 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_153
timestamp 1698175906
transform 1 0 18312 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_154
timestamp 1698175906
transform 1 0 4592 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_155
timestamp 1698175906
transform 1 0 8512 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_156
timestamp 1698175906
transform 1 0 12432 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_157
timestamp 1698175906
transform 1 0 16352 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_158
timestamp 1698175906
transform 1 0 2632 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_159
timestamp 1698175906
transform 1 0 6552 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_160
timestamp 1698175906
transform 1 0 10472 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_161
timestamp 1698175906
transform 1 0 14392 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_162
timestamp 1698175906
transform 1 0 18312 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_163
timestamp 1698175906
transform 1 0 4592 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_164
timestamp 1698175906
transform 1 0 8512 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_165
timestamp 1698175906
transform 1 0 12432 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_166
timestamp 1698175906
transform 1 0 16352 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_167
timestamp 1698175906
transform 1 0 2632 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_168
timestamp 1698175906
transform 1 0 6552 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_169
timestamp 1698175906
transform 1 0 10472 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_170
timestamp 1698175906
transform 1 0 14392 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_171
timestamp 1698175906
transform 1 0 18312 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_172
timestamp 1698175906
transform 1 0 4592 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_173
timestamp 1698175906
transform 1 0 8512 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_174
timestamp 1698175906
transform 1 0 12432 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_175
timestamp 1698175906
transform 1 0 16352 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_176
timestamp 1698175906
transform 1 0 2632 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_177
timestamp 1698175906
transform 1 0 6552 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_178
timestamp 1698175906
transform 1 0 10472 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_179
timestamp 1698175906
transform 1 0 14392 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_180
timestamp 1698175906
transform 1 0 18312 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_181
timestamp 1698175906
transform 1 0 4592 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_182
timestamp 1698175906
transform 1 0 8512 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_183
timestamp 1698175906
transform 1 0 12432 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_184
timestamp 1698175906
transform 1 0 16352 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_185
timestamp 1698175906
transform 1 0 2632 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_186
timestamp 1698175906
transform 1 0 6552 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_187
timestamp 1698175906
transform 1 0 10472 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_188
timestamp 1698175906
transform 1 0 14392 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_189
timestamp 1698175906
transform 1 0 18312 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_190
timestamp 1698175906
transform 1 0 4592 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_191
timestamp 1698175906
transform 1 0 8512 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_192
timestamp 1698175906
transform 1 0 12432 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_193
timestamp 1698175906
transform 1 0 16352 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_194
timestamp 1698175906
transform 1 0 2632 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_195
timestamp 1698175906
transform 1 0 6552 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_196
timestamp 1698175906
transform 1 0 10472 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_197
timestamp 1698175906
transform 1 0 14392 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_198
timestamp 1698175906
transform 1 0 18312 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_199
timestamp 1698175906
transform 1 0 4592 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_200
timestamp 1698175906
transform 1 0 8512 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_201
timestamp 1698175906
transform 1 0 12432 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_202
timestamp 1698175906
transform 1 0 16352 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_203
timestamp 1698175906
transform 1 0 2632 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_204
timestamp 1698175906
transform 1 0 6552 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_205
timestamp 1698175906
transform 1 0 10472 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_206
timestamp 1698175906
transform 1 0 14392 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_207
timestamp 1698175906
transform 1 0 18312 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_208
timestamp 1698175906
transform 1 0 4592 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_209
timestamp 1698175906
transform 1 0 8512 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_210
timestamp 1698175906
transform 1 0 12432 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_211
timestamp 1698175906
transform 1 0 16352 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_212
timestamp 1698175906
transform 1 0 2632 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_213
timestamp 1698175906
transform 1 0 6552 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_214
timestamp 1698175906
transform 1 0 10472 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_215
timestamp 1698175906
transform 1 0 14392 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_216
timestamp 1698175906
transform 1 0 18312 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_217
timestamp 1698175906
transform 1 0 4592 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_218
timestamp 1698175906
transform 1 0 8512 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_219
timestamp 1698175906
transform 1 0 12432 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_220
timestamp 1698175906
transform 1 0 16352 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_221
timestamp 1698175906
transform 1 0 2632 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_222
timestamp 1698175906
transform 1 0 6552 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_223
timestamp 1698175906
transform 1 0 10472 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_224
timestamp 1698175906
transform 1 0 14392 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_225
timestamp 1698175906
transform 1 0 18312 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_226
timestamp 1698175906
transform 1 0 4592 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_227
timestamp 1698175906
transform 1 0 8512 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_228
timestamp 1698175906
transform 1 0 12432 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_229
timestamp 1698175906
transform 1 0 16352 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_230
timestamp 1698175906
transform 1 0 2632 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_231
timestamp 1698175906
transform 1 0 6552 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_232
timestamp 1698175906
transform 1 0 10472 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_233
timestamp 1698175906
transform 1 0 14392 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_234
timestamp 1698175906
transform 1 0 18312 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_235
timestamp 1698175906
transform 1 0 4592 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_236
timestamp 1698175906
transform 1 0 8512 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_237
timestamp 1698175906
transform 1 0 12432 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_238
timestamp 1698175906
transform 1 0 16352 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_239
timestamp 1698175906
transform 1 0 2632 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_240
timestamp 1698175906
transform 1 0 6552 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_241
timestamp 1698175906
transform 1 0 10472 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_242
timestamp 1698175906
transform 1 0 14392 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_243
timestamp 1698175906
transform 1 0 18312 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_244
timestamp 1698175906
transform 1 0 4592 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_245
timestamp 1698175906
transform 1 0 8512 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_246
timestamp 1698175906
transform 1 0 12432 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_247
timestamp 1698175906
transform 1 0 16352 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_248
timestamp 1698175906
transform 1 0 2632 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_249
timestamp 1698175906
transform 1 0 6552 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_250
timestamp 1698175906
transform 1 0 10472 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_251
timestamp 1698175906
transform 1 0 14392 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_252
timestamp 1698175906
transform 1 0 18312 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_253
timestamp 1698175906
transform 1 0 4592 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_254
timestamp 1698175906
transform 1 0 8512 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_255
timestamp 1698175906
transform 1 0 12432 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_256
timestamp 1698175906
transform 1 0 16352 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_257
timestamp 1698175906
transform 1 0 2632 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_258
timestamp 1698175906
transform 1 0 6552 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_259
timestamp 1698175906
transform 1 0 10472 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_260
timestamp 1698175906
transform 1 0 14392 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_261
timestamp 1698175906
transform 1 0 18312 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_262
timestamp 1698175906
transform 1 0 4592 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_263
timestamp 1698175906
transform 1 0 8512 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_264
timestamp 1698175906
transform 1 0 12432 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_265
timestamp 1698175906
transform 1 0 16352 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_266
timestamp 1698175906
transform 1 0 2632 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_267
timestamp 1698175906
transform 1 0 6552 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_268
timestamp 1698175906
transform 1 0 10472 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_269
timestamp 1698175906
transform 1 0 14392 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_270
timestamp 1698175906
transform 1 0 18312 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_271
timestamp 1698175906
transform 1 0 4592 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_272
timestamp 1698175906
transform 1 0 8512 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_273
timestamp 1698175906
transform 1 0 12432 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_274
timestamp 1698175906
transform 1 0 16352 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_275
timestamp 1698175906
transform 1 0 2632 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_276
timestamp 1698175906
transform 1 0 6552 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_277
timestamp 1698175906
transform 1 0 10472 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_278
timestamp 1698175906
transform 1 0 14392 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_279
timestamp 1698175906
transform 1 0 18312 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_280
timestamp 1698175906
transform 1 0 4592 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_281
timestamp 1698175906
transform 1 0 8512 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_282
timestamp 1698175906
transform 1 0 12432 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_283
timestamp 1698175906
transform 1 0 16352 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_284
timestamp 1698175906
transform 1 0 2632 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_285
timestamp 1698175906
transform 1 0 6552 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_286
timestamp 1698175906
transform 1 0 10472 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_287
timestamp 1698175906
transform 1 0 14392 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_288
timestamp 1698175906
transform 1 0 18312 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_289
timestamp 1698175906
transform 1 0 4592 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_290
timestamp 1698175906
transform 1 0 8512 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_291
timestamp 1698175906
transform 1 0 12432 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_292
timestamp 1698175906
transform 1 0 16352 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_293
timestamp 1698175906
transform 1 0 2576 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_294
timestamp 1698175906
transform 1 0 4480 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_295
timestamp 1698175906
transform 1 0 6384 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_296
timestamp 1698175906
transform 1 0 8288 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_297
timestamp 1698175906
transform 1 0 10192 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_298
timestamp 1698175906
transform 1 0 12096 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_299
timestamp 1698175906
transform 1 0 14000 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_300
timestamp 1698175906
transform 1 0 15904 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_301
timestamp 1698175906
transform 1 0 17808 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_302
timestamp 1698175906
transform 1 0 19712 0 1 18816
box -43 -43 155 435
<< labels >>
flabel metal3 s 0 13776 400 13832 0 FreeSans 224 0 0 0 clk
port 0 nsew signal input
flabel metal2 s 5712 20600 5768 21000 0 FreeSans 224 90 0 0 segm[0]
port 1 nsew signal tristate
flabel metal3 s 20600 9744 21000 9800 0 FreeSans 224 0 0 0 segm[10]
port 2 nsew signal tristate
flabel metal2 s 9072 20600 9128 21000 0 FreeSans 224 90 0 0 segm[11]
port 3 nsew signal tristate
flabel metal3 s 0 7728 400 7784 0 FreeSans 224 0 0 0 segm[12]
port 4 nsew signal tristate
flabel metal2 s 8400 0 8456 400 0 FreeSans 224 90 0 0 segm[13]
port 5 nsew signal tristate
flabel metal3 s 20600 11424 21000 11480 0 FreeSans 224 0 0 0 segm[1]
port 6 nsew signal tristate
flabel metal2 s 10080 20600 10136 21000 0 FreeSans 224 90 0 0 segm[2]
port 7 nsew signal tristate
flabel metal3 s 0 18144 400 18200 0 FreeSans 224 0 0 0 segm[3]
port 8 nsew signal tristate
flabel metal3 s 20600 11760 21000 11816 0 FreeSans 224 0 0 0 segm[4]
port 9 nsew signal tristate
flabel metal2 s 17472 20600 17528 21000 0 FreeSans 224 90 0 0 segm[5]
port 10 nsew signal tristate
flabel metal3 s 20600 10752 21000 10808 0 FreeSans 224 0 0 0 segm[6]
port 11 nsew signal tristate
flabel metal3 s 0 10416 400 10472 0 FreeSans 224 0 0 0 segm[7]
port 12 nsew signal tristate
flabel metal3 s 20600 8400 21000 8456 0 FreeSans 224 0 0 0 segm[8]
port 13 nsew signal tristate
flabel metal3 s 20600 8736 21000 8792 0 FreeSans 224 0 0 0 segm[9]
port 14 nsew signal tristate
flabel metal3 s 0 10080 400 10136 0 FreeSans 224 0 0 0 sel[0]
port 15 nsew signal tristate
flabel metal3 s 20600 11088 21000 11144 0 FreeSans 224 0 0 0 sel[10]
port 16 nsew signal tristate
flabel metal2 s 12432 0 12488 400 0 FreeSans 224 90 0 0 sel[11]
port 17 nsew signal tristate
flabel metal2 s 11088 20600 11144 21000 0 FreeSans 224 90 0 0 sel[1]
port 18 nsew signal tristate
flabel metal2 s 13440 20600 13496 21000 0 FreeSans 224 90 0 0 sel[2]
port 19 nsew signal tristate
flabel metal2 s 10416 20600 10472 21000 0 FreeSans 224 90 0 0 sel[3]
port 20 nsew signal tristate
flabel metal2 s 11424 20600 11480 21000 0 FreeSans 224 90 0 0 sel[4]
port 21 nsew signal tristate
flabel metal2 s 11088 0 11144 400 0 FreeSans 224 90 0 0 sel[5]
port 22 nsew signal tristate
flabel metal2 s 9408 0 9464 400 0 FreeSans 224 90 0 0 sel[6]
port 23 nsew signal tristate
flabel metal3 s 0 12096 400 12152 0 FreeSans 224 0 0 0 sel[7]
port 24 nsew signal tristate
flabel metal3 s 20600 13104 21000 13160 0 FreeSans 224 0 0 0 sel[8]
port 25 nsew signal tristate
flabel metal2 s 11424 0 11480 400 0 FreeSans 224 90 0 0 sel[9]
port 26 nsew signal tristate
flabel metal4 s 2224 1538 2384 19238 0 FreeSans 640 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 17584 1538 17744 19238 0 FreeSans 640 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 9904 1538 10064 19238 0 FreeSans 640 90 0 0 vss
port 28 nsew ground bidirectional
rlabel metal1 10500 19208 10500 19208 0 vdd
rlabel metal1 10500 18816 10500 18816 0 vss
rlabel metal3 8764 7196 8764 7196 0 _000_
rlabel metal2 8092 9380 8092 9380 0 _001_
rlabel metal2 7840 8876 7840 8876 0 _002_
rlabel metal3 8540 11676 8540 11676 0 _003_
rlabel metal2 7980 11368 7980 11368 0 _004_
rlabel metal2 10864 6132 10864 6132 0 _005_
rlabel metal2 10668 13692 10668 13692 0 _006_
rlabel metal2 9212 13748 9212 13748 0 _007_
rlabel metal2 12348 13020 12348 13020 0 _008_
rlabel metal2 11060 12376 11060 12376 0 _009_
rlabel metal3 7000 10108 7000 10108 0 _010_
rlabel metal2 13468 11368 13468 11368 0 _011_
rlabel metal2 13020 10584 13020 10584 0 _012_
rlabel metal2 6076 10556 6076 10556 0 _013_
rlabel metal2 12964 12964 12964 12964 0 _014_
rlabel metal2 11956 11004 11956 11004 0 _015_
rlabel metal2 12264 7308 12264 7308 0 _016_
rlabel metal3 12348 8764 12348 8764 0 _017_
rlabel metal2 12124 9352 12124 9352 0 _018_
rlabel metal3 8288 13244 8288 13244 0 _019_
rlabel metal3 6664 7644 6664 7644 0 _020_
rlabel metal2 7252 7028 7252 7028 0 _021_
rlabel metal2 10640 6916 10640 6916 0 _022_
rlabel metal2 6692 12124 6692 12124 0 _023_
rlabel metal2 13552 11900 13552 11900 0 _024_
rlabel metal2 11396 10752 11396 10752 0 _025_
rlabel metal2 11116 12152 11116 12152 0 _026_
rlabel metal2 7476 10304 7476 10304 0 _027_
rlabel metal2 11340 9828 11340 9828 0 _028_
rlabel metal2 11116 9156 11116 9156 0 _029_
rlabel metal2 13356 11200 13356 11200 0 _030_
rlabel metal2 13524 11396 13524 11396 0 _031_
rlabel metal2 13188 10416 13188 10416 0 _032_
rlabel metal2 13468 10416 13468 10416 0 _033_
rlabel metal2 9996 8932 9996 8932 0 _034_
rlabel metal2 10052 8792 10052 8792 0 _035_
rlabel metal2 10304 8820 10304 8820 0 _036_
rlabel metal2 9940 8960 9940 8960 0 _037_
rlabel metal3 6608 10892 6608 10892 0 _038_
rlabel metal2 6860 10640 6860 10640 0 _039_
rlabel metal2 13328 12628 13328 12628 0 _040_
rlabel metal2 9492 10752 9492 10752 0 _041_
rlabel metal3 9548 10528 9548 10528 0 _042_
rlabel metal2 11788 10752 11788 10752 0 _043_
rlabel metal2 11956 10080 11956 10080 0 _044_
rlabel metal2 10444 7644 10444 7644 0 _045_
rlabel metal2 12488 8092 12488 8092 0 _046_
rlabel metal3 11312 8876 11312 8876 0 _047_
rlabel metal3 12264 8372 12264 8372 0 _048_
rlabel metal2 11424 10388 11424 10388 0 _049_
rlabel metal2 11956 9240 11956 9240 0 _050_
rlabel metal2 9100 11228 9100 11228 0 _051_
rlabel metal2 9436 13132 9436 13132 0 _052_
rlabel metal3 7238 7700 7238 7700 0 _053_
rlabel metal2 6860 7812 6860 7812 0 _054_
rlabel metal2 7700 7336 7700 7336 0 _055_
rlabel metal2 9128 9156 9128 9156 0 _056_
rlabel metal2 9660 8988 9660 8988 0 _057_
rlabel metal2 9268 9352 9268 9352 0 _058_
rlabel via2 9324 7980 9324 7980 0 _059_
rlabel metal2 10752 8036 10752 8036 0 _060_
rlabel metal2 10752 11956 10752 11956 0 _061_
rlabel metal2 10724 10500 10724 10500 0 _062_
rlabel metal2 10108 11144 10108 11144 0 _063_
rlabel metal2 11900 9968 11900 9968 0 _064_
rlabel metal2 9044 11312 9044 11312 0 _065_
rlabel metal2 9156 11004 9156 11004 0 _066_
rlabel metal3 10696 7196 10696 7196 0 _067_
rlabel metal2 11172 7462 11172 7462 0 _068_
rlabel metal2 9716 12124 9716 12124 0 _069_
rlabel metal2 7140 11984 7140 11984 0 _070_
rlabel metal2 6804 11816 6804 11816 0 _071_
rlabel metal3 9772 9548 9772 9548 0 _072_
rlabel metal2 8260 10976 8260 10976 0 _073_
rlabel metal2 11564 9072 11564 9072 0 _074_
rlabel metal2 9772 9156 9772 9156 0 _075_
rlabel metal2 8904 10780 8904 10780 0 _076_
rlabel metal3 6860 11816 6860 11816 0 _077_
rlabel metal2 9660 10052 9660 10052 0 _078_
rlabel metal2 10668 8904 10668 8904 0 _079_
rlabel metal2 9884 8876 9884 8876 0 _080_
rlabel metal2 9044 7252 9044 7252 0 _081_
rlabel metal2 7728 8428 7728 8428 0 _082_
rlabel metal3 10948 10276 10948 10276 0 _083_
rlabel metal2 10220 10556 10220 10556 0 _084_
rlabel metal3 8764 10052 8764 10052 0 _085_
rlabel metal2 7140 10220 7140 10220 0 _086_
rlabel metal2 9268 13706 9268 13706 0 _087_
rlabel metal2 10528 7252 10528 7252 0 _088_
rlabel metal2 7252 9968 7252 9968 0 _089_
rlabel metal2 10780 13300 10780 13300 0 _090_
rlabel metal2 13048 13916 13048 13916 0 _091_
rlabel metal2 10920 13468 10920 13468 0 _092_
rlabel metal2 9324 14140 9324 14140 0 _093_
rlabel metal2 9436 9436 9436 9436 0 _094_
rlabel metal2 12796 11312 12796 11312 0 _095_
rlabel metal3 12656 13804 12656 13804 0 _096_
rlabel metal3 1239 13804 1239 13804 0 clk
rlabel metal3 10080 9940 10080 9940 0 clknet_0_clk
rlabel metal2 11648 7308 11648 7308 0 clknet_1_0__leaf_clk
rlabel metal2 7084 10556 7084 10556 0 clknet_1_1__leaf_clk
rlabel metal2 7476 9184 7476 9184 0 dut51.count\[0\]
rlabel metal3 8484 9212 8484 9212 0 dut51.count\[1\]
rlabel metal2 9716 10864 9716 10864 0 dut51.count\[2\]
rlabel metal3 8764 11564 8764 11564 0 dut51.count\[3\]
rlabel metal2 13748 9996 13748 9996 0 net1
rlabel metal2 18956 8568 18956 8568 0 net10
rlabel metal2 13916 8736 13916 8736 0 net11
rlabel metal3 3178 10388 3178 10388 0 net12
rlabel metal3 15960 11116 15960 11116 0 net13
rlabel metal3 12488 7700 12488 7700 0 net14
rlabel metal2 12012 17486 12012 17486 0 net15
rlabel metal3 13216 14028 13216 14028 0 net16
rlabel metal2 10556 16324 10556 16324 0 net17
rlabel metal3 11956 13860 11956 13860 0 net18
rlabel metal2 10332 6552 10332 6552 0 net19
rlabel metal3 9128 13580 9128 13580 0 net2
rlabel metal3 9352 6916 9352 6916 0 net20
rlabel metal2 5628 12320 5628 12320 0 net21
rlabel metal2 18844 13300 18844 13300 0 net22
rlabel metal2 11620 6776 11620 6776 0 net23
rlabel metal2 5796 18956 5796 18956 0 net24
rlabel metal3 623 18172 623 18172 0 net25
rlabel metal2 17556 18956 17556 18956 0 net26
rlabel metal2 5236 7812 5236 7812 0 net3
rlabel metal2 8540 2982 8540 2982 0 net4
rlabel metal3 15302 11620 15302 11620 0 net5
rlabel metal2 10276 13860 10276 13860 0 net6
rlabel metal2 14532 11760 14532 11760 0 net7
rlabel metal2 13636 10528 13636 10528 0 net8
rlabel metal3 3178 10780 3178 10780 0 net9
rlabel metal2 20020 9828 20020 9828 0 segm[10]
rlabel metal2 9100 19845 9100 19845 0 segm[11]
rlabel metal3 679 7756 679 7756 0 segm[12]
rlabel metal2 8428 1043 8428 1043 0 segm[13]
rlabel metal3 20321 11452 20321 11452 0 segm[1]
rlabel metal2 10108 19481 10108 19481 0 segm[2]
rlabel metal2 20020 11900 20020 11900 0 segm[4]
rlabel metal2 20020 10752 20020 10752 0 segm[6]
rlabel metal3 679 10444 679 10444 0 segm[7]
rlabel metal2 20020 8400 20020 8400 0 segm[8]
rlabel metal2 20020 8820 20020 8820 0 segm[9]
rlabel metal3 707 10108 707 10108 0 sel[0]
rlabel metal2 20020 11172 20020 11172 0 sel[10]
rlabel metal2 12460 1211 12460 1211 0 sel[11]
rlabel metal2 11116 19845 11116 19845 0 sel[1]
rlabel metal2 13468 19677 13468 19677 0 sel[2]
rlabel metal2 10444 19677 10444 19677 0 sel[3]
rlabel metal2 11452 19873 11452 19873 0 sel[4]
rlabel metal2 11116 1015 11116 1015 0 sel[5]
rlabel metal2 9436 1211 9436 1211 0 sel[6]
rlabel metal3 679 12124 679 12124 0 sel[7]
rlabel metal2 20020 13356 20020 13356 0 sel[8]
rlabel metal2 11452 1099 11452 1099 0 sel[9]
<< properties >>
string FIXED_BBOX 0 0 21000 21000
<< end >>
