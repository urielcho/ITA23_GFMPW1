// This is the unpowered netlist.
module user_proj_example (wb_clk_i,
    wb_rst_i,
    wbs_ack_o,
    wbs_cyc_i,
    wbs_stb_i,
    wbs_we_i,
    io_in,
    io_oeb,
    io_out,
    irq,
    la_data_in,
    la_data_out,
    la_oenb,
    wbs_adr_i,
    wbs_dat_i,
    wbs_dat_o,
    wbs_sel_i);
 input wb_clk_i;
 input wb_rst_i;
 output wbs_ack_o;
 input wbs_cyc_i;
 input wbs_stb_i;
 input wbs_we_i;
 input [15:0] io_in;
 output [15:0] io_oeb;
 output [15:0] io_out;
 output [2:0] irq;
 input [63:0] la_data_in;
 output [63:0] la_data_out;
 input [63:0] la_oenb;
 input [31:0] wbs_adr_i;
 input [31:0] wbs_dat_i;
 output [31:0] wbs_dat_o;
 input [3:0] wbs_sel_i;

 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire \clknet_0_counter.clk ;
 wire \clknet_2_0__leaf_counter.clk ;
 wire \clknet_2_1__leaf_counter.clk ;
 wire \clknet_2_2__leaf_counter.clk ;
 wire \clknet_2_3__leaf_counter.clk ;
 wire \counter.clk ;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;

 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_1 (.I(net140));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__170__I0 (.I(net278));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__170__I1 (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__170__S (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__172__I1 (.I(wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__174__I (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__176__I (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__179__A1 (.I(net107));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__179__A2 (.I(_039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__180__A2 (.I(_040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__184__I (.I(_043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__186__A1 (.I(net107));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__186__A2 (.I(_039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__188__A2 (.I(_047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__194__A1 (.I(_052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__194__A2 (.I(_053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__195__B (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__197__A1 (.I(_055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__197__A2 (.I(_056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__198__I (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__199__I (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__205__B (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__206__A4 (.I(_065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__208__B (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__210__A1 (.I(_067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__210__A2 (.I(_068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__210__A3 (.I(_069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__210__A4 (.I(_045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__215__A1 (.I(_071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__215__A3 (.I(_073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__215__A4 (.I(_074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__217__A1 (.I(_040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__218__A1 (.I(_040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__218__A2 (.I(_047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__220__I (.I(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__222__A2 (.I(_045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__222__B2 (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__222__C2 (.I(_081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__225__I (.I(net82));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__226__A2 (.I(_084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__227__A2 (.I(_053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__227__C2 (.I(net46));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__229__A2 (.I(_084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__230__A1 (.I(net136));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__231__C2 (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__233__A2 (.I(_084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__233__A3 (.I(net136));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__234__A1 (.I(net135));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__235__C2 (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__237__I (.I(_043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__238__A1 (.I(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__238__A2 (.I(net82));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__238__A3 (.I(net137));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__238__A4 (.I(net135));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__239__A1 (.I(net133));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__241__A2 (.I(_055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__241__C2 (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__243__A1 (.I(net133));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__243__A2 (.I(net132));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__245__A1 (.I(net134));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__245__B (.I(net132));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__247__A2 (.I(_056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__247__C2 (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__249__A1 (.I(net130));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__250__A2 (.I(_052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__250__C2 (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__252__A1 (.I(net130));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__253__A1 (.I(net129));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__254__C2 (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__256__I (.I(_043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__258__A2 (.I(_109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__261__I (.I(net89));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__262__A1 (.I(net131));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__262__A2 (.I(net129));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__263__I (.I(_114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__265__A1 (.I(_040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__265__A2 (.I(_109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__267__A1 (.I(net262));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__267__A2 (.I(_068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__267__C1 (.I(_118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__270__A1 (.I(net89));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__270__A2 (.I(net128));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__271__A1 (.I(net128));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__272__A2 (.I(_069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__272__B1 (.I(_118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__277__A1 (.I(net270));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__277__A2 (.I(_074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__277__C2 (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__279__B (.I(net77));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__281__I (.I(net77));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__282__A3 (.I(_114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__283__A2 (.I(_131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__284__A1 (.I(net266));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__284__A2 (.I(_067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__286__A1 (.I(net124));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__286__A2 (.I(_131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__287__A1 (.I(net274));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__287__A2 (.I(_073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__287__C2 (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__289__I (.I(net79));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__290__A1 (.I(net124));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__290__A2 (.I(_131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__291__B2 (.I(_136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__292__A1 (.I(_136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__293__A2 (.I(_071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__293__B1 (.I(_118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__293__B2 (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__295__A1 (.I(net124));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__295__A2 (.I(net79));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__295__A3 (.I(net80));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__295__A4 (.I(_131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__296__I (.I(net80));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__297__A1 (.I(_136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__299__B1 (.I(_118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__299__B2 (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__300__B (.I(net142));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__301__A1 (.I(net81));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__302__A1 (.I(net258));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__302__A2 (.I(_065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__302__C2 (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__303__A1 (.I(_043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__306__A1 (.I(_081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__308__I1 (.I(_084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__310__I1 (.I(net136));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__312__I1 (.I(net135));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__314__I1 (.I(net133));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__317__I1 (.I(net132));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__319__I1 (.I(net130));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__321__I1 (.I(net129));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__325__I1 (.I(net128));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__333__I (.I(net124));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__337__A1 (.I(_136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__340__I1 (.I(net81));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__342__CLK (.I(\clknet_2_0__leaf_counter.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__343__CLK (.I(\clknet_2_2__leaf_counter.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__344__CLK (.I(\clknet_2_2__leaf_counter.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__345__CLK (.I(\clknet_2_2__leaf_counter.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__346__CLK (.I(\clknet_2_2__leaf_counter.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__347__CLK (.I(\clknet_2_2__leaf_counter.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__348__CLK (.I(\clknet_2_2__leaf_counter.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__349__CLK (.I(\clknet_2_2__leaf_counter.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__350__CLK (.I(\clknet_2_2__leaf_counter.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__352__CLK (.I(\clknet_2_1__leaf_counter.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__357__CLK (.I(\clknet_2_2__leaf_counter.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__359__CLK (.I(\clknet_2_0__leaf_counter.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__360__CLK (.I(\clknet_2_0__leaf_counter.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__361__CLK (.I(\clknet_2_0__leaf_counter.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__362__CLK (.I(\clknet_2_0__leaf_counter.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__363__CLK (.I(\clknet_2_0__leaf_counter.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__364__CLK (.I(\clknet_2_1__leaf_counter.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__365__CLK (.I(\clknet_2_0__leaf_counter.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__366__CLK (.I(\clknet_2_1__leaf_counter.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__367__CLK (.I(\clknet_2_0__leaf_counter.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__368__CLK (.I(\clknet_2_0__leaf_counter.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__369__CLK (.I(\clknet_2_1__leaf_counter.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__370__CLK (.I(\clknet_2_1__leaf_counter.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__371__CLK (.I(\clknet_2_1__leaf_counter.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__372__CLK (.I(\clknet_2_1__leaf_counter.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__373__CLK (.I(\clknet_2_1__leaf_counter.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__374__CLK (.I(\clknet_2_0__leaf_counter.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__442__I (.I(net142));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__443__I (.I(net142));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__444__I (.I(net142));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__445__I (.I(net143));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__446__I (.I(net143));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__447__I (.I(net143));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__450__I (.I(net140));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__451__I (.I(net140));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__454__I (.I(net138));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__455__I (.I(net138));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__456__I (.I(net138));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__457__I (.I(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__458__I (.I(net82));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__459__I (.I(net136));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__460__I (.I(net135));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__461__I (.I(net133));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__462__I (.I(net132));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__463__I (.I(net130));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__464__I (.I(net129));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__465__I (.I(net89));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__466__I (.I(net128));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__468__I (.I(net77));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__470__I (.I(net79));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__471__I (.I(net80));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__472__I (.I(net81));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_clkbuf_0_counter.clk_I  (.I(\counter.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_clkbuf_2_0__f_counter.clk_I  (.I(\clknet_0_counter.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_clkbuf_2_1__f_counter.clk_I  (.I(\clknet_0_counter.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_clkbuf_2_2__f_counter.clk_I  (.I(\clknet_0_counter.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_clkbuf_2_3__f_counter.clk_I  (.I(\clknet_0_counter.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout125_I (.I(net126));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout127_I (.I(net76));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout128_I (.I(net90));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout129_I (.I(net88));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout130_I (.I(net131));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout132_I (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout135_I (.I(net84));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout138_I (.I(net140));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout139_I (.I(net140));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout140_I (.I(net145));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout141_I (.I(net145));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout142_I (.I(net143));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout143_I (.I(net145));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout144_I (.I(net145));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold13_I (.I(la_data_in[47]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold17_I (.I(la_data_in[60]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold1_I (.I(la_data_in[53]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold21_I (.I(la_data_in[48]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold25_I (.I(la_data_in[46]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold29_I (.I(la_data_in[59]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold30_I (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold33_I (.I(la_data_in[50]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold37_I (.I(la_data_in[49]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold41_I (.I(la_data_in[55]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold42_I (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold45_I (.I(la_data_in[61]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold46_I (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold49_I (.I(la_data_in[54]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold50_I (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold53_I (.I(la_data_in[57]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold54_I (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold57_I (.I(la_data_in[56]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold58_I (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold5_I (.I(la_data_in[51]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold61_I (.I(la_data_in[58]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold62_I (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold65_I (.I(la_data_in[63]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold66_I (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold68_I (.I(la_oenb[60]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold71_I (.I(la_oenb[47]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold75_I (.I(la_oenb[52]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold76_I (.I(la_oenb[59]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold78_I (.I(la_oenb[48]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold79_I (.I(la_oenb[55]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold81_I (.I(la_oenb[51]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold82_I (.I(la_oenb[53]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold83_I (.I(la_oenb[46]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold84_I (.I(la_oenb[49]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold85_I (.I(la_oenb[56]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold86_I (.I(la_oenb[61]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold87_I (.I(la_oenb[50]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold88_I (.I(la_oenb[58]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold89_I (.I(la_oenb[57]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold90_I (.I(la_oenb[54]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold91_I (.I(la_oenb[63]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold9_I (.I(la_data_in[52]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input17_I (.I(la_data_in[62]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input35_I (.I(la_oenb[62]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input37_I (.I(wb_rst_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input38_I (.I(wbs_cyc_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input39_I (.I(wbs_dat_i[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input40_I (.I(wbs_dat_i[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input41_I (.I(wbs_dat_i[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input42_I (.I(wbs_dat_i[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input43_I (.I(wbs_dat_i[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input44_I (.I(wbs_dat_i[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input45_I (.I(wbs_dat_i[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input46_I (.I(wbs_dat_i[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input47_I (.I(wbs_dat_i[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input48_I (.I(wbs_dat_i[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input49_I (.I(wbs_dat_i[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input50_I (.I(wbs_dat_i[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input51_I (.I(wbs_dat_i[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input52_I (.I(wbs_dat_i[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input53_I (.I(wbs_dat_i[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input54_I (.I(wbs_dat_i[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input55_I (.I(wbs_sel_i[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input56_I (.I(wbs_sel_i[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input57_I (.I(wbs_stb_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input58_I (.I(wbs_we_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output107_I (.I(net107));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output65_I (.I(net138));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output75_I (.I(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output76_I (.I(net76));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output77_I (.I(net77));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output78_I (.I(net126));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output79_I (.I(net79));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output80_I (.I(net80));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output81_I (.I(net81));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output82_I (.I(net82));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output83_I (.I(net137));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output84_I (.I(net84));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output85_I (.I(net134));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output86_I (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output87_I (.I(net131));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output88_I (.I(net88));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output89_I (.I(net89));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output90_I (.I(net90));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_100_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_100_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_100_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_100_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_100_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_100_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_100_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_100_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_100_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_100_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_100_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_100_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_100_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_101_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_101_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_101_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_101_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_101_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_101_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_101_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_101_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_101_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_101_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_101_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_101_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_102_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_102_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_102_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_102_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_102_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_102_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_102_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_102_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_102_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_102_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_102_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_102_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_102_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_103_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_103_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_103_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_103_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_103_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_103_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_103_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_103_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_103_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_103_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_103_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_103_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_104_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_104_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_104_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_104_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_104_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_104_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_104_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_104_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_104_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_104_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_104_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_104_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_104_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_105_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_105_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_105_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_105_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_105_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_105_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_105_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_105_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_105_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_105_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_105_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_105_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_106_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_106_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_106_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_106_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_106_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_106_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_106_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_106_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_106_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_106_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_106_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_106_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_106_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_107_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_107_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_107_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_107_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_107_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_107_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_107_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_107_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_107_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_107_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_107_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_107_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_108_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_108_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_108_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_108_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_108_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_108_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_108_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_108_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_108_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_108_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_108_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_108_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_109_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_109_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_109_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_109_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_109_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_109_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_109_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_109_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_109_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_109_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_109_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_109_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_110_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_110_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_110_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_110_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_110_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_110_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_110_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_110_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_110_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_110_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_110_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_110_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_110_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_111_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_111_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_111_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_111_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_111_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_111_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_111_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_111_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_111_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_111_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_111_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_111_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_112_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_112_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_112_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_112_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_112_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_112_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_112_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_112_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_112_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_112_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_112_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_112_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_112_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_113_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_113_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_113_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_113_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_113_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_113_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_113_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_113_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_113_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_113_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_113_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_113_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_114_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_114_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_114_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_114_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_114_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_114_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_114_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_114_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_114_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_114_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_114_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_115_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_115_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_115_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_115_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_115_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_115_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_115_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_115_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_115_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_115_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_115_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_115_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_116_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_116_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_116_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_116_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_116_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_116_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_116_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_116_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_116_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_116_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_116_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_116_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_116_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_117_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_117_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_117_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_117_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_117_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_117_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_117_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_117_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_117_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_117_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_117_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_117_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_118_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_118_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_118_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_118_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_118_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_118_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_118_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_118_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_118_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_118_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_118_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_118_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_118_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_118_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_118_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_118_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_118_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_118_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_118_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_118_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_118_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_118_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_118_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_118_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_13_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_13_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_14_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_14_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_15_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_15_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_16_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_18_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_21_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_24_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_26_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_28_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_30_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_31_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_32_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_3_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_3_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_47_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_48_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_48_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_50_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_50_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_56_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_56_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_58_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_58_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_5_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_5_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_60_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_60_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_62_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_63_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_64_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_64_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_66_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_66_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_67_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_67_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_67_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_67_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_67_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_67_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_67_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_67_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_67_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_67_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_67_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_67_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_68_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_68_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_68_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_68_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_68_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_68_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_68_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_68_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_68_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_68_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_68_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_69_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_69_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_69_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_69_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_69_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_69_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_69_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_69_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_69_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_69_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_69_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_69_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_70_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_70_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_70_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_70_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_70_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_70_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_70_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_70_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_70_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_70_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_70_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_70_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_70_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_71_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_71_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_71_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_71_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_71_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_71_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_71_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_71_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_71_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_71_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_71_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_71_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_72_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_72_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_72_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_72_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_72_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_72_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_72_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_72_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_72_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_72_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_72_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_73_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_73_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_73_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_73_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_73_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_73_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_73_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_73_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_73_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_73_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_73_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_73_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_74_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_74_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_74_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_74_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_74_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_74_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_74_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_74_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_74_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_74_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_74_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_74_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_74_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_75_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_75_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_75_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_75_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_75_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_75_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_75_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_75_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_75_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_75_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_75_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_75_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_76_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_76_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_76_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_76_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_76_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_76_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_76_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_76_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_76_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_76_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_76_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_76_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_76_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_77_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_77_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_77_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_77_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_77_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_77_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_77_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_77_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_77_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_77_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_77_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_78_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_78_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_78_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_78_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_78_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_78_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_78_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_78_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_78_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_78_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_78_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_78_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_79_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_79_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_79_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_79_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_79_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_79_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_79_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_79_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_79_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_79_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_79_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_79_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_80_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_80_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_80_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_80_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_80_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_80_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_80_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_80_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_80_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_80_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_80_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_81_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_81_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_81_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_81_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_81_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_81_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_81_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_81_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_81_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_81_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_81_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_81_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_82_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_82_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_82_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_82_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_82_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_82_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_82_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_82_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_82_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_82_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_82_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_82_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_83_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_83_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_83_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_83_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_83_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_83_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_83_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_83_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_83_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_83_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_83_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_83_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_84_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_84_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_84_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_84_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_84_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_84_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_84_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_84_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_84_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_84_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_84_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_84_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_84_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_85_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_85_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_85_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_85_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_85_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_85_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_85_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_85_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_85_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_85_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_85_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_85_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_86_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_86_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_86_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_86_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_86_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_86_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_86_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_86_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_86_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_86_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_86_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_86_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_86_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_87_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_87_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_87_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_87_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_87_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_87_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_87_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_87_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_87_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_87_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_87_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_87_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_88_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_88_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_88_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_88_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_88_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_88_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_88_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_88_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_88_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_88_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_88_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_88_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_88_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_89_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_89_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_89_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_89_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_89_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_89_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_89_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_89_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_89_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_89_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_89_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_89_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_90_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_90_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_90_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_90_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_90_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_90_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_90_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_90_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_90_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_90_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_90_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_90_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_90_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_91_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_91_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_91_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_91_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_91_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_91_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_91_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_91_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_91_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_91_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_91_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_91_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_92_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_92_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_92_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_92_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_92_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_92_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_92_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_92_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_92_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_92_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_92_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_92_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_93_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_93_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_93_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_93_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_93_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_93_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_93_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_93_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_93_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_93_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_93_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_93_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_94_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_94_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_94_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_94_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_94_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_94_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_94_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_94_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_94_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_94_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_94_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_94_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_94_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_95_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_95_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_95_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_95_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_95_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_95_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_95_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_95_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_95_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_95_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_95_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_95_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_96_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_96_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_96_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_96_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_96_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_96_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_96_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_96_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_96_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_96_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_96_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_96_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_96_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_97_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_97_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_97_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_97_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_97_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_97_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_97_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_97_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_97_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_97_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_97_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_97_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_98_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_98_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_98_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_98_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_98_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_98_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_98_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_98_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_98_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_98_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_98_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_99_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_99_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_99_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_99_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_99_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_99_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_99_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_99_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_99_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_99_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_99_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_99_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_858 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Left_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_100_Left_219 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_100_Right_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_101_Left_220 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_101_Right_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_102_Left_221 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_102_Right_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_103_Left_222 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_103_Right_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_104_Left_223 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_104_Right_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_105_Left_224 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_105_Right_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_106_Left_225 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_106_Right_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_107_Left_226 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_107_Right_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_108_Left_227 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_108_Right_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_109_Left_228 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_109_Right_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Left_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_110_Left_229 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_110_Right_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_111_Left_230 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_111_Right_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_112_Left_231 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_112_Right_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_113_Left_232 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_113_Right_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_114_Left_233 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_114_Right_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_115_Left_234 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_115_Right_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_116_Left_235 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_116_Right_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_117_Left_236 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_117_Right_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_118_Left_237 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_118_Right_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Left_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Left_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Left_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Left_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Left_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Left_135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Left_136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Left_137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Left_138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Left_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Left_139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Left_140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Left_141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Left_142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Left_143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Left_144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Left_145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Right_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Left_146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Right_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Left_147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Right_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Left_148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Right_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Left_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Left_149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Right_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Left_150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Right_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Left_151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Right_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Left_152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Right_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Left_153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Right_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Left_154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Right_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Left_155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Right_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Left_156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Right_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Left_157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Right_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Left_158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Right_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Left_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Left_159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Right_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Left_160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Right_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Left_161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Right_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Left_162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Right_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Left_163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Right_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Left_164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Right_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Left_165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Right_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_Left_166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_Right_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_Left_167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_Right_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_Left_168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_Right_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Left_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_Left_169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_Right_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_Left_170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_Right_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_Left_171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_Right_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_Left_172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_Right_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_Left_173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_Right_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_Left_174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_Right_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_Left_175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_Right_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_Left_176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_Right_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_Left_177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_Right_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_Left_178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_Right_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Left_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_Left_179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_Right_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_Left_180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_Right_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_Left_181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_Right_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_Left_182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_Right_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_Left_183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_Right_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_Left_184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_Right_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_Left_185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_Right_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_Left_186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_Right_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_Left_187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_Right_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_Left_188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_Right_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Left_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_Left_189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_Right_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_Left_190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_Right_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_Left_191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_Right_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_Left_192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_Right_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_Left_193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_Right_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_Left_194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_Right_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_Left_195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_Right_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_Left_196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_Right_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_Left_197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_Right_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_Left_198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_Right_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Left_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_Left_199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_Right_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_Left_200 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_Right_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_Left_201 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_Right_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_83_Left_202 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_83_Right_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_84_Left_203 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_84_Right_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_85_Left_204 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_85_Right_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_86_Left_205 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_86_Right_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_87_Left_206 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_87_Right_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_88_Left_207 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_88_Right_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_89_Left_208 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_89_Right_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Left_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_90_Left_209 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_90_Right_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_91_Left_210 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_91_Right_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_92_Left_211 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_92_Right_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_93_Left_212 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_93_Right_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_94_Left_213 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_94_Right_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_95_Left_214 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_95_Right_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_96_Left_215 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_96_Right_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_97_Left_216 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_97_Right_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_98_Left_217 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_98_Right_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_99_Left_218 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_99_Right_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Left_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_370 ();
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _170_ (.I0(net278),
    .I1(net37),
    .S(net36),
    .Z(_033_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _171_ (.I(_033_),
    .Z(net65));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _172_ (.I0(net17),
    .I1(wb_clk_i),
    .S(net35),
    .Z(_034_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _173_ (.I(_034_),
    .Z(\counter.clk ));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _174_ (.I(net57),
    .Z(_035_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _175_ (.I(_035_),
    .Z(_036_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _176_ (.I(net38),
    .Z(_037_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _177_ (.I(_037_),
    .Z(_038_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _178_ (.A1(_036_),
    .A2(_038_),
    .ZN(_039_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _179_ (.A1(net107),
    .A2(_039_),
    .Z(_040_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _180_ (.A1(net279),
    .A2(_040_),
    .ZN(_041_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _181_ (.I(_041_),
    .Z(_042_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _182_ (.I(_042_),
    .Z(_000_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _183_ (.I(net279),
    .Z(_043_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _184_ (.I(_043_),
    .Z(_044_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _185_ (.A1(_036_),
    .A2(_038_),
    .B(net19),
    .ZN(_045_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _186_ (.A1(net107),
    .A2(_039_),
    .ZN(_046_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _187_ (.A1(net58),
    .A2(net55),
    .Z(_047_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _188_ (.A1(_046_),
    .A2(_047_),
    .Z(_048_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _189_ (.I(_048_),
    .Z(_049_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _190_ (.I(_035_),
    .Z(_050_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _191_ (.I(_037_),
    .Z(_051_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _192_ (.A1(_050_),
    .A2(_051_),
    .B(net25),
    .ZN(_052_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _193_ (.A1(_050_),
    .A2(_051_),
    .B(net20),
    .ZN(_053_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _194_ (.A1(_052_),
    .A2(_053_),
    .ZN(_054_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _195_ (.A1(_050_),
    .A2(_051_),
    .B(net23),
    .ZN(_055_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _196_ (.A1(_050_),
    .A2(_051_),
    .B(net24),
    .ZN(_056_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _197_ (.A1(_055_),
    .A2(_056_),
    .ZN(_057_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _198_ (.I(net57),
    .Z(_058_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _199_ (.I(net38),
    .Z(_059_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _200_ (.A1(_058_),
    .A2(_059_),
    .B(net22),
    .ZN(_060_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _201_ (.A1(_035_),
    .A2(_037_),
    .B(net21),
    .ZN(_061_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _202_ (.A1(_058_),
    .A2(_059_),
    .B(net33),
    .ZN(_062_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _203_ (.I(_035_),
    .Z(_063_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _204_ (.I(_037_),
    .Z(_064_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _205_ (.A1(_063_),
    .A2(_064_),
    .B(net34),
    .ZN(_065_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _206_ (.A1(_060_),
    .A2(_061_),
    .A3(_062_),
    .A4(_065_),
    .ZN(_066_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _207_ (.A1(_063_),
    .A2(_064_),
    .B(net30),
    .ZN(_067_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _208_ (.A1(_058_),
    .A2(_059_),
    .B(net27),
    .ZN(_068_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _209_ (.A1(_058_),
    .A2(_059_),
    .B(net28),
    .ZN(_069_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _210_ (.A1(_067_),
    .A2(_068_),
    .A3(_069_),
    .A4(_045_),
    .ZN(_070_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _211_ (.A1(_063_),
    .A2(_038_),
    .B(net32),
    .ZN(_071_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _212_ (.A1(_063_),
    .A2(_064_),
    .B(net26),
    .ZN(_072_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _213_ (.A1(_036_),
    .A2(_064_),
    .B(net31),
    .ZN(_073_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _214_ (.A1(_036_),
    .A2(_038_),
    .B(net29),
    .ZN(_074_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _215_ (.A1(_071_),
    .A2(_072_),
    .A3(_073_),
    .A4(_074_),
    .ZN(_075_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _216_ (.A1(_066_),
    .A2(_070_),
    .A3(_075_),
    .Z(_076_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _217_ (.A1(_040_),
    .A2(net284),
    .A3(_057_),
    .A4(_076_),
    .ZN(_077_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _218_ (.A1(_040_),
    .A2(_047_),
    .B(_077_),
    .ZN(_078_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _219_ (.I(_078_),
    .Z(_079_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _220_ (.I(net75),
    .Z(_080_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _221_ (.I(_080_),
    .ZN(_081_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _222_ (.A1(net238),
    .A2(_045_),
    .B1(_049_),
    .B2(net39),
    .C1(_079_),
    .C2(_081_),
    .ZN(_082_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _223_ (.A1(_044_),
    .A2(net239),
    .ZN(_001_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _224_ (.I(_078_),
    .Z(_083_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _225_ (.I(net82),
    .Z(_084_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _226_ (.A1(_080_),
    .A2(_084_),
    .Z(_085_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _227_ (.A1(net226),
    .A2(_053_),
    .B1(_083_),
    .B2(_085_),
    .C1(_049_),
    .C2(net46),
    .ZN(_086_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _228_ (.A1(_044_),
    .A2(net227),
    .ZN(_002_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _229_ (.A1(_080_),
    .A2(_084_),
    .ZN(_087_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _230_ (.A1(net136),
    .A2(_087_),
    .ZN(_088_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _231_ (.A1(net234),
    .A2(_061_),
    .B1(_083_),
    .B2(_088_),
    .C1(_049_),
    .C2(net47),
    .ZN(_089_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _232_ (.A1(_044_),
    .A2(net235),
    .ZN(_003_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _233_ (.A1(_080_),
    .A2(_084_),
    .A3(net136),
    .ZN(_090_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _234_ (.A1(net135),
    .A2(_090_),
    .ZN(_091_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _235_ (.A1(net250),
    .A2(_060_),
    .B1(_083_),
    .B2(_091_),
    .C1(_049_),
    .C2(net48),
    .ZN(_092_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _236_ (.A1(_044_),
    .A2(net251),
    .ZN(_004_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _237_ (.I(_043_),
    .Z(_093_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _238_ (.A1(net75),
    .A2(net82),
    .A3(net137),
    .A4(net135),
    .Z(_094_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _239_ (.A1(net133),
    .A2(_094_),
    .Z(_095_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _240_ (.I(_048_),
    .Z(_096_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _241_ (.A1(net246),
    .A2(_055_),
    .B1(_083_),
    .B2(_095_),
    .C1(_096_),
    .C2(net49),
    .ZN(_097_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _242_ (.A1(_093_),
    .A2(net247),
    .ZN(_005_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _243_ (.A1(net133),
    .A2(net132),
    .Z(_098_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _244_ (.A1(_094_),
    .A2(_098_),
    .Z(_099_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _245_ (.A1(net134),
    .A2(_094_),
    .B(net132),
    .ZN(_100_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _246_ (.A1(_099_),
    .A2(_100_),
    .ZN(_101_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _247_ (.A1(net218),
    .A2(_056_),
    .B1(_079_),
    .B2(_101_),
    .C1(_096_),
    .C2(net50),
    .ZN(_102_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _248_ (.A1(_093_),
    .A2(net219),
    .ZN(_006_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _249_ (.A1(net130),
    .A2(_099_),
    .Z(_103_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _250_ (.A1(net222),
    .A2(_052_),
    .B1(_079_),
    .B2(_103_),
    .C1(_096_),
    .C2(net51),
    .ZN(_104_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _251_ (.A1(_093_),
    .A2(net223),
    .ZN(_007_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _252_ (.A1(net130),
    .A2(_099_),
    .ZN(_105_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _253_ (.A1(net129),
    .A2(_105_),
    .ZN(_106_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _254_ (.A1(net214),
    .A2(_072_),
    .B1(_079_),
    .B2(_106_),
    .C1(_096_),
    .C2(net52),
    .ZN(_107_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _255_ (.A1(_093_),
    .A2(net215),
    .ZN(_008_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _256_ (.I(_043_),
    .Z(_108_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _257_ (.A1(net58),
    .A2(net56),
    .ZN(_109_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _258_ (.A1(_046_),
    .A2(_109_),
    .ZN(_110_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _259_ (.A1(net285),
    .A2(_110_),
    .ZN(_111_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _260_ (.I(_111_),
    .Z(_112_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _261_ (.I(net89),
    .ZN(_113_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _262_ (.A1(net131),
    .A2(net129),
    .A3(_094_),
    .A4(_098_),
    .ZN(_114_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _263_ (.I(_114_),
    .Z(_115_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _264_ (.A1(_113_),
    .A2(_115_),
    .Z(_116_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _265_ (.A1(_040_),
    .A2(_109_),
    .ZN(_117_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _266_ (.I(_117_),
    .Z(_118_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _267_ (.A1(net262),
    .A2(_068_),
    .B1(_112_),
    .B2(_116_),
    .C1(_118_),
    .C2(net53),
    .ZN(_119_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _268_ (.A1(_108_),
    .A2(net263),
    .ZN(_009_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _269_ (.A1(_113_),
    .A2(_115_),
    .ZN(_120_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _270_ (.A1(net89),
    .A2(net128),
    .ZN(_121_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _271_ (.A1(net128),
    .A2(_120_),
    .B1(_121_),
    .B2(_115_),
    .C(_111_),
    .ZN(_122_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _272_ (.A1(net254),
    .A2(_069_),
    .B1(_118_),
    .B2(net54),
    .ZN(_123_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _273_ (.A1(_122_),
    .A2(net255),
    .B(net139),
    .ZN(_010_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _274_ (.A1(_115_),
    .A2(_121_),
    .ZN(_124_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _275_ (.A1(net127),
    .A2(_124_),
    .Z(_125_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _276_ (.I(_117_),
    .Z(_126_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _277_ (.A1(net270),
    .A2(_074_),
    .B1(_112_),
    .B2(_125_),
    .C1(_126_),
    .C2(net40),
    .ZN(_127_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _278_ (.A1(_108_),
    .A2(net271),
    .ZN(_011_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _279_ (.A1(net127),
    .A2(_124_),
    .B(net77),
    .ZN(_128_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _280_ (.I(net127),
    .ZN(_129_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _281_ (.I(net77),
    .ZN(_130_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _282_ (.A1(_129_),
    .A2(_130_),
    .A3(_114_),
    .A4(_121_),
    .ZN(_131_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _283_ (.A1(_128_),
    .A2(_131_),
    .ZN(_132_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _284_ (.A1(net266),
    .A2(_067_),
    .B1(_112_),
    .B2(_132_),
    .C1(_126_),
    .C2(net41),
    .ZN(_133_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _285_ (.A1(_108_),
    .A2(net267),
    .ZN(_012_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _286_ (.A1(net124),
    .A2(_131_),
    .Z(_134_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _287_ (.A1(net274),
    .A2(_073_),
    .B1(_111_),
    .B2(_134_),
    .C1(_126_),
    .C2(net42),
    .ZN(_135_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _288_ (.A1(_108_),
    .A2(net275),
    .ZN(_013_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _289_ (.I(net79),
    .ZN(_136_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _290_ (.A1(net124),
    .A2(_131_),
    .ZN(_137_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _291_ (.A1(net285),
    .A2(_110_),
    .B1(_137_),
    .B2(_136_),
    .ZN(_138_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _292_ (.A1(_136_),
    .A2(_137_),
    .B(_138_),
    .ZN(_139_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _293_ (.A1(net242),
    .A2(_071_),
    .B1(_118_),
    .B2(net43),
    .ZN(_140_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _294_ (.A1(_139_),
    .A2(net243),
    .B(net139),
    .ZN(_014_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _295_ (.A1(net124),
    .A2(net79),
    .A3(net80),
    .A4(_131_),
    .ZN(_141_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _296_ (.I(net80),
    .ZN(_142_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _297_ (.A1(_136_),
    .A2(_137_),
    .B(_142_),
    .ZN(_143_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _298_ (.A1(_112_),
    .A2(_141_),
    .A3(_143_),
    .ZN(_144_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _299_ (.A1(net230),
    .A2(_062_),
    .B1(_118_),
    .B2(net44),
    .ZN(_145_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _300_ (.A1(_144_),
    .A2(net231),
    .B(net142),
    .ZN(_015_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _301_ (.A1(net81),
    .A2(_141_),
    .ZN(_146_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _302_ (.A1(net258),
    .A2(_065_),
    .B1(_111_),
    .B2(_146_),
    .C1(_126_),
    .C2(net45),
    .ZN(_147_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _303_ (.A1(_043_),
    .A2(net259),
    .ZN(_016_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _304_ (.I(_041_),
    .Z(_148_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _305_ (.A1(net108),
    .A2(_148_),
    .ZN(_149_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _306_ (.A1(_081_),
    .A2(_000_),
    .B(_149_),
    .ZN(_017_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _307_ (.I(_042_),
    .Z(_150_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _308_ (.I0(net115),
    .I1(_084_),
    .S(_150_),
    .Z(_151_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _309_ (.I(_151_),
    .Z(_018_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _310_ (.I0(net116),
    .I1(net136),
    .S(_150_),
    .Z(_152_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _311_ (.I(_152_),
    .Z(_019_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _312_ (.I0(net117),
    .I1(net135),
    .S(_150_),
    .Z(_153_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _313_ (.I(_153_),
    .Z(_020_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _314_ (.I0(net118),
    .I1(net133),
    .S(_150_),
    .Z(_154_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _315_ (.I(_154_),
    .Z(_021_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _316_ (.I(_042_),
    .Z(_155_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _317_ (.I0(net119),
    .I1(net132),
    .S(_155_),
    .Z(_156_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _318_ (.I(_156_),
    .Z(_022_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _319_ (.I0(net120),
    .I1(net130),
    .S(_155_),
    .Z(_157_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _320_ (.I(_157_),
    .Z(_023_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _321_ (.I0(net121),
    .I1(net129),
    .S(_155_),
    .Z(_158_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _322_ (.I(_158_),
    .Z(_024_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _323_ (.A1(net122),
    .A2(_148_),
    .ZN(_159_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _324_ (.A1(_113_),
    .A2(_000_),
    .B(_159_),
    .ZN(_025_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _325_ (.I0(net123),
    .I1(net128),
    .S(_155_),
    .Z(_160_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _326_ (.I(_160_),
    .Z(_026_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _327_ (.A1(net109),
    .A2(_148_),
    .ZN(_161_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _328_ (.A1(_129_),
    .A2(_000_),
    .B(_161_),
    .ZN(_027_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _329_ (.I(_041_),
    .Z(_162_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _330_ (.I(_162_),
    .Z(_163_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _331_ (.A1(net110),
    .A2(_148_),
    .ZN(_164_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _332_ (.A1(_130_),
    .A2(_163_),
    .B(_164_),
    .ZN(_028_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _333_ (.I(net124),
    .ZN(_165_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _334_ (.A1(net111),
    .A2(net281),
    .ZN(_166_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _335_ (.A1(_165_),
    .A2(_163_),
    .B(_166_),
    .ZN(_029_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _336_ (.A1(net112),
    .A2(net281),
    .ZN(_167_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _337_ (.A1(_136_),
    .A2(_163_),
    .B(_167_),
    .ZN(_030_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _338_ (.A1(net113),
    .A2(net281),
    .ZN(_168_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _339_ (.A1(_142_),
    .A2(_163_),
    .B(_168_),
    .ZN(_031_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _340_ (.I0(net114),
    .I1(net81),
    .S(_042_),
    .Z(_169_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _341_ (.I(_169_),
    .Z(_032_));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _342_ (.D(_000_),
    .CLK(\clknet_2_0__leaf_counter.clk ),
    .Q(net107));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _343_ (.D(net240),
    .CLK(\clknet_2_2__leaf_counter.clk ),
    .Q(net75));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _344_ (.D(net228),
    .CLK(\clknet_2_2__leaf_counter.clk ),
    .Q(net82));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _345_ (.D(net236),
    .CLK(\clknet_2_2__leaf_counter.clk ),
    .Q(net83));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _346_ (.D(net252),
    .CLK(\clknet_2_2__leaf_counter.clk ),
    .Q(net84));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _347_ (.D(net248),
    .CLK(\clknet_2_2__leaf_counter.clk ),
    .Q(net85));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _348_ (.D(net220),
    .CLK(\clknet_2_2__leaf_counter.clk ),
    .Q(net86));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _349_ (.D(net224),
    .CLK(\clknet_2_2__leaf_counter.clk ),
    .Q(net87));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _350_ (.D(net216),
    .CLK(\clknet_2_2__leaf_counter.clk ),
    .Q(net88));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _351_ (.D(net264),
    .CLK(\clknet_2_3__leaf_counter.clk ),
    .Q(net89));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _352_ (.D(net256),
    .CLK(\clknet_2_1__leaf_counter.clk ),
    .Q(net90));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _353_ (.D(net272),
    .CLK(\clknet_2_3__leaf_counter.clk ),
    .Q(net76));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _354_ (.D(net268),
    .CLK(\clknet_2_3__leaf_counter.clk ),
    .Q(net77));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _355_ (.D(net276),
    .CLK(\clknet_2_3__leaf_counter.clk ),
    .Q(net78));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _356_ (.D(net244),
    .CLK(\clknet_2_3__leaf_counter.clk ),
    .Q(net79));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _357_ (.D(net232),
    .CLK(\clknet_2_2__leaf_counter.clk ),
    .Q(net80));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _358_ (.D(net260),
    .CLK(\clknet_2_3__leaf_counter.clk ),
    .Q(net81));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _359_ (.D(_017_),
    .CLK(\clknet_2_0__leaf_counter.clk ),
    .Q(net108));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _360_ (.D(_018_),
    .CLK(\clknet_2_0__leaf_counter.clk ),
    .Q(net115));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _361_ (.D(_019_),
    .CLK(\clknet_2_0__leaf_counter.clk ),
    .Q(net116));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _362_ (.D(_020_),
    .CLK(\clknet_2_0__leaf_counter.clk ),
    .Q(net117));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _363_ (.D(_021_),
    .CLK(\clknet_2_0__leaf_counter.clk ),
    .Q(net118));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _364_ (.D(_022_),
    .CLK(\clknet_2_1__leaf_counter.clk ),
    .Q(net119));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _365_ (.D(_023_),
    .CLK(\clknet_2_0__leaf_counter.clk ),
    .Q(net120));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _366_ (.D(_024_),
    .CLK(\clknet_2_1__leaf_counter.clk ),
    .Q(net121));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _367_ (.D(_025_),
    .CLK(\clknet_2_0__leaf_counter.clk ),
    .Q(net122));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _368_ (.D(_026_),
    .CLK(\clknet_2_0__leaf_counter.clk ),
    .Q(net123));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _369_ (.D(_027_),
    .CLK(\clknet_2_1__leaf_counter.clk ),
    .Q(net109));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _370_ (.D(_028_),
    .CLK(\clknet_2_1__leaf_counter.clk ),
    .Q(net110));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _371_ (.D(_029_),
    .CLK(\clknet_2_1__leaf_counter.clk ),
    .Q(net111));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _372_ (.D(_030_),
    .CLK(\clknet_2_1__leaf_counter.clk ),
    .Q(net112));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _373_ (.D(_031_),
    .CLK(\clknet_2_1__leaf_counter.clk ),
    .Q(net113));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _374_ (.D(_032_),
    .CLK(\clknet_2_0__leaf_counter.clk ),
    .Q(net114));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _442_ (.I(net142),
    .Z(net59));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _443_ (.I(net142),
    .Z(net66));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _444_ (.I(net142),
    .Z(net67));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _445_ (.I(net143),
    .Z(net68));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _446_ (.I(net143),
    .Z(net69));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _447_ (.I(net143),
    .Z(net70));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _448_ (.I(net144),
    .Z(net71));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _449_ (.I(net144),
    .Z(net72));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _450_ (.I(net140),
    .Z(net73));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _451_ (.I(net140),
    .Z(net74));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _452_ (.I(net141),
    .Z(net60));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _453_ (.I(net141),
    .Z(net61));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _454_ (.I(net138),
    .Z(net62));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _455_ (.I(net138),
    .Z(net63));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _456_ (.I(net138),
    .Z(net64));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _457_ (.I(net75),
    .Z(net91));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _458_ (.I(net82),
    .Z(net98));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _459_ (.I(net136),
    .Z(net99));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _460_ (.I(net135),
    .Z(net100));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _461_ (.I(net133),
    .Z(net101));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _462_ (.I(net132),
    .Z(net102));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _463_ (.I(net130),
    .Z(net103));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _464_ (.I(net129),
    .Z(net104));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _465_ (.I(net89),
    .Z(net105));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _466_ (.I(net128),
    .Z(net106));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _467_ (.I(net127),
    .Z(net92));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _468_ (.I(net77),
    .Z(net93));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _469_ (.I(net125),
    .Z(net94));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _470_ (.I(net79),
    .Z(net95));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _471_ (.I(net80),
    .Z(net96));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _472_ (.I(net81),
    .Z(net97));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \clkbuf_0_counter.clk  (.I(\counter.clk ),
    .Z(\clknet_0_counter.clk ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \clkbuf_2_0__f_counter.clk  (.I(\clknet_0_counter.clk ),
    .Z(\clknet_2_0__leaf_counter.clk ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \clkbuf_2_1__f_counter.clk  (.I(\clknet_0_counter.clk ),
    .Z(\clknet_2_1__leaf_counter.clk ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \clkbuf_2_2__f_counter.clk  (.I(\clknet_0_counter.clk ),
    .Z(\clknet_2_2__leaf_counter.clk ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \clkbuf_2_3__f_counter.clk  (.I(\clknet_0_counter.clk ),
    .Z(\clknet_2_3__leaf_counter.clk ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 fanout124 (.I(net125),
    .Z(net124));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout125 (.I(net126),
    .Z(net125));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 fanout126 (.I(net78),
    .Z(net126));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout127 (.I(net76),
    .Z(net127));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 fanout128 (.I(net90),
    .Z(net128));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 fanout129 (.I(net88),
    .Z(net129));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 fanout130 (.I(net131),
    .Z(net130));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 fanout131 (.I(net87),
    .Z(net131));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 fanout132 (.I(net86),
    .Z(net132));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 fanout133 (.I(net85),
    .Z(net133));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 fanout134 (.I(net85),
    .Z(net134));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 fanout135 (.I(net84),
    .Z(net135));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 fanout136 (.I(net83),
    .Z(net136));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 fanout137 (.I(net83),
    .Z(net137));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 fanout138 (.I(net140),
    .Z(net138));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout139 (.I(net140),
    .Z(net139));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 fanout140 (.I(net145),
    .Z(net140));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout141 (.I(net145),
    .Z(net141));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 fanout142 (.I(net143),
    .Z(net142));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 fanout143 (.I(net145),
    .Z(net143));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout144 (.I(net145),
    .Z(net144));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 fanout145 (.I(net65),
    .Z(net145));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold1 (.I(la_data_in[53]),
    .Z(net213));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold10 (.I(net7),
    .Z(net222));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold11 (.I(_104_),
    .Z(net223));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold12 (.I(_007_),
    .Z(net224));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold13 (.I(la_data_in[47]),
    .Z(net225));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold14 (.I(net2),
    .Z(net226));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold15 (.I(_086_),
    .Z(net227));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold16 (.I(_002_),
    .Z(net228));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold17 (.I(la_data_in[60]),
    .Z(net229));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold18 (.I(net15),
    .Z(net230));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold19 (.I(_145_),
    .Z(net231));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold2 (.I(net8),
    .Z(net214));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold20 (.I(net286),
    .Z(net232));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold21 (.I(la_data_in[48]),
    .Z(net233));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold22 (.I(net3),
    .Z(net234));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold23 (.I(_089_),
    .Z(net235));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold24 (.I(_003_),
    .Z(net236));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold25 (.I(la_data_in[46]),
    .Z(net237));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold26 (.I(net1),
    .Z(net238));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold27 (.I(_082_),
    .Z(net239));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold28 (.I(_001_),
    .Z(net240));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold29 (.I(la_data_in[59]),
    .Z(net241));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold3 (.I(_107_),
    .Z(net215));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold30 (.I(net14),
    .Z(net242));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold31 (.I(_140_),
    .Z(net243));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold32 (.I(net289),
    .Z(net244));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold33 (.I(la_data_in[50]),
    .Z(net245));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold34 (.I(net5),
    .Z(net246));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold35 (.I(_097_),
    .Z(net247));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold36 (.I(_005_),
    .Z(net248));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold37 (.I(la_data_in[49]),
    .Z(net249));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold38 (.I(net4),
    .Z(net250));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold39 (.I(_092_),
    .Z(net251));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold4 (.I(_008_),
    .Z(net216));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold40 (.I(_004_),
    .Z(net252));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold41 (.I(la_data_in[55]),
    .Z(net253));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold42 (.I(net10),
    .Z(net254));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold43 (.I(_123_),
    .Z(net255));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold44 (.I(net292),
    .Z(net256));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold45 (.I(la_data_in[61]),
    .Z(net257));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold46 (.I(net16),
    .Z(net258));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold47 (.I(_147_),
    .Z(net259));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold48 (.I(_016_),
    .Z(net260));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold49 (.I(la_data_in[54]),
    .Z(net261));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold5 (.I(la_data_in[51]),
    .Z(net217));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold50 (.I(net9),
    .Z(net262));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold51 (.I(_119_),
    .Z(net263));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold52 (.I(_009_),
    .Z(net264));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold53 (.I(la_data_in[57]),
    .Z(net265));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold54 (.I(net12),
    .Z(net266));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold55 (.I(_133_),
    .Z(net267));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold56 (.I(_012_),
    .Z(net268));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold57 (.I(la_data_in[56]),
    .Z(net269));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold58 (.I(net11),
    .Z(net270));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold59 (.I(_127_),
    .Z(net271));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold6 (.I(net6),
    .Z(net218));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold60 (.I(_011_),
    .Z(net272));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold61 (.I(la_data_in[58]),
    .Z(net273));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 hold62 (.I(net13),
    .Z(net274));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold63 (.I(_135_),
    .Z(net275));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold64 (.I(_013_),
    .Z(net276));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold65 (.I(la_data_in[63]),
    .Z(net277));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold66 (.I(net18),
    .Z(net278));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold67 (.I(_033_),
    .Z(net279));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold68 (.I(la_oenb[60]),
    .Z(net280));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold69 (.I(_162_),
    .Z(net281));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold7 (.I(_102_),
    .Z(net219));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold70 (.I(net303),
    .Z(net282));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold71 (.I(la_oenb[47]),
    .Z(net283));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold72 (.I(_054_),
    .Z(net284));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 hold73 (.I(_077_),
    .Z(net285));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold74 (.I(_015_),
    .Z(net286));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold75 (.I(la_oenb[52]),
    .Z(net287));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold76 (.I(la_oenb[59]),
    .Z(net288));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold77 (.I(_014_),
    .Z(net289));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold78 (.I(la_oenb[48]),
    .Z(net290));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold79 (.I(la_oenb[55]),
    .Z(net291));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold8 (.I(_006_),
    .Z(net220));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold80 (.I(_010_),
    .Z(net292));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold81 (.I(la_oenb[51]),
    .Z(net293));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold82 (.I(la_oenb[53]),
    .Z(net294));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold83 (.I(la_oenb[46]),
    .Z(net295));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold84 (.I(la_oenb[49]),
    .Z(net296));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold85 (.I(la_oenb[56]),
    .Z(net297));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold86 (.I(la_oenb[61]),
    .Z(net298));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold87 (.I(la_oenb[50]),
    .Z(net299));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold88 (.I(la_oenb[58]),
    .Z(net300));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold89 (.I(la_oenb[57]),
    .Z(net301));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold9 (.I(la_data_in[52]),
    .Z(net221));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold90 (.I(la_oenb[54]),
    .Z(net302));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold91 (.I(la_oenb[63]),
    .Z(net303));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1 (.I(net237),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input10 (.I(net253),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input11 (.I(net269),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input12 (.I(net265),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input13 (.I(net273),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input14 (.I(net241),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input15 (.I(net229),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input16 (.I(net257),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input17 (.I(la_data_in[62]),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input18 (.I(net277),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input19 (.I(net295),
    .Z(net19));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input2 (.I(net225),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input20 (.I(net283),
    .Z(net20));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input21 (.I(net290),
    .Z(net21));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input22 (.I(net296),
    .Z(net22));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input23 (.I(net299),
    .Z(net23));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input24 (.I(net293),
    .Z(net24));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input25 (.I(net287),
    .Z(net25));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input26 (.I(net294),
    .Z(net26));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input27 (.I(net302),
    .Z(net27));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input28 (.I(net291),
    .Z(net28));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input29 (.I(net297),
    .Z(net29));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input3 (.I(net233),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input30 (.I(net301),
    .Z(net30));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input31 (.I(net300),
    .Z(net31));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input32 (.I(net288),
    .Z(net32));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input33 (.I(net280),
    .Z(net33));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input34 (.I(net298),
    .Z(net34));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input35 (.I(la_oenb[62]),
    .Z(net35));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input36 (.I(net282),
    .Z(net36));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input37 (.I(wb_rst_i),
    .Z(net37));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input38 (.I(wbs_cyc_i),
    .Z(net38));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input39 (.I(wbs_dat_i[0]),
    .Z(net39));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input4 (.I(net249),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input40 (.I(wbs_dat_i[10]),
    .Z(net40));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input41 (.I(wbs_dat_i[11]),
    .Z(net41));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input42 (.I(wbs_dat_i[12]),
    .Z(net42));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input43 (.I(wbs_dat_i[13]),
    .Z(net43));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input44 (.I(wbs_dat_i[14]),
    .Z(net44));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input45 (.I(wbs_dat_i[15]),
    .Z(net45));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input46 (.I(wbs_dat_i[1]),
    .Z(net46));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input47 (.I(wbs_dat_i[2]),
    .Z(net47));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input48 (.I(wbs_dat_i[3]),
    .Z(net48));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input49 (.I(wbs_dat_i[4]),
    .Z(net49));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input5 (.I(net245),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input50 (.I(wbs_dat_i[5]),
    .Z(net50));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input51 (.I(wbs_dat_i[6]),
    .Z(net51));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input52 (.I(wbs_dat_i[7]),
    .Z(net52));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input53 (.I(wbs_dat_i[8]),
    .Z(net53));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input54 (.I(wbs_dat_i[9]),
    .Z(net54));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input55 (.I(wbs_sel_i[0]),
    .Z(net55));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input56 (.I(wbs_sel_i[1]),
    .Z(net56));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input57 (.I(wbs_stb_i),
    .Z(net57));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input58 (.I(wbs_we_i),
    .Z(net58));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input6 (.I(net217),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input7 (.I(net221),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input8 (.I(net213),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input9 (.I(net261),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output100 (.I(net100),
    .Z(la_data_out[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output101 (.I(net101),
    .Z(la_data_out[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output102 (.I(net102),
    .Z(la_data_out[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output103 (.I(net103),
    .Z(la_data_out[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output104 (.I(net104),
    .Z(la_data_out[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output105 (.I(net105),
    .Z(la_data_out[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output106 (.I(net106),
    .Z(la_data_out[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output107 (.I(net107),
    .Z(wbs_ack_o));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output108 (.I(net108),
    .Z(wbs_dat_o[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output109 (.I(net109),
    .Z(wbs_dat_o[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output110 (.I(net110),
    .Z(wbs_dat_o[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output111 (.I(net111),
    .Z(wbs_dat_o[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output112 (.I(net112),
    .Z(wbs_dat_o[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output113 (.I(net113),
    .Z(wbs_dat_o[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output114 (.I(net114),
    .Z(wbs_dat_o[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output115 (.I(net115),
    .Z(wbs_dat_o[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output116 (.I(net116),
    .Z(wbs_dat_o[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output117 (.I(net117),
    .Z(wbs_dat_o[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output118 (.I(net118),
    .Z(wbs_dat_o[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output119 (.I(net119),
    .Z(wbs_dat_o[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output120 (.I(net120),
    .Z(wbs_dat_o[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output121 (.I(net121),
    .Z(wbs_dat_o[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output122 (.I(net122),
    .Z(wbs_dat_o[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output123 (.I(net123),
    .Z(wbs_dat_o[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output59 (.I(net59),
    .Z(io_oeb[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output60 (.I(net60),
    .Z(io_oeb[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output61 (.I(net61),
    .Z(io_oeb[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output62 (.I(net62),
    .Z(io_oeb[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output63 (.I(net63),
    .Z(io_oeb[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output64 (.I(net64),
    .Z(io_oeb[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output65 (.I(net138),
    .Z(io_oeb[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output66 (.I(net66),
    .Z(io_oeb[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output67 (.I(net67),
    .Z(io_oeb[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output68 (.I(net68),
    .Z(io_oeb[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output69 (.I(net69),
    .Z(io_oeb[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output70 (.I(net70),
    .Z(io_oeb[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output71 (.I(net71),
    .Z(io_oeb[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output72 (.I(net72),
    .Z(io_oeb[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output73 (.I(net73),
    .Z(io_oeb[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output74 (.I(net74),
    .Z(io_oeb[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output75 (.I(net75),
    .Z(io_out[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output76 (.I(net76),
    .Z(io_out[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output77 (.I(net77),
    .Z(io_out[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output78 (.I(net126),
    .Z(io_out[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output79 (.I(net79),
    .Z(io_out[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output80 (.I(net80),
    .Z(io_out[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output81 (.I(net81),
    .Z(io_out[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output82 (.I(net82),
    .Z(io_out[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output83 (.I(net137),
    .Z(io_out[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output84 (.I(net84),
    .Z(io_out[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output85 (.I(net134),
    .Z(io_out[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output86 (.I(net86),
    .Z(io_out[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output87 (.I(net131),
    .Z(io_out[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output88 (.I(net88),
    .Z(io_out[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output89 (.I(net89),
    .Z(io_out[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output90 (.I(net90),
    .Z(io_out[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output91 (.I(net91),
    .Z(la_data_out[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output92 (.I(net92),
    .Z(la_data_out[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output93 (.I(net93),
    .Z(la_data_out[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output94 (.I(net94),
    .Z(la_data_out[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output95 (.I(net95),
    .Z(la_data_out[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output96 (.I(net96),
    .Z(la_data_out[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output97 (.I(net97),
    .Z(la_data_out[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output98 (.I(net98),
    .Z(la_data_out[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output99 (.I(net99),
    .Z(la_data_out[2]));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_146 (.ZN(net146));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_147 (.ZN(net147));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_148 (.ZN(net148));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_149 (.ZN(net149));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_150 (.ZN(net150));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_151 (.ZN(net151));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_152 (.ZN(net152));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_153 (.ZN(net153));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_154 (.ZN(net154));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_155 (.ZN(net155));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_156 (.ZN(net156));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_157 (.ZN(net157));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_158 (.ZN(net158));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_159 (.ZN(net159));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_160 (.ZN(net160));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_161 (.ZN(net161));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_162 (.ZN(net162));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_163 (.ZN(net163));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_164 (.ZN(net164));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_165 (.ZN(net165));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_166 (.ZN(net166));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_167 (.ZN(net167));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_168 (.ZN(net168));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_169 (.ZN(net169));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_170 (.ZN(net170));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_171 (.ZN(net171));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_172 (.ZN(net172));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_173 (.ZN(net173));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_174 (.ZN(net174));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_175 (.ZN(net175));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_176 (.ZN(net176));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_177 (.ZN(net177));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_178 (.ZN(net178));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_179 (.ZN(net179));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_180 (.ZN(net180));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_181 (.ZN(net181));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_182 (.ZN(net182));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_183 (.ZN(net183));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_184 (.ZN(net184));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_185 (.ZN(net185));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_186 (.ZN(net186));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_187 (.ZN(net187));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_188 (.ZN(net188));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_189 (.ZN(net189));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_190 (.ZN(net190));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_191 (.ZN(net191));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_192 (.ZN(net192));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_193 (.ZN(net193));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_194 (.ZN(net194));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_195 (.ZN(net195));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_196 (.ZN(net196));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_197 (.ZN(net197));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_198 (.ZN(net198));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_199 (.ZN(net199));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_200 (.ZN(net200));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_201 (.ZN(net201));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_202 (.ZN(net202));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_203 (.ZN(net203));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_204 (.ZN(net204));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_205 (.ZN(net205));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_206 (.ZN(net206));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_207 (.ZN(net207));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_208 (.ZN(net208));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_209 (.ZN(net209));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_210 (.ZN(net210));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_211 (.ZN(net211));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_212 (.ZN(net212));
 assign irq[0] = net194;
 assign irq[1] = net195;
 assign irq[2] = net196;
 assign la_data_out[16] = net197;
 assign la_data_out[17] = net198;
 assign la_data_out[18] = net199;
 assign la_data_out[19] = net200;
 assign la_data_out[20] = net201;
 assign la_data_out[21] = net202;
 assign la_data_out[22] = net203;
 assign la_data_out[23] = net204;
 assign la_data_out[24] = net205;
 assign la_data_out[25] = net206;
 assign la_data_out[26] = net207;
 assign la_data_out[27] = net208;
 assign la_data_out[28] = net209;
 assign la_data_out[29] = net210;
 assign la_data_out[30] = net211;
 assign la_data_out[31] = net212;
 assign la_data_out[32] = net146;
 assign la_data_out[33] = net147;
 assign la_data_out[34] = net148;
 assign la_data_out[35] = net149;
 assign la_data_out[36] = net150;
 assign la_data_out[37] = net151;
 assign la_data_out[38] = net152;
 assign la_data_out[39] = net153;
 assign la_data_out[40] = net154;
 assign la_data_out[41] = net155;
 assign la_data_out[42] = net156;
 assign la_data_out[43] = net157;
 assign la_data_out[44] = net158;
 assign la_data_out[45] = net159;
 assign la_data_out[46] = net160;
 assign la_data_out[47] = net161;
 assign la_data_out[48] = net162;
 assign la_data_out[49] = net163;
 assign la_data_out[50] = net164;
 assign la_data_out[51] = net165;
 assign la_data_out[52] = net166;
 assign la_data_out[53] = net167;
 assign la_data_out[54] = net168;
 assign la_data_out[55] = net169;
 assign la_data_out[56] = net170;
 assign la_data_out[57] = net171;
 assign la_data_out[58] = net172;
 assign la_data_out[59] = net173;
 assign la_data_out[60] = net174;
 assign la_data_out[61] = net175;
 assign la_data_out[62] = net176;
 assign la_data_out[63] = net177;
 assign wbs_dat_o[16] = net178;
 assign wbs_dat_o[17] = net179;
 assign wbs_dat_o[18] = net180;
 assign wbs_dat_o[19] = net181;
 assign wbs_dat_o[20] = net182;
 assign wbs_dat_o[21] = net183;
 assign wbs_dat_o[22] = net184;
 assign wbs_dat_o[23] = net185;
 assign wbs_dat_o[24] = net186;
 assign wbs_dat_o[25] = net187;
 assign wbs_dat_o[26] = net188;
 assign wbs_dat_o[27] = net189;
 assign wbs_dat_o[28] = net190;
 assign wbs_dat_o[29] = net191;
 assign wbs_dat_o[30] = net192;
 assign wbs_dat_o[31] = net193;
endmodule

