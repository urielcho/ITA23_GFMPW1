VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO ita
  CLASS BLOCK ;
  FOREIGN ita ;
  ORIGIN 0.000 0.000 ;
  SIZE 320.000 BY 2702.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 10.080 0.000 10.640 4.000 ;
    END
  END clk
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 106.400 2698.000 106.960 2702.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 162.400 2698.000 162.960 2702.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 168.000 2698.000 168.560 2702.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 173.600 2698.000 174.160 2702.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 179.200 2698.000 179.760 2702.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 184.800 2698.000 185.360 2702.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 190.400 2698.000 190.960 2702.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 196.000 2698.000 196.560 2702.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 201.600 2698.000 202.160 2702.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 207.200 2698.000 207.760 2702.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 212.800 2698.000 213.360 2702.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 112.000 2698.000 112.560 2702.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 218.400 2698.000 218.960 2702.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 224.000 2698.000 224.560 2702.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 229.600 2698.000 230.160 2702.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 235.200 2698.000 235.760 2702.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 240.800 2698.000 241.360 2702.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 246.400 2698.000 246.960 2702.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 252.000 2698.000 252.560 2702.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 257.600 2698.000 258.160 2702.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 263.200 2698.000 263.760 2702.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 268.800 2698.000 269.360 2702.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 117.600 2698.000 118.160 2702.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 274.400 2698.000 274.960 2702.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 280.000 2698.000 280.560 2702.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 285.600 2698.000 286.160 2702.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 291.200 2698.000 291.760 2702.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 296.800 2698.000 297.360 2702.000 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 302.400 2698.000 302.960 2702.000 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 308.000 2698.000 308.560 2702.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 313.600 2698.000 314.160 2702.000 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 123.200 2698.000 123.760 2702.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 128.800 2698.000 129.360 2702.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 134.400 2698.000 134.960 2702.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 140.000 2698.000 140.560 2702.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 145.600 2698.000 146.160 2702.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 151.200 2698.000 151.760 2702.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 156.800 2698.000 157.360 2702.000 ;
    END
  END io_oeb[9]
  PIN itasegm[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 319.200 4.000 319.760 ;
    END
  END itasegm[0]
  PIN itasegm[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 442.400 320.000 442.960 ;
    END
  END itasegm[100]
  PIN itasegm[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 445.200 320.000 445.760 ;
    END
  END itasegm[101]
  PIN itasegm[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 448.000 320.000 448.560 ;
    END
  END itasegm[102]
  PIN itasegm[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 450.800 320.000 451.360 ;
    END
  END itasegm[103]
  PIN itasegm[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 453.600 320.000 454.160 ;
    END
  END itasegm[104]
  PIN itasegm[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 456.400 320.000 456.960 ;
    END
  END itasegm[105]
  PIN itasegm[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 459.200 320.000 459.760 ;
    END
  END itasegm[106]
  PIN itasegm[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 462.000 320.000 462.560 ;
    END
  END itasegm[107]
  PIN itasegm[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 464.800 320.000 465.360 ;
    END
  END itasegm[108]
  PIN itasegm[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 467.600 320.000 468.160 ;
    END
  END itasegm[109]
  PIN itasegm[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 347.200 4.000 347.760 ;
    END
  END itasegm[10]
  PIN itasegm[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 470.400 320.000 470.960 ;
    END
  END itasegm[110]
  PIN itasegm[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 473.200 320.000 473.760 ;
    END
  END itasegm[111]
  PIN itasegm[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 610.400 4.000 610.960 ;
    END
  END itasegm[112]
  PIN itasegm[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 613.200 4.000 613.760 ;
    END
  END itasegm[113]
  PIN itasegm[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 616.000 4.000 616.560 ;
    END
  END itasegm[114]
  PIN itasegm[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 618.800 4.000 619.360 ;
    END
  END itasegm[115]
  PIN itasegm[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 621.600 4.000 622.160 ;
    END
  END itasegm[116]
  PIN itasegm[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 624.400 4.000 624.960 ;
    END
  END itasegm[117]
  PIN itasegm[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 627.200 4.000 627.760 ;
    END
  END itasegm[118]
  PIN itasegm[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 630.000 4.000 630.560 ;
    END
  END itasegm[119]
  PIN itasegm[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 350.000 4.000 350.560 ;
    END
  END itasegm[11]
  PIN itasegm[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 632.800 4.000 633.360 ;
    END
  END itasegm[120]
  PIN itasegm[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 635.600 4.000 636.160 ;
    END
  END itasegm[121]
  PIN itasegm[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 638.400 4.000 638.960 ;
    END
  END itasegm[122]
  PIN itasegm[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 641.200 4.000 641.760 ;
    END
  END itasegm[123]
  PIN itasegm[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 644.000 4.000 644.560 ;
    END
  END itasegm[124]
  PIN itasegm[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 646.800 4.000 647.360 ;
    END
  END itasegm[125]
  PIN itasegm[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 649.600 4.000 650.160 ;
    END
  END itasegm[126]
  PIN itasegm[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 652.400 4.000 652.960 ;
    END
  END itasegm[127]
  PIN itasegm[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 655.200 4.000 655.760 ;
    END
  END itasegm[128]
  PIN itasegm[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 658.000 4.000 658.560 ;
    END
  END itasegm[129]
  PIN itasegm[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 352.800 4.000 353.360 ;
    END
  END itasegm[12]
  PIN itasegm[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 660.800 4.000 661.360 ;
    END
  END itasegm[130]
  PIN itasegm[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 663.600 4.000 664.160 ;
    END
  END itasegm[131]
  PIN itasegm[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 666.400 4.000 666.960 ;
    END
  END itasegm[132]
  PIN itasegm[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 669.200 4.000 669.760 ;
    END
  END itasegm[133]
  PIN itasegm[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 672.000 4.000 672.560 ;
    END
  END itasegm[134]
  PIN itasegm[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 674.800 4.000 675.360 ;
    END
  END itasegm[135]
  PIN itasegm[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 677.600 4.000 678.160 ;
    END
  END itasegm[136]
  PIN itasegm[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 680.400 4.000 680.960 ;
    END
  END itasegm[137]
  PIN itasegm[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 683.200 4.000 683.760 ;
    END
  END itasegm[138]
  PIN itasegm[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 686.000 4.000 686.560 ;
    END
  END itasegm[139]
  PIN itasegm[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 355.600 4.000 356.160 ;
    END
  END itasegm[13]
  PIN itasegm[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 688.800 4.000 689.360 ;
    END
  END itasegm[140]
  PIN itasegm[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 691.600 4.000 692.160 ;
    END
  END itasegm[141]
  PIN itasegm[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 694.400 4.000 694.960 ;
    END
  END itasegm[142]
  PIN itasegm[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 697.200 4.000 697.760 ;
    END
  END itasegm[143]
  PIN itasegm[144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 700.000 4.000 700.560 ;
    END
  END itasegm[144]
  PIN itasegm[145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 702.800 4.000 703.360 ;
    END
  END itasegm[145]
  PIN itasegm[146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 705.600 4.000 706.160 ;
    END
  END itasegm[146]
  PIN itasegm[147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 708.400 4.000 708.960 ;
    END
  END itasegm[147]
  PIN itasegm[148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 711.200 4.000 711.760 ;
    END
  END itasegm[148]
  PIN itasegm[149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 714.000 4.000 714.560 ;
    END
  END itasegm[149]
  PIN itasegm[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 358.400 4.000 358.960 ;
    END
  END itasegm[14]
  PIN itasegm[150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 716.800 4.000 717.360 ;
    END
  END itasegm[150]
  PIN itasegm[151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 719.600 4.000 720.160 ;
    END
  END itasegm[151]
  PIN itasegm[152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 722.400 4.000 722.960 ;
    END
  END itasegm[152]
  PIN itasegm[153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 725.200 4.000 725.760 ;
    END
  END itasegm[153]
  PIN itasegm[154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 728.000 4.000 728.560 ;
    END
  END itasegm[154]
  PIN itasegm[155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 730.800 4.000 731.360 ;
    END
  END itasegm[155]
  PIN itasegm[156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 733.600 4.000 734.160 ;
    END
  END itasegm[156]
  PIN itasegm[157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 736.400 4.000 736.960 ;
    END
  END itasegm[157]
  PIN itasegm[158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 739.200 4.000 739.760 ;
    END
  END itasegm[158]
  PIN itasegm[159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 742.000 4.000 742.560 ;
    END
  END itasegm[159]
  PIN itasegm[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 361.200 4.000 361.760 ;
    END
  END itasegm[15]
  PIN itasegm[160]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 744.800 4.000 745.360 ;
    END
  END itasegm[160]
  PIN itasegm[161]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 747.600 4.000 748.160 ;
    END
  END itasegm[161]
  PIN itasegm[162]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 750.400 4.000 750.960 ;
    END
  END itasegm[162]
  PIN itasegm[163]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 753.200 4.000 753.760 ;
    END
  END itasegm[163]
  PIN itasegm[164]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 756.000 4.000 756.560 ;
    END
  END itasegm[164]
  PIN itasegm[165]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 758.800 4.000 759.360 ;
    END
  END itasegm[165]
  PIN itasegm[166]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 761.600 4.000 762.160 ;
    END
  END itasegm[166]
  PIN itasegm[167]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 764.400 4.000 764.960 ;
    END
  END itasegm[167]
  PIN itasegm[168]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 610.400 320.000 610.960 ;
    END
  END itasegm[168]
  PIN itasegm[169]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 613.200 320.000 613.760 ;
    END
  END itasegm[169]
  PIN itasegm[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 364.000 4.000 364.560 ;
    END
  END itasegm[16]
  PIN itasegm[170]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 616.000 320.000 616.560 ;
    END
  END itasegm[170]
  PIN itasegm[171]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 618.800 320.000 619.360 ;
    END
  END itasegm[171]
  PIN itasegm[172]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 621.600 320.000 622.160 ;
    END
  END itasegm[172]
  PIN itasegm[173]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 624.400 320.000 624.960 ;
    END
  END itasegm[173]
  PIN itasegm[174]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 627.200 320.000 627.760 ;
    END
  END itasegm[174]
  PIN itasegm[175]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 630.000 320.000 630.560 ;
    END
  END itasegm[175]
  PIN itasegm[176]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 632.800 320.000 633.360 ;
    END
  END itasegm[176]
  PIN itasegm[177]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 635.600 320.000 636.160 ;
    END
  END itasegm[177]
  PIN itasegm[178]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 638.400 320.000 638.960 ;
    END
  END itasegm[178]
  PIN itasegm[179]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 641.200 320.000 641.760 ;
    END
  END itasegm[179]
  PIN itasegm[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 366.800 4.000 367.360 ;
    END
  END itasegm[17]
  PIN itasegm[180]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 644.000 320.000 644.560 ;
    END
  END itasegm[180]
  PIN itasegm[181]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 646.800 320.000 647.360 ;
    END
  END itasegm[181]
  PIN itasegm[182]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 649.600 320.000 650.160 ;
    END
  END itasegm[182]
  PIN itasegm[183]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 652.400 320.000 652.960 ;
    END
  END itasegm[183]
  PIN itasegm[184]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 655.200 320.000 655.760 ;
    END
  END itasegm[184]
  PIN itasegm[185]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 658.000 320.000 658.560 ;
    END
  END itasegm[185]
  PIN itasegm[186]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 660.800 320.000 661.360 ;
    END
  END itasegm[186]
  PIN itasegm[187]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 663.600 320.000 664.160 ;
    END
  END itasegm[187]
  PIN itasegm[188]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 666.400 320.000 666.960 ;
    END
  END itasegm[188]
  PIN itasegm[189]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 669.200 320.000 669.760 ;
    END
  END itasegm[189]
  PIN itasegm[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 369.600 4.000 370.160 ;
    END
  END itasegm[18]
  PIN itasegm[190]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 672.000 320.000 672.560 ;
    END
  END itasegm[190]
  PIN itasegm[191]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 674.800 320.000 675.360 ;
    END
  END itasegm[191]
  PIN itasegm[192]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 677.600 320.000 678.160 ;
    END
  END itasegm[192]
  PIN itasegm[193]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 680.400 320.000 680.960 ;
    END
  END itasegm[193]
  PIN itasegm[194]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 683.200 320.000 683.760 ;
    END
  END itasegm[194]
  PIN itasegm[195]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 686.000 320.000 686.560 ;
    END
  END itasegm[195]
  PIN itasegm[196]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 688.800 320.000 689.360 ;
    END
  END itasegm[196]
  PIN itasegm[197]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 691.600 320.000 692.160 ;
    END
  END itasegm[197]
  PIN itasegm[198]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 694.400 320.000 694.960 ;
    END
  END itasegm[198]
  PIN itasegm[199]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 697.200 320.000 697.760 ;
    END
  END itasegm[199]
  PIN itasegm[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 372.400 4.000 372.960 ;
    END
  END itasegm[19]
  PIN itasegm[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 322.000 4.000 322.560 ;
    END
  END itasegm[1]
  PIN itasegm[200]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 700.000 320.000 700.560 ;
    END
  END itasegm[200]
  PIN itasegm[201]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 702.800 320.000 703.360 ;
    END
  END itasegm[201]
  PIN itasegm[202]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 705.600 320.000 706.160 ;
    END
  END itasegm[202]
  PIN itasegm[203]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 708.400 320.000 708.960 ;
    END
  END itasegm[203]
  PIN itasegm[204]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 711.200 320.000 711.760 ;
    END
  END itasegm[204]
  PIN itasegm[205]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 714.000 320.000 714.560 ;
    END
  END itasegm[205]
  PIN itasegm[206]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 716.800 320.000 717.360 ;
    END
  END itasegm[206]
  PIN itasegm[207]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 719.600 320.000 720.160 ;
    END
  END itasegm[207]
  PIN itasegm[208]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 722.400 320.000 722.960 ;
    END
  END itasegm[208]
  PIN itasegm[209]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 725.200 320.000 725.760 ;
    END
  END itasegm[209]
  PIN itasegm[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 375.200 4.000 375.760 ;
    END
  END itasegm[20]
  PIN itasegm[210]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 728.000 320.000 728.560 ;
    END
  END itasegm[210]
  PIN itasegm[211]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 730.800 320.000 731.360 ;
    END
  END itasegm[211]
  PIN itasegm[212]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 733.600 320.000 734.160 ;
    END
  END itasegm[212]
  PIN itasegm[213]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 736.400 320.000 736.960 ;
    END
  END itasegm[213]
  PIN itasegm[214]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 739.200 320.000 739.760 ;
    END
  END itasegm[214]
  PIN itasegm[215]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 742.000 320.000 742.560 ;
    END
  END itasegm[215]
  PIN itasegm[216]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 744.800 320.000 745.360 ;
    END
  END itasegm[216]
  PIN itasegm[217]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 747.600 320.000 748.160 ;
    END
  END itasegm[217]
  PIN itasegm[218]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 750.400 320.000 750.960 ;
    END
  END itasegm[218]
  PIN itasegm[219]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 753.200 320.000 753.760 ;
    END
  END itasegm[219]
  PIN itasegm[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 378.000 4.000 378.560 ;
    END
  END itasegm[21]
  PIN itasegm[220]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 756.000 320.000 756.560 ;
    END
  END itasegm[220]
  PIN itasegm[221]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 758.800 320.000 759.360 ;
    END
  END itasegm[221]
  PIN itasegm[222]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 761.600 320.000 762.160 ;
    END
  END itasegm[222]
  PIN itasegm[223]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 764.400 320.000 764.960 ;
    END
  END itasegm[223]
  PIN itasegm[224]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 901.600 4.000 902.160 ;
    END
  END itasegm[224]
  PIN itasegm[225]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 904.400 4.000 904.960 ;
    END
  END itasegm[225]
  PIN itasegm[226]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 907.200 4.000 907.760 ;
    END
  END itasegm[226]
  PIN itasegm[227]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 910.000 4.000 910.560 ;
    END
  END itasegm[227]
  PIN itasegm[228]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 912.800 4.000 913.360 ;
    END
  END itasegm[228]
  PIN itasegm[229]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 915.600 4.000 916.160 ;
    END
  END itasegm[229]
  PIN itasegm[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 380.800 4.000 381.360 ;
    END
  END itasegm[22]
  PIN itasegm[230]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 918.400 4.000 918.960 ;
    END
  END itasegm[230]
  PIN itasegm[231]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 921.200 4.000 921.760 ;
    END
  END itasegm[231]
  PIN itasegm[232]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 924.000 4.000 924.560 ;
    END
  END itasegm[232]
  PIN itasegm[233]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 926.800 4.000 927.360 ;
    END
  END itasegm[233]
  PIN itasegm[234]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 929.600 4.000 930.160 ;
    END
  END itasegm[234]
  PIN itasegm[235]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 932.400 4.000 932.960 ;
    END
  END itasegm[235]
  PIN itasegm[236]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 935.200 4.000 935.760 ;
    END
  END itasegm[236]
  PIN itasegm[237]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 938.000 4.000 938.560 ;
    END
  END itasegm[237]
  PIN itasegm[238]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 940.800 4.000 941.360 ;
    END
  END itasegm[238]
  PIN itasegm[239]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 943.600 4.000 944.160 ;
    END
  END itasegm[239]
  PIN itasegm[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 383.600 4.000 384.160 ;
    END
  END itasegm[23]
  PIN itasegm[240]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 946.400 4.000 946.960 ;
    END
  END itasegm[240]
  PIN itasegm[241]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 949.200 4.000 949.760 ;
    END
  END itasegm[241]
  PIN itasegm[242]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 952.000 4.000 952.560 ;
    END
  END itasegm[242]
  PIN itasegm[243]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 954.800 4.000 955.360 ;
    END
  END itasegm[243]
  PIN itasegm[244]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 957.600 4.000 958.160 ;
    END
  END itasegm[244]
  PIN itasegm[245]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 960.400 4.000 960.960 ;
    END
  END itasegm[245]
  PIN itasegm[246]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 963.200 4.000 963.760 ;
    END
  END itasegm[246]
  PIN itasegm[247]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 966.000 4.000 966.560 ;
    END
  END itasegm[247]
  PIN itasegm[248]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 968.800 4.000 969.360 ;
    END
  END itasegm[248]
  PIN itasegm[249]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 971.600 4.000 972.160 ;
    END
  END itasegm[249]
  PIN itasegm[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 386.400 4.000 386.960 ;
    END
  END itasegm[24]
  PIN itasegm[250]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 974.400 4.000 974.960 ;
    END
  END itasegm[250]
  PIN itasegm[251]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 977.200 4.000 977.760 ;
    END
  END itasegm[251]
  PIN itasegm[252]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 980.000 4.000 980.560 ;
    END
  END itasegm[252]
  PIN itasegm[253]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 982.800 4.000 983.360 ;
    END
  END itasegm[253]
  PIN itasegm[254]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 985.600 4.000 986.160 ;
    END
  END itasegm[254]
  PIN itasegm[255]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 988.400 4.000 988.960 ;
    END
  END itasegm[255]
  PIN itasegm[256]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 991.200 4.000 991.760 ;
    END
  END itasegm[256]
  PIN itasegm[257]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 994.000 4.000 994.560 ;
    END
  END itasegm[257]
  PIN itasegm[258]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 996.800 4.000 997.360 ;
    END
  END itasegm[258]
  PIN itasegm[259]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 999.600 4.000 1000.160 ;
    END
  END itasegm[259]
  PIN itasegm[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 389.200 4.000 389.760 ;
    END
  END itasegm[25]
  PIN itasegm[260]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1002.400 4.000 1002.960 ;
    END
  END itasegm[260]
  PIN itasegm[261]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1005.200 4.000 1005.760 ;
    END
  END itasegm[261]
  PIN itasegm[262]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1008.000 4.000 1008.560 ;
    END
  END itasegm[262]
  PIN itasegm[263]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1010.800 4.000 1011.360 ;
    END
  END itasegm[263]
  PIN itasegm[264]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1013.600 4.000 1014.160 ;
    END
  END itasegm[264]
  PIN itasegm[265]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1016.400 4.000 1016.960 ;
    END
  END itasegm[265]
  PIN itasegm[266]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1019.200 4.000 1019.760 ;
    END
  END itasegm[266]
  PIN itasegm[267]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1022.000 4.000 1022.560 ;
    END
  END itasegm[267]
  PIN itasegm[268]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1024.800 4.000 1025.360 ;
    END
  END itasegm[268]
  PIN itasegm[269]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1027.600 4.000 1028.160 ;
    END
  END itasegm[269]
  PIN itasegm[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 392.000 4.000 392.560 ;
    END
  END itasegm[26]
  PIN itasegm[270]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1030.400 4.000 1030.960 ;
    END
  END itasegm[270]
  PIN itasegm[271]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1033.200 4.000 1033.760 ;
    END
  END itasegm[271]
  PIN itasegm[272]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1036.000 4.000 1036.560 ;
    END
  END itasegm[272]
  PIN itasegm[273]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1038.800 4.000 1039.360 ;
    END
  END itasegm[273]
  PIN itasegm[274]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1041.600 4.000 1042.160 ;
    END
  END itasegm[274]
  PIN itasegm[275]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1044.400 4.000 1044.960 ;
    END
  END itasegm[275]
  PIN itasegm[276]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1047.200 4.000 1047.760 ;
    END
  END itasegm[276]
  PIN itasegm[277]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1050.000 4.000 1050.560 ;
    END
  END itasegm[277]
  PIN itasegm[278]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1052.800 4.000 1053.360 ;
    END
  END itasegm[278]
  PIN itasegm[279]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1055.600 4.000 1056.160 ;
    END
  END itasegm[279]
  PIN itasegm[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 394.800 4.000 395.360 ;
    END
  END itasegm[27]
  PIN itasegm[280]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 901.600 320.000 902.160 ;
    END
  END itasegm[280]
  PIN itasegm[281]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 904.400 320.000 904.960 ;
    END
  END itasegm[281]
  PIN itasegm[282]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 907.200 320.000 907.760 ;
    END
  END itasegm[282]
  PIN itasegm[283]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 910.000 320.000 910.560 ;
    END
  END itasegm[283]
  PIN itasegm[284]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 912.800 320.000 913.360 ;
    END
  END itasegm[284]
  PIN itasegm[285]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 915.600 320.000 916.160 ;
    END
  END itasegm[285]
  PIN itasegm[286]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 918.400 320.000 918.960 ;
    END
  END itasegm[286]
  PIN itasegm[287]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 921.200 320.000 921.760 ;
    END
  END itasegm[287]
  PIN itasegm[288]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 924.000 320.000 924.560 ;
    END
  END itasegm[288]
  PIN itasegm[289]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 926.800 320.000 927.360 ;
    END
  END itasegm[289]
  PIN itasegm[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 397.600 4.000 398.160 ;
    END
  END itasegm[28]
  PIN itasegm[290]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 929.600 320.000 930.160 ;
    END
  END itasegm[290]
  PIN itasegm[291]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 932.400 320.000 932.960 ;
    END
  END itasegm[291]
  PIN itasegm[292]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 935.200 320.000 935.760 ;
    END
  END itasegm[292]
  PIN itasegm[293]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 938.000 320.000 938.560 ;
    END
  END itasegm[293]
  PIN itasegm[294]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 940.800 320.000 941.360 ;
    END
  END itasegm[294]
  PIN itasegm[295]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 943.600 320.000 944.160 ;
    END
  END itasegm[295]
  PIN itasegm[296]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 946.400 320.000 946.960 ;
    END
  END itasegm[296]
  PIN itasegm[297]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 949.200 320.000 949.760 ;
    END
  END itasegm[297]
  PIN itasegm[298]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 952.000 320.000 952.560 ;
    END
  END itasegm[298]
  PIN itasegm[299]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 954.800 320.000 955.360 ;
    END
  END itasegm[299]
  PIN itasegm[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 400.400 4.000 400.960 ;
    END
  END itasegm[29]
  PIN itasegm[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 324.800 4.000 325.360 ;
    END
  END itasegm[2]
  PIN itasegm[300]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 957.600 320.000 958.160 ;
    END
  END itasegm[300]
  PIN itasegm[301]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 960.400 320.000 960.960 ;
    END
  END itasegm[301]
  PIN itasegm[302]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 963.200 320.000 963.760 ;
    END
  END itasegm[302]
  PIN itasegm[303]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 966.000 320.000 966.560 ;
    END
  END itasegm[303]
  PIN itasegm[304]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 968.800 320.000 969.360 ;
    END
  END itasegm[304]
  PIN itasegm[305]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 971.600 320.000 972.160 ;
    END
  END itasegm[305]
  PIN itasegm[306]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 974.400 320.000 974.960 ;
    END
  END itasegm[306]
  PIN itasegm[307]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 977.200 320.000 977.760 ;
    END
  END itasegm[307]
  PIN itasegm[308]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 980.000 320.000 980.560 ;
    END
  END itasegm[308]
  PIN itasegm[309]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 982.800 320.000 983.360 ;
    END
  END itasegm[309]
  PIN itasegm[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 403.200 4.000 403.760 ;
    END
  END itasegm[30]
  PIN itasegm[310]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 985.600 320.000 986.160 ;
    END
  END itasegm[310]
  PIN itasegm[311]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 988.400 320.000 988.960 ;
    END
  END itasegm[311]
  PIN itasegm[312]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 991.200 320.000 991.760 ;
    END
  END itasegm[312]
  PIN itasegm[313]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 994.000 320.000 994.560 ;
    END
  END itasegm[313]
  PIN itasegm[314]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 996.800 320.000 997.360 ;
    END
  END itasegm[314]
  PIN itasegm[315]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 999.600 320.000 1000.160 ;
    END
  END itasegm[315]
  PIN itasegm[316]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1002.400 320.000 1002.960 ;
    END
  END itasegm[316]
  PIN itasegm[317]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1005.200 320.000 1005.760 ;
    END
  END itasegm[317]
  PIN itasegm[318]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1008.000 320.000 1008.560 ;
    END
  END itasegm[318]
  PIN itasegm[319]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1010.800 320.000 1011.360 ;
    END
  END itasegm[319]
  PIN itasegm[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 406.000 4.000 406.560 ;
    END
  END itasegm[31]
  PIN itasegm[320]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1013.600 320.000 1014.160 ;
    END
  END itasegm[320]
  PIN itasegm[321]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1016.400 320.000 1016.960 ;
    END
  END itasegm[321]
  PIN itasegm[322]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1019.200 320.000 1019.760 ;
    END
  END itasegm[322]
  PIN itasegm[323]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1022.000 320.000 1022.560 ;
    END
  END itasegm[323]
  PIN itasegm[324]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1024.800 320.000 1025.360 ;
    END
  END itasegm[324]
  PIN itasegm[325]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1027.600 320.000 1028.160 ;
    END
  END itasegm[325]
  PIN itasegm[326]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1030.400 320.000 1030.960 ;
    END
  END itasegm[326]
  PIN itasegm[327]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1033.200 320.000 1033.760 ;
    END
  END itasegm[327]
  PIN itasegm[328]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1036.000 320.000 1036.560 ;
    END
  END itasegm[328]
  PIN itasegm[329]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1038.800 320.000 1039.360 ;
    END
  END itasegm[329]
  PIN itasegm[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 408.800 4.000 409.360 ;
    END
  END itasegm[32]
  PIN itasegm[330]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1041.600 320.000 1042.160 ;
    END
  END itasegm[330]
  PIN itasegm[331]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1044.400 320.000 1044.960 ;
    END
  END itasegm[331]
  PIN itasegm[332]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1047.200 320.000 1047.760 ;
    END
  END itasegm[332]
  PIN itasegm[333]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1050.000 320.000 1050.560 ;
    END
  END itasegm[333]
  PIN itasegm[334]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1052.800 320.000 1053.360 ;
    END
  END itasegm[334]
  PIN itasegm[335]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1055.600 320.000 1056.160 ;
    END
  END itasegm[335]
  PIN itasegm[336]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1192.800 4.000 1193.360 ;
    END
  END itasegm[336]
  PIN itasegm[337]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1195.600 4.000 1196.160 ;
    END
  END itasegm[337]
  PIN itasegm[338]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1198.400 4.000 1198.960 ;
    END
  END itasegm[338]
  PIN itasegm[339]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1201.200 4.000 1201.760 ;
    END
  END itasegm[339]
  PIN itasegm[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 411.600 4.000 412.160 ;
    END
  END itasegm[33]
  PIN itasegm[340]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1204.000 4.000 1204.560 ;
    END
  END itasegm[340]
  PIN itasegm[341]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1206.800 4.000 1207.360 ;
    END
  END itasegm[341]
  PIN itasegm[342]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1209.600 4.000 1210.160 ;
    END
  END itasegm[342]
  PIN itasegm[343]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1212.400 4.000 1212.960 ;
    END
  END itasegm[343]
  PIN itasegm[344]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1215.200 4.000 1215.760 ;
    END
  END itasegm[344]
  PIN itasegm[345]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1218.000 4.000 1218.560 ;
    END
  END itasegm[345]
  PIN itasegm[346]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1220.800 4.000 1221.360 ;
    END
  END itasegm[346]
  PIN itasegm[347]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1223.600 4.000 1224.160 ;
    END
  END itasegm[347]
  PIN itasegm[348]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1226.400 4.000 1226.960 ;
    END
  END itasegm[348]
  PIN itasegm[349]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1229.200 4.000 1229.760 ;
    END
  END itasegm[349]
  PIN itasegm[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 414.400 4.000 414.960 ;
    END
  END itasegm[34]
  PIN itasegm[350]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1232.000 4.000 1232.560 ;
    END
  END itasegm[350]
  PIN itasegm[351]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1234.800 4.000 1235.360 ;
    END
  END itasegm[351]
  PIN itasegm[352]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1237.600 4.000 1238.160 ;
    END
  END itasegm[352]
  PIN itasegm[353]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1240.400 4.000 1240.960 ;
    END
  END itasegm[353]
  PIN itasegm[354]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1243.200 4.000 1243.760 ;
    END
  END itasegm[354]
  PIN itasegm[355]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1246.000 4.000 1246.560 ;
    END
  END itasegm[355]
  PIN itasegm[356]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1248.800 4.000 1249.360 ;
    END
  END itasegm[356]
  PIN itasegm[357]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1251.600 4.000 1252.160 ;
    END
  END itasegm[357]
  PIN itasegm[358]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1254.400 4.000 1254.960 ;
    END
  END itasegm[358]
  PIN itasegm[359]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1257.200 4.000 1257.760 ;
    END
  END itasegm[359]
  PIN itasegm[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 417.200 4.000 417.760 ;
    END
  END itasegm[35]
  PIN itasegm[360]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1260.000 4.000 1260.560 ;
    END
  END itasegm[360]
  PIN itasegm[361]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1262.800 4.000 1263.360 ;
    END
  END itasegm[361]
  PIN itasegm[362]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1265.600 4.000 1266.160 ;
    END
  END itasegm[362]
  PIN itasegm[363]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1268.400 4.000 1268.960 ;
    END
  END itasegm[363]
  PIN itasegm[364]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1271.200 4.000 1271.760 ;
    END
  END itasegm[364]
  PIN itasegm[365]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1274.000 4.000 1274.560 ;
    END
  END itasegm[365]
  PIN itasegm[366]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1276.800 4.000 1277.360 ;
    END
  END itasegm[366]
  PIN itasegm[367]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1279.600 4.000 1280.160 ;
    END
  END itasegm[367]
  PIN itasegm[368]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1282.400 4.000 1282.960 ;
    END
  END itasegm[368]
  PIN itasegm[369]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1285.200 4.000 1285.760 ;
    END
  END itasegm[369]
  PIN itasegm[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 420.000 4.000 420.560 ;
    END
  END itasegm[36]
  PIN itasegm[370]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1288.000 4.000 1288.560 ;
    END
  END itasegm[370]
  PIN itasegm[371]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1290.800 4.000 1291.360 ;
    END
  END itasegm[371]
  PIN itasegm[372]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1293.600 4.000 1294.160 ;
    END
  END itasegm[372]
  PIN itasegm[373]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1296.400 4.000 1296.960 ;
    END
  END itasegm[373]
  PIN itasegm[374]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1299.200 4.000 1299.760 ;
    END
  END itasegm[374]
  PIN itasegm[375]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1302.000 4.000 1302.560 ;
    END
  END itasegm[375]
  PIN itasegm[376]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1304.800 4.000 1305.360 ;
    END
  END itasegm[376]
  PIN itasegm[377]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1307.600 4.000 1308.160 ;
    END
  END itasegm[377]
  PIN itasegm[378]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1310.400 4.000 1310.960 ;
    END
  END itasegm[378]
  PIN itasegm[379]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1313.200 4.000 1313.760 ;
    END
  END itasegm[379]
  PIN itasegm[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 422.800 4.000 423.360 ;
    END
  END itasegm[37]
  PIN itasegm[380]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1316.000 4.000 1316.560 ;
    END
  END itasegm[380]
  PIN itasegm[381]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1318.800 4.000 1319.360 ;
    END
  END itasegm[381]
  PIN itasegm[382]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1321.600 4.000 1322.160 ;
    END
  END itasegm[382]
  PIN itasegm[383]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1324.400 4.000 1324.960 ;
    END
  END itasegm[383]
  PIN itasegm[384]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1327.200 4.000 1327.760 ;
    END
  END itasegm[384]
  PIN itasegm[385]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1330.000 4.000 1330.560 ;
    END
  END itasegm[385]
  PIN itasegm[386]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1332.800 4.000 1333.360 ;
    END
  END itasegm[386]
  PIN itasegm[387]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1335.600 4.000 1336.160 ;
    END
  END itasegm[387]
  PIN itasegm[388]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1338.400 4.000 1338.960 ;
    END
  END itasegm[388]
  PIN itasegm[389]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1341.200 4.000 1341.760 ;
    END
  END itasegm[389]
  PIN itasegm[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 425.600 4.000 426.160 ;
    END
  END itasegm[38]
  PIN itasegm[390]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1344.000 4.000 1344.560 ;
    END
  END itasegm[390]
  PIN itasegm[391]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1346.800 4.000 1347.360 ;
    END
  END itasegm[391]
  PIN itasegm[392]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1192.800 320.000 1193.360 ;
    END
  END itasegm[392]
  PIN itasegm[393]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1195.600 320.000 1196.160 ;
    END
  END itasegm[393]
  PIN itasegm[394]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1198.400 320.000 1198.960 ;
    END
  END itasegm[394]
  PIN itasegm[395]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1201.200 320.000 1201.760 ;
    END
  END itasegm[395]
  PIN itasegm[396]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1204.000 320.000 1204.560 ;
    END
  END itasegm[396]
  PIN itasegm[397]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1206.800 320.000 1207.360 ;
    END
  END itasegm[397]
  PIN itasegm[398]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1209.600 320.000 1210.160 ;
    END
  END itasegm[398]
  PIN itasegm[399]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1212.400 320.000 1212.960 ;
    END
  END itasegm[399]
  PIN itasegm[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 428.400 4.000 428.960 ;
    END
  END itasegm[39]
  PIN itasegm[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 327.600 4.000 328.160 ;
    END
  END itasegm[3]
  PIN itasegm[400]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1215.200 320.000 1215.760 ;
    END
  END itasegm[400]
  PIN itasegm[401]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1218.000 320.000 1218.560 ;
    END
  END itasegm[401]
  PIN itasegm[402]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1220.800 320.000 1221.360 ;
    END
  END itasegm[402]
  PIN itasegm[403]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1223.600 320.000 1224.160 ;
    END
  END itasegm[403]
  PIN itasegm[404]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1226.400 320.000 1226.960 ;
    END
  END itasegm[404]
  PIN itasegm[405]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1229.200 320.000 1229.760 ;
    END
  END itasegm[405]
  PIN itasegm[406]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1232.000 320.000 1232.560 ;
    END
  END itasegm[406]
  PIN itasegm[407]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1234.800 320.000 1235.360 ;
    END
  END itasegm[407]
  PIN itasegm[408]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1237.600 320.000 1238.160 ;
    END
  END itasegm[408]
  PIN itasegm[409]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1240.400 320.000 1240.960 ;
    END
  END itasegm[409]
  PIN itasegm[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 431.200 4.000 431.760 ;
    END
  END itasegm[40]
  PIN itasegm[410]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1243.200 320.000 1243.760 ;
    END
  END itasegm[410]
  PIN itasegm[411]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1246.000 320.000 1246.560 ;
    END
  END itasegm[411]
  PIN itasegm[412]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1248.800 320.000 1249.360 ;
    END
  END itasegm[412]
  PIN itasegm[413]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1251.600 320.000 1252.160 ;
    END
  END itasegm[413]
  PIN itasegm[414]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1254.400 320.000 1254.960 ;
    END
  END itasegm[414]
  PIN itasegm[415]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1257.200 320.000 1257.760 ;
    END
  END itasegm[415]
  PIN itasegm[416]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1260.000 320.000 1260.560 ;
    END
  END itasegm[416]
  PIN itasegm[417]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1262.800 320.000 1263.360 ;
    END
  END itasegm[417]
  PIN itasegm[418]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1265.600 320.000 1266.160 ;
    END
  END itasegm[418]
  PIN itasegm[419]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1268.400 320.000 1268.960 ;
    END
  END itasegm[419]
  PIN itasegm[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 434.000 4.000 434.560 ;
    END
  END itasegm[41]
  PIN itasegm[420]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1271.200 320.000 1271.760 ;
    END
  END itasegm[420]
  PIN itasegm[421]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1274.000 320.000 1274.560 ;
    END
  END itasegm[421]
  PIN itasegm[422]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1276.800 320.000 1277.360 ;
    END
  END itasegm[422]
  PIN itasegm[423]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1279.600 320.000 1280.160 ;
    END
  END itasegm[423]
  PIN itasegm[424]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1282.400 320.000 1282.960 ;
    END
  END itasegm[424]
  PIN itasegm[425]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1285.200 320.000 1285.760 ;
    END
  END itasegm[425]
  PIN itasegm[426]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1288.000 320.000 1288.560 ;
    END
  END itasegm[426]
  PIN itasegm[427]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1290.800 320.000 1291.360 ;
    END
  END itasegm[427]
  PIN itasegm[428]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1293.600 320.000 1294.160 ;
    END
  END itasegm[428]
  PIN itasegm[429]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1296.400 320.000 1296.960 ;
    END
  END itasegm[429]
  PIN itasegm[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 436.800 4.000 437.360 ;
    END
  END itasegm[42]
  PIN itasegm[430]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1299.200 320.000 1299.760 ;
    END
  END itasegm[430]
  PIN itasegm[431]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1302.000 320.000 1302.560 ;
    END
  END itasegm[431]
  PIN itasegm[432]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1304.800 320.000 1305.360 ;
    END
  END itasegm[432]
  PIN itasegm[433]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1307.600 320.000 1308.160 ;
    END
  END itasegm[433]
  PIN itasegm[434]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1310.400 320.000 1310.960 ;
    END
  END itasegm[434]
  PIN itasegm[435]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1313.200 320.000 1313.760 ;
    END
  END itasegm[435]
  PIN itasegm[436]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1316.000 320.000 1316.560 ;
    END
  END itasegm[436]
  PIN itasegm[437]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1318.800 320.000 1319.360 ;
    END
  END itasegm[437]
  PIN itasegm[438]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1321.600 320.000 1322.160 ;
    END
  END itasegm[438]
  PIN itasegm[439]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1324.400 320.000 1324.960 ;
    END
  END itasegm[439]
  PIN itasegm[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 439.600 4.000 440.160 ;
    END
  END itasegm[43]
  PIN itasegm[440]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1327.200 320.000 1327.760 ;
    END
  END itasegm[440]
  PIN itasegm[441]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1330.000 320.000 1330.560 ;
    END
  END itasegm[441]
  PIN itasegm[442]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1332.800 320.000 1333.360 ;
    END
  END itasegm[442]
  PIN itasegm[443]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1335.600 320.000 1336.160 ;
    END
  END itasegm[443]
  PIN itasegm[444]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1338.400 320.000 1338.960 ;
    END
  END itasegm[444]
  PIN itasegm[445]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1341.200 320.000 1341.760 ;
    END
  END itasegm[445]
  PIN itasegm[446]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1344.000 320.000 1344.560 ;
    END
  END itasegm[446]
  PIN itasegm[447]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1346.800 320.000 1347.360 ;
    END
  END itasegm[447]
  PIN itasegm[448]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1484.000 4.000 1484.560 ;
    END
  END itasegm[448]
  PIN itasegm[449]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1486.800 4.000 1487.360 ;
    END
  END itasegm[449]
  PIN itasegm[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 442.400 4.000 442.960 ;
    END
  END itasegm[44]
  PIN itasegm[450]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1489.600 4.000 1490.160 ;
    END
  END itasegm[450]
  PIN itasegm[451]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1492.400 4.000 1492.960 ;
    END
  END itasegm[451]
  PIN itasegm[452]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1495.200 4.000 1495.760 ;
    END
  END itasegm[452]
  PIN itasegm[453]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1498.000 4.000 1498.560 ;
    END
  END itasegm[453]
  PIN itasegm[454]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1500.800 4.000 1501.360 ;
    END
  END itasegm[454]
  PIN itasegm[455]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1503.600 4.000 1504.160 ;
    END
  END itasegm[455]
  PIN itasegm[456]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1506.400 4.000 1506.960 ;
    END
  END itasegm[456]
  PIN itasegm[457]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1509.200 4.000 1509.760 ;
    END
  END itasegm[457]
  PIN itasegm[458]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1512.000 4.000 1512.560 ;
    END
  END itasegm[458]
  PIN itasegm[459]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1514.800 4.000 1515.360 ;
    END
  END itasegm[459]
  PIN itasegm[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 445.200 4.000 445.760 ;
    END
  END itasegm[45]
  PIN itasegm[460]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1517.600 4.000 1518.160 ;
    END
  END itasegm[460]
  PIN itasegm[461]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1520.400 4.000 1520.960 ;
    END
  END itasegm[461]
  PIN itasegm[462]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1523.200 4.000 1523.760 ;
    END
  END itasegm[462]
  PIN itasegm[463]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1526.000 4.000 1526.560 ;
    END
  END itasegm[463]
  PIN itasegm[464]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1528.800 4.000 1529.360 ;
    END
  END itasegm[464]
  PIN itasegm[465]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1531.600 4.000 1532.160 ;
    END
  END itasegm[465]
  PIN itasegm[466]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1534.400 4.000 1534.960 ;
    END
  END itasegm[466]
  PIN itasegm[467]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1537.200 4.000 1537.760 ;
    END
  END itasegm[467]
  PIN itasegm[468]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1540.000 4.000 1540.560 ;
    END
  END itasegm[468]
  PIN itasegm[469]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1542.800 4.000 1543.360 ;
    END
  END itasegm[469]
  PIN itasegm[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 448.000 4.000 448.560 ;
    END
  END itasegm[46]
  PIN itasegm[470]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1545.600 4.000 1546.160 ;
    END
  END itasegm[470]
  PIN itasegm[471]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1548.400 4.000 1548.960 ;
    END
  END itasegm[471]
  PIN itasegm[472]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1551.200 4.000 1551.760 ;
    END
  END itasegm[472]
  PIN itasegm[473]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1554.000 4.000 1554.560 ;
    END
  END itasegm[473]
  PIN itasegm[474]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1556.800 4.000 1557.360 ;
    END
  END itasegm[474]
  PIN itasegm[475]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1559.600 4.000 1560.160 ;
    END
  END itasegm[475]
  PIN itasegm[476]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1562.400 4.000 1562.960 ;
    END
  END itasegm[476]
  PIN itasegm[477]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1565.200 4.000 1565.760 ;
    END
  END itasegm[477]
  PIN itasegm[478]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1568.000 4.000 1568.560 ;
    END
  END itasegm[478]
  PIN itasegm[479]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1570.800 4.000 1571.360 ;
    END
  END itasegm[479]
  PIN itasegm[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 450.800 4.000 451.360 ;
    END
  END itasegm[47]
  PIN itasegm[480]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1573.600 4.000 1574.160 ;
    END
  END itasegm[480]
  PIN itasegm[481]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1576.400 4.000 1576.960 ;
    END
  END itasegm[481]
  PIN itasegm[482]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1579.200 4.000 1579.760 ;
    END
  END itasegm[482]
  PIN itasegm[483]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1582.000 4.000 1582.560 ;
    END
  END itasegm[483]
  PIN itasegm[484]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1584.800 4.000 1585.360 ;
    END
  END itasegm[484]
  PIN itasegm[485]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1587.600 4.000 1588.160 ;
    END
  END itasegm[485]
  PIN itasegm[486]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1590.400 4.000 1590.960 ;
    END
  END itasegm[486]
  PIN itasegm[487]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1593.200 4.000 1593.760 ;
    END
  END itasegm[487]
  PIN itasegm[488]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1596.000 4.000 1596.560 ;
    END
  END itasegm[488]
  PIN itasegm[489]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1598.800 4.000 1599.360 ;
    END
  END itasegm[489]
  PIN itasegm[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 453.600 4.000 454.160 ;
    END
  END itasegm[48]
  PIN itasegm[490]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1601.600 4.000 1602.160 ;
    END
  END itasegm[490]
  PIN itasegm[491]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1604.400 4.000 1604.960 ;
    END
  END itasegm[491]
  PIN itasegm[492]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1607.200 4.000 1607.760 ;
    END
  END itasegm[492]
  PIN itasegm[493]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1610.000 4.000 1610.560 ;
    END
  END itasegm[493]
  PIN itasegm[494]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1612.800 4.000 1613.360 ;
    END
  END itasegm[494]
  PIN itasegm[495]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1615.600 4.000 1616.160 ;
    END
  END itasegm[495]
  PIN itasegm[496]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1618.400 4.000 1618.960 ;
    END
  END itasegm[496]
  PIN itasegm[497]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1621.200 4.000 1621.760 ;
    END
  END itasegm[497]
  PIN itasegm[498]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1624.000 4.000 1624.560 ;
    END
  END itasegm[498]
  PIN itasegm[499]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1626.800 4.000 1627.360 ;
    END
  END itasegm[499]
  PIN itasegm[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 456.400 4.000 456.960 ;
    END
  END itasegm[49]
  PIN itasegm[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 330.400 4.000 330.960 ;
    END
  END itasegm[4]
  PIN itasegm[500]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1629.600 4.000 1630.160 ;
    END
  END itasegm[500]
  PIN itasegm[501]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1632.400 4.000 1632.960 ;
    END
  END itasegm[501]
  PIN itasegm[502]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1635.200 4.000 1635.760 ;
    END
  END itasegm[502]
  PIN itasegm[503]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1638.000 4.000 1638.560 ;
    END
  END itasegm[503]
  PIN itasegm[504]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1484.000 320.000 1484.560 ;
    END
  END itasegm[504]
  PIN itasegm[505]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1486.800 320.000 1487.360 ;
    END
  END itasegm[505]
  PIN itasegm[506]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1489.600 320.000 1490.160 ;
    END
  END itasegm[506]
  PIN itasegm[507]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1492.400 320.000 1492.960 ;
    END
  END itasegm[507]
  PIN itasegm[508]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1495.200 320.000 1495.760 ;
    END
  END itasegm[508]
  PIN itasegm[509]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1498.000 320.000 1498.560 ;
    END
  END itasegm[509]
  PIN itasegm[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 459.200 4.000 459.760 ;
    END
  END itasegm[50]
  PIN itasegm[510]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1500.800 320.000 1501.360 ;
    END
  END itasegm[510]
  PIN itasegm[511]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1503.600 320.000 1504.160 ;
    END
  END itasegm[511]
  PIN itasegm[512]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1506.400 320.000 1506.960 ;
    END
  END itasegm[512]
  PIN itasegm[513]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1509.200 320.000 1509.760 ;
    END
  END itasegm[513]
  PIN itasegm[514]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1512.000 320.000 1512.560 ;
    END
  END itasegm[514]
  PIN itasegm[515]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1514.800 320.000 1515.360 ;
    END
  END itasegm[515]
  PIN itasegm[516]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1517.600 320.000 1518.160 ;
    END
  END itasegm[516]
  PIN itasegm[517]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1520.400 320.000 1520.960 ;
    END
  END itasegm[517]
  PIN itasegm[518]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1523.200 320.000 1523.760 ;
    END
  END itasegm[518]
  PIN itasegm[519]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1526.000 320.000 1526.560 ;
    END
  END itasegm[519]
  PIN itasegm[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 462.000 4.000 462.560 ;
    END
  END itasegm[51]
  PIN itasegm[520]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1528.800 320.000 1529.360 ;
    END
  END itasegm[520]
  PIN itasegm[521]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1531.600 320.000 1532.160 ;
    END
  END itasegm[521]
  PIN itasegm[522]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1534.400 320.000 1534.960 ;
    END
  END itasegm[522]
  PIN itasegm[523]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1537.200 320.000 1537.760 ;
    END
  END itasegm[523]
  PIN itasegm[524]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1540.000 320.000 1540.560 ;
    END
  END itasegm[524]
  PIN itasegm[525]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1542.800 320.000 1543.360 ;
    END
  END itasegm[525]
  PIN itasegm[526]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1545.600 320.000 1546.160 ;
    END
  END itasegm[526]
  PIN itasegm[527]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1548.400 320.000 1548.960 ;
    END
  END itasegm[527]
  PIN itasegm[528]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1551.200 320.000 1551.760 ;
    END
  END itasegm[528]
  PIN itasegm[529]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1554.000 320.000 1554.560 ;
    END
  END itasegm[529]
  PIN itasegm[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 464.800 4.000 465.360 ;
    END
  END itasegm[52]
  PIN itasegm[530]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1556.800 320.000 1557.360 ;
    END
  END itasegm[530]
  PIN itasegm[531]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1559.600 320.000 1560.160 ;
    END
  END itasegm[531]
  PIN itasegm[532]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1562.400 320.000 1562.960 ;
    END
  END itasegm[532]
  PIN itasegm[533]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1565.200 320.000 1565.760 ;
    END
  END itasegm[533]
  PIN itasegm[534]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1568.000 320.000 1568.560 ;
    END
  END itasegm[534]
  PIN itasegm[535]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1570.800 320.000 1571.360 ;
    END
  END itasegm[535]
  PIN itasegm[536]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1573.600 320.000 1574.160 ;
    END
  END itasegm[536]
  PIN itasegm[537]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1576.400 320.000 1576.960 ;
    END
  END itasegm[537]
  PIN itasegm[538]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1579.200 320.000 1579.760 ;
    END
  END itasegm[538]
  PIN itasegm[539]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1582.000 320.000 1582.560 ;
    END
  END itasegm[539]
  PIN itasegm[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 467.600 4.000 468.160 ;
    END
  END itasegm[53]
  PIN itasegm[540]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1584.800 320.000 1585.360 ;
    END
  END itasegm[540]
  PIN itasegm[541]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1587.600 320.000 1588.160 ;
    END
  END itasegm[541]
  PIN itasegm[542]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1590.400 320.000 1590.960 ;
    END
  END itasegm[542]
  PIN itasegm[543]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1593.200 320.000 1593.760 ;
    END
  END itasegm[543]
  PIN itasegm[544]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1596.000 320.000 1596.560 ;
    END
  END itasegm[544]
  PIN itasegm[545]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1598.800 320.000 1599.360 ;
    END
  END itasegm[545]
  PIN itasegm[546]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1601.600 320.000 1602.160 ;
    END
  END itasegm[546]
  PIN itasegm[547]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1604.400 320.000 1604.960 ;
    END
  END itasegm[547]
  PIN itasegm[548]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1607.200 320.000 1607.760 ;
    END
  END itasegm[548]
  PIN itasegm[549]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1610.000 320.000 1610.560 ;
    END
  END itasegm[549]
  PIN itasegm[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 470.400 4.000 470.960 ;
    END
  END itasegm[54]
  PIN itasegm[550]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1612.800 320.000 1613.360 ;
    END
  END itasegm[550]
  PIN itasegm[551]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1615.600 320.000 1616.160 ;
    END
  END itasegm[551]
  PIN itasegm[552]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1618.400 320.000 1618.960 ;
    END
  END itasegm[552]
  PIN itasegm[553]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1621.200 320.000 1621.760 ;
    END
  END itasegm[553]
  PIN itasegm[554]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1624.000 320.000 1624.560 ;
    END
  END itasegm[554]
  PIN itasegm[555]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1626.800 320.000 1627.360 ;
    END
  END itasegm[555]
  PIN itasegm[556]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1629.600 320.000 1630.160 ;
    END
  END itasegm[556]
  PIN itasegm[557]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1632.400 320.000 1632.960 ;
    END
  END itasegm[557]
  PIN itasegm[558]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1635.200 320.000 1635.760 ;
    END
  END itasegm[558]
  PIN itasegm[559]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1638.000 320.000 1638.560 ;
    END
  END itasegm[559]
  PIN itasegm[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 473.200 4.000 473.760 ;
    END
  END itasegm[55]
  PIN itasegm[560]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1775.200 4.000 1775.760 ;
    END
  END itasegm[560]
  PIN itasegm[561]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1778.000 4.000 1778.560 ;
    END
  END itasegm[561]
  PIN itasegm[562]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1780.800 4.000 1781.360 ;
    END
  END itasegm[562]
  PIN itasegm[563]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1783.600 4.000 1784.160 ;
    END
  END itasegm[563]
  PIN itasegm[564]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1786.400 4.000 1786.960 ;
    END
  END itasegm[564]
  PIN itasegm[565]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1789.200 4.000 1789.760 ;
    END
  END itasegm[565]
  PIN itasegm[566]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1792.000 4.000 1792.560 ;
    END
  END itasegm[566]
  PIN itasegm[567]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1794.800 4.000 1795.360 ;
    END
  END itasegm[567]
  PIN itasegm[568]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1797.600 4.000 1798.160 ;
    END
  END itasegm[568]
  PIN itasegm[569]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1800.400 4.000 1800.960 ;
    END
  END itasegm[569]
  PIN itasegm[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 319.200 320.000 319.760 ;
    END
  END itasegm[56]
  PIN itasegm[570]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1803.200 4.000 1803.760 ;
    END
  END itasegm[570]
  PIN itasegm[571]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1806.000 4.000 1806.560 ;
    END
  END itasegm[571]
  PIN itasegm[572]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1808.800 4.000 1809.360 ;
    END
  END itasegm[572]
  PIN itasegm[573]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1811.600 4.000 1812.160 ;
    END
  END itasegm[573]
  PIN itasegm[574]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1814.400 4.000 1814.960 ;
    END
  END itasegm[574]
  PIN itasegm[575]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1817.200 4.000 1817.760 ;
    END
  END itasegm[575]
  PIN itasegm[576]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1820.000 4.000 1820.560 ;
    END
  END itasegm[576]
  PIN itasegm[577]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1822.800 4.000 1823.360 ;
    END
  END itasegm[577]
  PIN itasegm[578]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1825.600 4.000 1826.160 ;
    END
  END itasegm[578]
  PIN itasegm[579]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1828.400 4.000 1828.960 ;
    END
  END itasegm[579]
  PIN itasegm[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 322.000 320.000 322.560 ;
    END
  END itasegm[57]
  PIN itasegm[580]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1831.200 4.000 1831.760 ;
    END
  END itasegm[580]
  PIN itasegm[581]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1834.000 4.000 1834.560 ;
    END
  END itasegm[581]
  PIN itasegm[582]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1836.800 4.000 1837.360 ;
    END
  END itasegm[582]
  PIN itasegm[583]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1839.600 4.000 1840.160 ;
    END
  END itasegm[583]
  PIN itasegm[584]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1842.400 4.000 1842.960 ;
    END
  END itasegm[584]
  PIN itasegm[585]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1845.200 4.000 1845.760 ;
    END
  END itasegm[585]
  PIN itasegm[586]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1848.000 4.000 1848.560 ;
    END
  END itasegm[586]
  PIN itasegm[587]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1850.800 4.000 1851.360 ;
    END
  END itasegm[587]
  PIN itasegm[588]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1853.600 4.000 1854.160 ;
    END
  END itasegm[588]
  PIN itasegm[589]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1856.400 4.000 1856.960 ;
    END
  END itasegm[589]
  PIN itasegm[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 324.800 320.000 325.360 ;
    END
  END itasegm[58]
  PIN itasegm[590]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1859.200 4.000 1859.760 ;
    END
  END itasegm[590]
  PIN itasegm[591]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1862.000 4.000 1862.560 ;
    END
  END itasegm[591]
  PIN itasegm[592]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1864.800 4.000 1865.360 ;
    END
  END itasegm[592]
  PIN itasegm[593]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1867.600 4.000 1868.160 ;
    END
  END itasegm[593]
  PIN itasegm[594]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1870.400 4.000 1870.960 ;
    END
  END itasegm[594]
  PIN itasegm[595]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1873.200 4.000 1873.760 ;
    END
  END itasegm[595]
  PIN itasegm[596]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1876.000 4.000 1876.560 ;
    END
  END itasegm[596]
  PIN itasegm[597]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1878.800 4.000 1879.360 ;
    END
  END itasegm[597]
  PIN itasegm[598]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1881.600 4.000 1882.160 ;
    END
  END itasegm[598]
  PIN itasegm[599]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1884.400 4.000 1884.960 ;
    END
  END itasegm[599]
  PIN itasegm[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 327.600 320.000 328.160 ;
    END
  END itasegm[59]
  PIN itasegm[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 333.200 4.000 333.760 ;
    END
  END itasegm[5]
  PIN itasegm[600]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1887.200 4.000 1887.760 ;
    END
  END itasegm[600]
  PIN itasegm[601]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1890.000 4.000 1890.560 ;
    END
  END itasegm[601]
  PIN itasegm[602]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1892.800 4.000 1893.360 ;
    END
  END itasegm[602]
  PIN itasegm[603]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1895.600 4.000 1896.160 ;
    END
  END itasegm[603]
  PIN itasegm[604]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1898.400 4.000 1898.960 ;
    END
  END itasegm[604]
  PIN itasegm[605]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1901.200 4.000 1901.760 ;
    END
  END itasegm[605]
  PIN itasegm[606]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1904.000 4.000 1904.560 ;
    END
  END itasegm[606]
  PIN itasegm[607]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1906.800 4.000 1907.360 ;
    END
  END itasegm[607]
  PIN itasegm[608]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1909.600 4.000 1910.160 ;
    END
  END itasegm[608]
  PIN itasegm[609]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1912.400 4.000 1912.960 ;
    END
  END itasegm[609]
  PIN itasegm[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 330.400 320.000 330.960 ;
    END
  END itasegm[60]
  PIN itasegm[610]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1915.200 4.000 1915.760 ;
    END
  END itasegm[610]
  PIN itasegm[611]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1918.000 4.000 1918.560 ;
    END
  END itasegm[611]
  PIN itasegm[612]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1920.800 4.000 1921.360 ;
    END
  END itasegm[612]
  PIN itasegm[613]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1923.600 4.000 1924.160 ;
    END
  END itasegm[613]
  PIN itasegm[614]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1926.400 4.000 1926.960 ;
    END
  END itasegm[614]
  PIN itasegm[615]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1929.200 4.000 1929.760 ;
    END
  END itasegm[615]
  PIN itasegm[616]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1775.200 320.000 1775.760 ;
    END
  END itasegm[616]
  PIN itasegm[617]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1778.000 320.000 1778.560 ;
    END
  END itasegm[617]
  PIN itasegm[618]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1780.800 320.000 1781.360 ;
    END
  END itasegm[618]
  PIN itasegm[619]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1783.600 320.000 1784.160 ;
    END
  END itasegm[619]
  PIN itasegm[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 333.200 320.000 333.760 ;
    END
  END itasegm[61]
  PIN itasegm[620]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1786.400 320.000 1786.960 ;
    END
  END itasegm[620]
  PIN itasegm[621]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1789.200 320.000 1789.760 ;
    END
  END itasegm[621]
  PIN itasegm[622]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1792.000 320.000 1792.560 ;
    END
  END itasegm[622]
  PIN itasegm[623]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1794.800 320.000 1795.360 ;
    END
  END itasegm[623]
  PIN itasegm[624]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1797.600 320.000 1798.160 ;
    END
  END itasegm[624]
  PIN itasegm[625]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1800.400 320.000 1800.960 ;
    END
  END itasegm[625]
  PIN itasegm[626]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1803.200 320.000 1803.760 ;
    END
  END itasegm[626]
  PIN itasegm[627]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1806.000 320.000 1806.560 ;
    END
  END itasegm[627]
  PIN itasegm[628]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1808.800 320.000 1809.360 ;
    END
  END itasegm[628]
  PIN itasegm[629]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1811.600 320.000 1812.160 ;
    END
  END itasegm[629]
  PIN itasegm[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 336.000 320.000 336.560 ;
    END
  END itasegm[62]
  PIN itasegm[630]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1814.400 320.000 1814.960 ;
    END
  END itasegm[630]
  PIN itasegm[631]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1817.200 320.000 1817.760 ;
    END
  END itasegm[631]
  PIN itasegm[632]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1820.000 320.000 1820.560 ;
    END
  END itasegm[632]
  PIN itasegm[633]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1822.800 320.000 1823.360 ;
    END
  END itasegm[633]
  PIN itasegm[634]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1825.600 320.000 1826.160 ;
    END
  END itasegm[634]
  PIN itasegm[635]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1828.400 320.000 1828.960 ;
    END
  END itasegm[635]
  PIN itasegm[636]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1831.200 320.000 1831.760 ;
    END
  END itasegm[636]
  PIN itasegm[637]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1834.000 320.000 1834.560 ;
    END
  END itasegm[637]
  PIN itasegm[638]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1836.800 320.000 1837.360 ;
    END
  END itasegm[638]
  PIN itasegm[639]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1839.600 320.000 1840.160 ;
    END
  END itasegm[639]
  PIN itasegm[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 338.800 320.000 339.360 ;
    END
  END itasegm[63]
  PIN itasegm[640]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1842.400 320.000 1842.960 ;
    END
  END itasegm[640]
  PIN itasegm[641]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1845.200 320.000 1845.760 ;
    END
  END itasegm[641]
  PIN itasegm[642]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1848.000 320.000 1848.560 ;
    END
  END itasegm[642]
  PIN itasegm[643]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1850.800 320.000 1851.360 ;
    END
  END itasegm[643]
  PIN itasegm[644]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1853.600 320.000 1854.160 ;
    END
  END itasegm[644]
  PIN itasegm[645]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1856.400 320.000 1856.960 ;
    END
  END itasegm[645]
  PIN itasegm[646]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1859.200 320.000 1859.760 ;
    END
  END itasegm[646]
  PIN itasegm[647]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1862.000 320.000 1862.560 ;
    END
  END itasegm[647]
  PIN itasegm[648]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1864.800 320.000 1865.360 ;
    END
  END itasegm[648]
  PIN itasegm[649]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1867.600 320.000 1868.160 ;
    END
  END itasegm[649]
  PIN itasegm[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 341.600 320.000 342.160 ;
    END
  END itasegm[64]
  PIN itasegm[650]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1870.400 320.000 1870.960 ;
    END
  END itasegm[650]
  PIN itasegm[651]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1873.200 320.000 1873.760 ;
    END
  END itasegm[651]
  PIN itasegm[652]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1876.000 320.000 1876.560 ;
    END
  END itasegm[652]
  PIN itasegm[653]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1878.800 320.000 1879.360 ;
    END
  END itasegm[653]
  PIN itasegm[654]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1881.600 320.000 1882.160 ;
    END
  END itasegm[654]
  PIN itasegm[655]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1884.400 320.000 1884.960 ;
    END
  END itasegm[655]
  PIN itasegm[656]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1887.200 320.000 1887.760 ;
    END
  END itasegm[656]
  PIN itasegm[657]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1890.000 320.000 1890.560 ;
    END
  END itasegm[657]
  PIN itasegm[658]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1892.800 320.000 1893.360 ;
    END
  END itasegm[658]
  PIN itasegm[659]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1895.600 320.000 1896.160 ;
    END
  END itasegm[659]
  PIN itasegm[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 344.400 320.000 344.960 ;
    END
  END itasegm[65]
  PIN itasegm[660]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1898.400 320.000 1898.960 ;
    END
  END itasegm[660]
  PIN itasegm[661]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1901.200 320.000 1901.760 ;
    END
  END itasegm[661]
  PIN itasegm[662]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1904.000 320.000 1904.560 ;
    END
  END itasegm[662]
  PIN itasegm[663]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1906.800 320.000 1907.360 ;
    END
  END itasegm[663]
  PIN itasegm[664]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1909.600 320.000 1910.160 ;
    END
  END itasegm[664]
  PIN itasegm[665]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1912.400 320.000 1912.960 ;
    END
  END itasegm[665]
  PIN itasegm[666]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1915.200 320.000 1915.760 ;
    END
  END itasegm[666]
  PIN itasegm[667]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1918.000 320.000 1918.560 ;
    END
  END itasegm[667]
  PIN itasegm[668]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1920.800 320.000 1921.360 ;
    END
  END itasegm[668]
  PIN itasegm[669]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1923.600 320.000 1924.160 ;
    END
  END itasegm[669]
  PIN itasegm[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 347.200 320.000 347.760 ;
    END
  END itasegm[66]
  PIN itasegm[670]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1926.400 320.000 1926.960 ;
    END
  END itasegm[670]
  PIN itasegm[671]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1929.200 320.000 1929.760 ;
    END
  END itasegm[671]
  PIN itasegm[672]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2066.400 4.000 2066.960 ;
    END
  END itasegm[672]
  PIN itasegm[673]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2069.200 4.000 2069.760 ;
    END
  END itasegm[673]
  PIN itasegm[674]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2072.000 4.000 2072.560 ;
    END
  END itasegm[674]
  PIN itasegm[675]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2074.800 4.000 2075.360 ;
    END
  END itasegm[675]
  PIN itasegm[676]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2077.600 4.000 2078.160 ;
    END
  END itasegm[676]
  PIN itasegm[677]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2080.400 4.000 2080.960 ;
    END
  END itasegm[677]
  PIN itasegm[678]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2083.200 4.000 2083.760 ;
    END
  END itasegm[678]
  PIN itasegm[679]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2086.000 4.000 2086.560 ;
    END
  END itasegm[679]
  PIN itasegm[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 350.000 320.000 350.560 ;
    END
  END itasegm[67]
  PIN itasegm[680]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2088.800 4.000 2089.360 ;
    END
  END itasegm[680]
  PIN itasegm[681]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2091.600 4.000 2092.160 ;
    END
  END itasegm[681]
  PIN itasegm[682]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2094.400 4.000 2094.960 ;
    END
  END itasegm[682]
  PIN itasegm[683]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2097.200 4.000 2097.760 ;
    END
  END itasegm[683]
  PIN itasegm[684]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2100.000 4.000 2100.560 ;
    END
  END itasegm[684]
  PIN itasegm[685]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2102.800 4.000 2103.360 ;
    END
  END itasegm[685]
  PIN itasegm[686]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2105.600 4.000 2106.160 ;
    END
  END itasegm[686]
  PIN itasegm[687]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2108.400 4.000 2108.960 ;
    END
  END itasegm[687]
  PIN itasegm[688]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2111.200 4.000 2111.760 ;
    END
  END itasegm[688]
  PIN itasegm[689]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2114.000 4.000 2114.560 ;
    END
  END itasegm[689]
  PIN itasegm[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 352.800 320.000 353.360 ;
    END
  END itasegm[68]
  PIN itasegm[690]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2116.800 4.000 2117.360 ;
    END
  END itasegm[690]
  PIN itasegm[691]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2119.600 4.000 2120.160 ;
    END
  END itasegm[691]
  PIN itasegm[692]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2122.400 4.000 2122.960 ;
    END
  END itasegm[692]
  PIN itasegm[693]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2125.200 4.000 2125.760 ;
    END
  END itasegm[693]
  PIN itasegm[694]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2128.000 4.000 2128.560 ;
    END
  END itasegm[694]
  PIN itasegm[695]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2130.800 4.000 2131.360 ;
    END
  END itasegm[695]
  PIN itasegm[696]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2133.600 4.000 2134.160 ;
    END
  END itasegm[696]
  PIN itasegm[697]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2136.400 4.000 2136.960 ;
    END
  END itasegm[697]
  PIN itasegm[698]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2139.200 4.000 2139.760 ;
    END
  END itasegm[698]
  PIN itasegm[699]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2142.000 4.000 2142.560 ;
    END
  END itasegm[699]
  PIN itasegm[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 355.600 320.000 356.160 ;
    END
  END itasegm[69]
  PIN itasegm[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 336.000 4.000 336.560 ;
    END
  END itasegm[6]
  PIN itasegm[700]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2144.800 4.000 2145.360 ;
    END
  END itasegm[700]
  PIN itasegm[701]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2147.600 4.000 2148.160 ;
    END
  END itasegm[701]
  PIN itasegm[702]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2150.400 4.000 2150.960 ;
    END
  END itasegm[702]
  PIN itasegm[703]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2153.200 4.000 2153.760 ;
    END
  END itasegm[703]
  PIN itasegm[704]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2156.000 4.000 2156.560 ;
    END
  END itasegm[704]
  PIN itasegm[705]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2158.800 4.000 2159.360 ;
    END
  END itasegm[705]
  PIN itasegm[706]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2161.600 4.000 2162.160 ;
    END
  END itasegm[706]
  PIN itasegm[707]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2164.400 4.000 2164.960 ;
    END
  END itasegm[707]
  PIN itasegm[708]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2167.200 4.000 2167.760 ;
    END
  END itasegm[708]
  PIN itasegm[709]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2170.000 4.000 2170.560 ;
    END
  END itasegm[709]
  PIN itasegm[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 358.400 320.000 358.960 ;
    END
  END itasegm[70]
  PIN itasegm[710]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2172.800 4.000 2173.360 ;
    END
  END itasegm[710]
  PIN itasegm[711]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2175.600 4.000 2176.160 ;
    END
  END itasegm[711]
  PIN itasegm[712]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2178.400 4.000 2178.960 ;
    END
  END itasegm[712]
  PIN itasegm[713]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2181.200 4.000 2181.760 ;
    END
  END itasegm[713]
  PIN itasegm[714]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2184.000 4.000 2184.560 ;
    END
  END itasegm[714]
  PIN itasegm[715]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2186.800 4.000 2187.360 ;
    END
  END itasegm[715]
  PIN itasegm[716]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2189.600 4.000 2190.160 ;
    END
  END itasegm[716]
  PIN itasegm[717]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2192.400 4.000 2192.960 ;
    END
  END itasegm[717]
  PIN itasegm[718]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2195.200 4.000 2195.760 ;
    END
  END itasegm[718]
  PIN itasegm[719]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2198.000 4.000 2198.560 ;
    END
  END itasegm[719]
  PIN itasegm[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 361.200 320.000 361.760 ;
    END
  END itasegm[71]
  PIN itasegm[720]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2200.800 4.000 2201.360 ;
    END
  END itasegm[720]
  PIN itasegm[721]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2203.600 4.000 2204.160 ;
    END
  END itasegm[721]
  PIN itasegm[722]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2206.400 4.000 2206.960 ;
    END
  END itasegm[722]
  PIN itasegm[723]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2209.200 4.000 2209.760 ;
    END
  END itasegm[723]
  PIN itasegm[724]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2212.000 4.000 2212.560 ;
    END
  END itasegm[724]
  PIN itasegm[725]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2214.800 4.000 2215.360 ;
    END
  END itasegm[725]
  PIN itasegm[726]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2217.600 4.000 2218.160 ;
    END
  END itasegm[726]
  PIN itasegm[727]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2220.400 4.000 2220.960 ;
    END
  END itasegm[727]
  PIN itasegm[728]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2066.400 320.000 2066.960 ;
    END
  END itasegm[728]
  PIN itasegm[729]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2069.200 320.000 2069.760 ;
    END
  END itasegm[729]
  PIN itasegm[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 364.000 320.000 364.560 ;
    END
  END itasegm[72]
  PIN itasegm[730]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2072.000 320.000 2072.560 ;
    END
  END itasegm[730]
  PIN itasegm[731]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2074.800 320.000 2075.360 ;
    END
  END itasegm[731]
  PIN itasegm[732]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2077.600 320.000 2078.160 ;
    END
  END itasegm[732]
  PIN itasegm[733]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2080.400 320.000 2080.960 ;
    END
  END itasegm[733]
  PIN itasegm[734]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2083.200 320.000 2083.760 ;
    END
  END itasegm[734]
  PIN itasegm[735]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2086.000 320.000 2086.560 ;
    END
  END itasegm[735]
  PIN itasegm[736]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2088.800 320.000 2089.360 ;
    END
  END itasegm[736]
  PIN itasegm[737]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2091.600 320.000 2092.160 ;
    END
  END itasegm[737]
  PIN itasegm[738]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2094.400 320.000 2094.960 ;
    END
  END itasegm[738]
  PIN itasegm[739]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2097.200 320.000 2097.760 ;
    END
  END itasegm[739]
  PIN itasegm[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 366.800 320.000 367.360 ;
    END
  END itasegm[73]
  PIN itasegm[740]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2100.000 320.000 2100.560 ;
    END
  END itasegm[740]
  PIN itasegm[741]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2102.800 320.000 2103.360 ;
    END
  END itasegm[741]
  PIN itasegm[742]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2105.600 320.000 2106.160 ;
    END
  END itasegm[742]
  PIN itasegm[743]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2108.400 320.000 2108.960 ;
    END
  END itasegm[743]
  PIN itasegm[744]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2111.200 320.000 2111.760 ;
    END
  END itasegm[744]
  PIN itasegm[745]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2114.000 320.000 2114.560 ;
    END
  END itasegm[745]
  PIN itasegm[746]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2116.800 320.000 2117.360 ;
    END
  END itasegm[746]
  PIN itasegm[747]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2119.600 320.000 2120.160 ;
    END
  END itasegm[747]
  PIN itasegm[748]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2122.400 320.000 2122.960 ;
    END
  END itasegm[748]
  PIN itasegm[749]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2125.200 320.000 2125.760 ;
    END
  END itasegm[749]
  PIN itasegm[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 369.600 320.000 370.160 ;
    END
  END itasegm[74]
  PIN itasegm[750]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2128.000 320.000 2128.560 ;
    END
  END itasegm[750]
  PIN itasegm[751]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2130.800 320.000 2131.360 ;
    END
  END itasegm[751]
  PIN itasegm[752]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2133.600 320.000 2134.160 ;
    END
  END itasegm[752]
  PIN itasegm[753]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2136.400 320.000 2136.960 ;
    END
  END itasegm[753]
  PIN itasegm[754]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2139.200 320.000 2139.760 ;
    END
  END itasegm[754]
  PIN itasegm[755]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2142.000 320.000 2142.560 ;
    END
  END itasegm[755]
  PIN itasegm[756]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2144.800 320.000 2145.360 ;
    END
  END itasegm[756]
  PIN itasegm[757]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2147.600 320.000 2148.160 ;
    END
  END itasegm[757]
  PIN itasegm[758]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2150.400 320.000 2150.960 ;
    END
  END itasegm[758]
  PIN itasegm[759]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2153.200 320.000 2153.760 ;
    END
  END itasegm[759]
  PIN itasegm[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 372.400 320.000 372.960 ;
    END
  END itasegm[75]
  PIN itasegm[760]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2156.000 320.000 2156.560 ;
    END
  END itasegm[760]
  PIN itasegm[761]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2158.800 320.000 2159.360 ;
    END
  END itasegm[761]
  PIN itasegm[762]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2161.600 320.000 2162.160 ;
    END
  END itasegm[762]
  PIN itasegm[763]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2164.400 320.000 2164.960 ;
    END
  END itasegm[763]
  PIN itasegm[764]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2167.200 320.000 2167.760 ;
    END
  END itasegm[764]
  PIN itasegm[765]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2170.000 320.000 2170.560 ;
    END
  END itasegm[765]
  PIN itasegm[766]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2172.800 320.000 2173.360 ;
    END
  END itasegm[766]
  PIN itasegm[767]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2175.600 320.000 2176.160 ;
    END
  END itasegm[767]
  PIN itasegm[768]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2178.400 320.000 2178.960 ;
    END
  END itasegm[768]
  PIN itasegm[769]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2181.200 320.000 2181.760 ;
    END
  END itasegm[769]
  PIN itasegm[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 375.200 320.000 375.760 ;
    END
  END itasegm[76]
  PIN itasegm[770]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2184.000 320.000 2184.560 ;
    END
  END itasegm[770]
  PIN itasegm[771]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2186.800 320.000 2187.360 ;
    END
  END itasegm[771]
  PIN itasegm[772]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.408000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2189.600 320.000 2190.160 ;
    END
  END itasegm[772]
  PIN itasegm[773]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.408000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2192.400 320.000 2192.960 ;
    END
  END itasegm[773]
  PIN itasegm[774]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2195.200 320.000 2195.760 ;
    END
  END itasegm[774]
  PIN itasegm[775]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.408000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2198.000 320.000 2198.560 ;
    END
  END itasegm[775]
  PIN itasegm[776]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2200.800 320.000 2201.360 ;
    END
  END itasegm[776]
  PIN itasegm[777]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2203.600 320.000 2204.160 ;
    END
  END itasegm[777]
  PIN itasegm[778]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2206.400 320.000 2206.960 ;
    END
  END itasegm[778]
  PIN itasegm[779]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2209.200 320.000 2209.760 ;
    END
  END itasegm[779]
  PIN itasegm[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 378.000 320.000 378.560 ;
    END
  END itasegm[77]
  PIN itasegm[780]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2212.000 320.000 2212.560 ;
    END
  END itasegm[780]
  PIN itasegm[781]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2214.800 320.000 2215.360 ;
    END
  END itasegm[781]
  PIN itasegm[782]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2217.600 320.000 2218.160 ;
    END
  END itasegm[782]
  PIN itasegm[783]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2220.400 320.000 2220.960 ;
    END
  END itasegm[783]
  PIN itasegm[784]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2357.600 4.000 2358.160 ;
    END
  END itasegm[784]
  PIN itasegm[785]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2360.400 4.000 2360.960 ;
    END
  END itasegm[785]
  PIN itasegm[786]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2363.200 4.000 2363.760 ;
    END
  END itasegm[786]
  PIN itasegm[787]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2366.000 4.000 2366.560 ;
    END
  END itasegm[787]
  PIN itasegm[788]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2368.800 4.000 2369.360 ;
    END
  END itasegm[788]
  PIN itasegm[789]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2371.600 4.000 2372.160 ;
    END
  END itasegm[789]
  PIN itasegm[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 380.800 320.000 381.360 ;
    END
  END itasegm[78]
  PIN itasegm[790]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2374.400 4.000 2374.960 ;
    END
  END itasegm[790]
  PIN itasegm[791]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2377.200 4.000 2377.760 ;
    END
  END itasegm[791]
  PIN itasegm[792]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2380.000 4.000 2380.560 ;
    END
  END itasegm[792]
  PIN itasegm[793]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2382.800 4.000 2383.360 ;
    END
  END itasegm[793]
  PIN itasegm[794]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2385.600 4.000 2386.160 ;
    END
  END itasegm[794]
  PIN itasegm[795]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2388.400 4.000 2388.960 ;
    END
  END itasegm[795]
  PIN itasegm[796]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2391.200 4.000 2391.760 ;
    END
  END itasegm[796]
  PIN itasegm[797]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2394.000 4.000 2394.560 ;
    END
  END itasegm[797]
  PIN itasegm[798]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2396.800 4.000 2397.360 ;
    END
  END itasegm[798]
  PIN itasegm[799]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2399.600 4.000 2400.160 ;
    END
  END itasegm[799]
  PIN itasegm[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 383.600 320.000 384.160 ;
    END
  END itasegm[79]
  PIN itasegm[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 338.800 4.000 339.360 ;
    END
  END itasegm[7]
  PIN itasegm[800]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2402.400 4.000 2402.960 ;
    END
  END itasegm[800]
  PIN itasegm[801]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2405.200 4.000 2405.760 ;
    END
  END itasegm[801]
  PIN itasegm[802]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2408.000 4.000 2408.560 ;
    END
  END itasegm[802]
  PIN itasegm[803]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2410.800 4.000 2411.360 ;
    END
  END itasegm[803]
  PIN itasegm[804]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2413.600 4.000 2414.160 ;
    END
  END itasegm[804]
  PIN itasegm[805]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2416.400 4.000 2416.960 ;
    END
  END itasegm[805]
  PIN itasegm[806]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2419.200 4.000 2419.760 ;
    END
  END itasegm[806]
  PIN itasegm[807]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2422.000 4.000 2422.560 ;
    END
  END itasegm[807]
  PIN itasegm[808]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2424.800 4.000 2425.360 ;
    END
  END itasegm[808]
  PIN itasegm[809]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2427.600 4.000 2428.160 ;
    END
  END itasegm[809]
  PIN itasegm[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 386.400 320.000 386.960 ;
    END
  END itasegm[80]
  PIN itasegm[810]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2430.400 4.000 2430.960 ;
    END
  END itasegm[810]
  PIN itasegm[811]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2433.200 4.000 2433.760 ;
    END
  END itasegm[811]
  PIN itasegm[812]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2436.000 4.000 2436.560 ;
    END
  END itasegm[812]
  PIN itasegm[813]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2438.800 4.000 2439.360 ;
    END
  END itasegm[813]
  PIN itasegm[814]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2441.600 4.000 2442.160 ;
    END
  END itasegm[814]
  PIN itasegm[815]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2444.400 4.000 2444.960 ;
    END
  END itasegm[815]
  PIN itasegm[816]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2447.200 4.000 2447.760 ;
    END
  END itasegm[816]
  PIN itasegm[817]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2450.000 4.000 2450.560 ;
    END
  END itasegm[817]
  PIN itasegm[818]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2452.800 4.000 2453.360 ;
    END
  END itasegm[818]
  PIN itasegm[819]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2455.600 4.000 2456.160 ;
    END
  END itasegm[819]
  PIN itasegm[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 389.200 320.000 389.760 ;
    END
  END itasegm[81]
  PIN itasegm[820]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2458.400 4.000 2458.960 ;
    END
  END itasegm[820]
  PIN itasegm[821]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2461.200 4.000 2461.760 ;
    END
  END itasegm[821]
  PIN itasegm[822]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2464.000 4.000 2464.560 ;
    END
  END itasegm[822]
  PIN itasegm[823]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2466.800 4.000 2467.360 ;
    END
  END itasegm[823]
  PIN itasegm[824]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2469.600 4.000 2470.160 ;
    END
  END itasegm[824]
  PIN itasegm[825]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2472.400 4.000 2472.960 ;
    END
  END itasegm[825]
  PIN itasegm[826]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2475.200 4.000 2475.760 ;
    END
  END itasegm[826]
  PIN itasegm[827]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2478.000 4.000 2478.560 ;
    END
  END itasegm[827]
  PIN itasegm[828]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2480.800 4.000 2481.360 ;
    END
  END itasegm[828]
  PIN itasegm[829]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2483.600 4.000 2484.160 ;
    END
  END itasegm[829]
  PIN itasegm[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 392.000 320.000 392.560 ;
    END
  END itasegm[82]
  PIN itasegm[830]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2486.400 4.000 2486.960 ;
    END
  END itasegm[830]
  PIN itasegm[831]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2489.200 4.000 2489.760 ;
    END
  END itasegm[831]
  PIN itasegm[832]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2492.000 4.000 2492.560 ;
    END
  END itasegm[832]
  PIN itasegm[833]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2494.800 4.000 2495.360 ;
    END
  END itasegm[833]
  PIN itasegm[834]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2497.600 4.000 2498.160 ;
    END
  END itasegm[834]
  PIN itasegm[835]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2500.400 4.000 2500.960 ;
    END
  END itasegm[835]
  PIN itasegm[836]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2503.200 4.000 2503.760 ;
    END
  END itasegm[836]
  PIN itasegm[837]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2506.000 4.000 2506.560 ;
    END
  END itasegm[837]
  PIN itasegm[838]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2508.800 4.000 2509.360 ;
    END
  END itasegm[838]
  PIN itasegm[839]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2511.600 4.000 2512.160 ;
    END
  END itasegm[839]
  PIN itasegm[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 394.800 320.000 395.360 ;
    END
  END itasegm[83]
  PIN itasegm[840]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2357.600 320.000 2358.160 ;
    END
  END itasegm[840]
  PIN itasegm[841]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2360.400 320.000 2360.960 ;
    END
  END itasegm[841]
  PIN itasegm[842]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2363.200 320.000 2363.760 ;
    END
  END itasegm[842]
  PIN itasegm[843]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2366.000 320.000 2366.560 ;
    END
  END itasegm[843]
  PIN itasegm[844]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2368.800 320.000 2369.360 ;
    END
  END itasegm[844]
  PIN itasegm[845]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2371.600 320.000 2372.160 ;
    END
  END itasegm[845]
  PIN itasegm[846]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2374.400 320.000 2374.960 ;
    END
  END itasegm[846]
  PIN itasegm[847]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2377.200 320.000 2377.760 ;
    END
  END itasegm[847]
  PIN itasegm[848]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2380.000 320.000 2380.560 ;
    END
  END itasegm[848]
  PIN itasegm[849]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2382.800 320.000 2383.360 ;
    END
  END itasegm[849]
  PIN itasegm[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 397.600 320.000 398.160 ;
    END
  END itasegm[84]
  PIN itasegm[850]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2385.600 320.000 2386.160 ;
    END
  END itasegm[850]
  PIN itasegm[851]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2388.400 320.000 2388.960 ;
    END
  END itasegm[851]
  PIN itasegm[852]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2391.200 320.000 2391.760 ;
    END
  END itasegm[852]
  PIN itasegm[853]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2394.000 320.000 2394.560 ;
    END
  END itasegm[853]
  PIN itasegm[854]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2396.800 320.000 2397.360 ;
    END
  END itasegm[854]
  PIN itasegm[855]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2399.600 320.000 2400.160 ;
    END
  END itasegm[855]
  PIN itasegm[856]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2402.400 320.000 2402.960 ;
    END
  END itasegm[856]
  PIN itasegm[857]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2405.200 320.000 2405.760 ;
    END
  END itasegm[857]
  PIN itasegm[858]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2408.000 320.000 2408.560 ;
    END
  END itasegm[858]
  PIN itasegm[859]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2410.800 320.000 2411.360 ;
    END
  END itasegm[859]
  PIN itasegm[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 400.400 320.000 400.960 ;
    END
  END itasegm[85]
  PIN itasegm[860]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2413.600 320.000 2414.160 ;
    END
  END itasegm[860]
  PIN itasegm[861]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2416.400 320.000 2416.960 ;
    END
  END itasegm[861]
  PIN itasegm[862]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2419.200 320.000 2419.760 ;
    END
  END itasegm[862]
  PIN itasegm[863]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2422.000 320.000 2422.560 ;
    END
  END itasegm[863]
  PIN itasegm[864]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2424.800 320.000 2425.360 ;
    END
  END itasegm[864]
  PIN itasegm[865]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2427.600 320.000 2428.160 ;
    END
  END itasegm[865]
  PIN itasegm[866]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2430.400 320.000 2430.960 ;
    END
  END itasegm[866]
  PIN itasegm[867]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2433.200 320.000 2433.760 ;
    END
  END itasegm[867]
  PIN itasegm[868]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2436.000 320.000 2436.560 ;
    END
  END itasegm[868]
  PIN itasegm[869]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2438.800 320.000 2439.360 ;
    END
  END itasegm[869]
  PIN itasegm[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 403.200 320.000 403.760 ;
    END
  END itasegm[86]
  PIN itasegm[870]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2441.600 320.000 2442.160 ;
    END
  END itasegm[870]
  PIN itasegm[871]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2444.400 320.000 2444.960 ;
    END
  END itasegm[871]
  PIN itasegm[872]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2447.200 320.000 2447.760 ;
    END
  END itasegm[872]
  PIN itasegm[873]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2450.000 320.000 2450.560 ;
    END
  END itasegm[873]
  PIN itasegm[874]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2452.800 320.000 2453.360 ;
    END
  END itasegm[874]
  PIN itasegm[875]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2455.600 320.000 2456.160 ;
    END
  END itasegm[875]
  PIN itasegm[876]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2458.400 320.000 2458.960 ;
    END
  END itasegm[876]
  PIN itasegm[877]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2461.200 320.000 2461.760 ;
    END
  END itasegm[877]
  PIN itasegm[878]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2464.000 320.000 2464.560 ;
    END
  END itasegm[878]
  PIN itasegm[879]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2466.800 320.000 2467.360 ;
    END
  END itasegm[879]
  PIN itasegm[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 406.000 320.000 406.560 ;
    END
  END itasegm[87]
  PIN itasegm[880]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2469.600 320.000 2470.160 ;
    END
  END itasegm[880]
  PIN itasegm[881]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2472.400 320.000 2472.960 ;
    END
  END itasegm[881]
  PIN itasegm[882]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2475.200 320.000 2475.760 ;
    END
  END itasegm[882]
  PIN itasegm[883]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2478.000 320.000 2478.560 ;
    END
  END itasegm[883]
  PIN itasegm[884]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2480.800 320.000 2481.360 ;
    END
  END itasegm[884]
  PIN itasegm[885]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2483.600 320.000 2484.160 ;
    END
  END itasegm[885]
  PIN itasegm[886]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2486.400 320.000 2486.960 ;
    END
  END itasegm[886]
  PIN itasegm[887]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2489.200 320.000 2489.760 ;
    END
  END itasegm[887]
  PIN itasegm[888]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2492.000 320.000 2492.560 ;
    END
  END itasegm[888]
  PIN itasegm[889]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2494.800 320.000 2495.360 ;
    END
  END itasegm[889]
  PIN itasegm[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 408.800 320.000 409.360 ;
    END
  END itasegm[88]
  PIN itasegm[890]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2497.600 320.000 2498.160 ;
    END
  END itasegm[890]
  PIN itasegm[891]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2500.400 320.000 2500.960 ;
    END
  END itasegm[891]
  PIN itasegm[892]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2503.200 320.000 2503.760 ;
    END
  END itasegm[892]
  PIN itasegm[893]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2506.000 320.000 2506.560 ;
    END
  END itasegm[893]
  PIN itasegm[894]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2508.800 320.000 2509.360 ;
    END
  END itasegm[894]
  PIN itasegm[895]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2511.600 320.000 2512.160 ;
    END
  END itasegm[895]
  PIN itasegm[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 411.600 320.000 412.160 ;
    END
  END itasegm[89]
  PIN itasegm[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 341.600 4.000 342.160 ;
    END
  END itasegm[8]
  PIN itasegm[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 414.400 320.000 414.960 ;
    END
  END itasegm[90]
  PIN itasegm[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 417.200 320.000 417.760 ;
    END
  END itasegm[91]
  PIN itasegm[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 420.000 320.000 420.560 ;
    END
  END itasegm[92]
  PIN itasegm[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 422.800 320.000 423.360 ;
    END
  END itasegm[93]
  PIN itasegm[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 425.600 320.000 426.160 ;
    END
  END itasegm[94]
  PIN itasegm[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 428.400 320.000 428.960 ;
    END
  END itasegm[95]
  PIN itasegm[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 431.200 320.000 431.760 ;
    END
  END itasegm[96]
  PIN itasegm[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 434.000 320.000 434.560 ;
    END
  END itasegm[97]
  PIN itasegm[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 436.800 320.000 437.360 ;
    END
  END itasegm[98]
  PIN itasegm[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 439.600 320.000 440.160 ;
    END
  END itasegm[99]
  PIN itasegm[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 344.400 4.000 344.960 ;
    END
  END itasegm[9]
  PIN itasel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 184.800 4.000 185.360 ;
    END
  END itasel[0]
  PIN itasel[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 487.200 4.000 487.760 ;
    END
  END itasel[100]
  PIN itasel[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 490.000 4.000 490.560 ;
    END
  END itasel[101]
  PIN itasel[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 492.800 4.000 493.360 ;
    END
  END itasel[102]
  PIN itasel[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 495.600 4.000 496.160 ;
    END
  END itasel[103]
  PIN itasel[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 498.400 4.000 498.960 ;
    END
  END itasel[104]
  PIN itasel[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 501.200 4.000 501.760 ;
    END
  END itasel[105]
  PIN itasel[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 504.000 4.000 504.560 ;
    END
  END itasel[106]
  PIN itasel[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 506.800 4.000 507.360 ;
    END
  END itasel[107]
  PIN itasel[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 509.600 4.000 510.160 ;
    END
  END itasel[108]
  PIN itasel[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 512.400 4.000 512.960 ;
    END
  END itasel[109]
  PIN itasel[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 212.800 4.000 213.360 ;
    END
  END itasel[10]
  PIN itasel[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 515.200 4.000 515.760 ;
    END
  END itasel[110]
  PIN itasel[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 518.000 4.000 518.560 ;
    END
  END itasel[111]
  PIN itasel[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 520.800 4.000 521.360 ;
    END
  END itasel[112]
  PIN itasel[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 523.600 4.000 524.160 ;
    END
  END itasel[113]
  PIN itasel[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 526.400 4.000 526.960 ;
    END
  END itasel[114]
  PIN itasel[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 529.200 4.000 529.760 ;
    END
  END itasel[115]
  PIN itasel[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 532.000 4.000 532.560 ;
    END
  END itasel[116]
  PIN itasel[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 534.800 4.000 535.360 ;
    END
  END itasel[117]
  PIN itasel[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 537.600 4.000 538.160 ;
    END
  END itasel[118]
  PIN itasel[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 540.400 4.000 540.960 ;
    END
  END itasel[119]
  PIN itasel[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 215.600 4.000 216.160 ;
    END
  END itasel[11]
  PIN itasel[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 543.200 4.000 543.760 ;
    END
  END itasel[120]
  PIN itasel[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 546.000 4.000 546.560 ;
    END
  END itasel[121]
  PIN itasel[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 548.800 4.000 549.360 ;
    END
  END itasel[122]
  PIN itasel[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 551.600 4.000 552.160 ;
    END
  END itasel[123]
  PIN itasel[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 554.400 4.000 554.960 ;
    END
  END itasel[124]
  PIN itasel[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 557.200 4.000 557.760 ;
    END
  END itasel[125]
  PIN itasel[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 560.000 4.000 560.560 ;
    END
  END itasel[126]
  PIN itasel[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 562.800 4.000 563.360 ;
    END
  END itasel[127]
  PIN itasel[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 565.600 4.000 566.160 ;
    END
  END itasel[128]
  PIN itasel[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 568.400 4.000 568.960 ;
    END
  END itasel[129]
  PIN itasel[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 218.400 4.000 218.960 ;
    END
  END itasel[12]
  PIN itasel[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 571.200 4.000 571.760 ;
    END
  END itasel[130]
  PIN itasel[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 574.000 4.000 574.560 ;
    END
  END itasel[131]
  PIN itasel[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 576.800 4.000 577.360 ;
    END
  END itasel[132]
  PIN itasel[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 579.600 4.000 580.160 ;
    END
  END itasel[133]
  PIN itasel[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 582.400 4.000 582.960 ;
    END
  END itasel[134]
  PIN itasel[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 585.200 4.000 585.760 ;
    END
  END itasel[135]
  PIN itasel[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 588.000 4.000 588.560 ;
    END
  END itasel[136]
  PIN itasel[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 590.800 4.000 591.360 ;
    END
  END itasel[137]
  PIN itasel[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 593.600 4.000 594.160 ;
    END
  END itasel[138]
  PIN itasel[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 596.400 4.000 596.960 ;
    END
  END itasel[139]
  PIN itasel[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 221.200 4.000 221.760 ;
    END
  END itasel[13]
  PIN itasel[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 599.200 4.000 599.760 ;
    END
  END itasel[140]
  PIN itasel[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 602.000 4.000 602.560 ;
    END
  END itasel[141]
  PIN itasel[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 604.800 4.000 605.360 ;
    END
  END itasel[142]
  PIN itasel[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 607.600 4.000 608.160 ;
    END
  END itasel[143]
  PIN itasel[144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 476.000 320.000 476.560 ;
    END
  END itasel[144]
  PIN itasel[145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 478.800 320.000 479.360 ;
    END
  END itasel[145]
  PIN itasel[146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 481.600 320.000 482.160 ;
    END
  END itasel[146]
  PIN itasel[147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 484.400 320.000 484.960 ;
    END
  END itasel[147]
  PIN itasel[148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 487.200 320.000 487.760 ;
    END
  END itasel[148]
  PIN itasel[149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 490.000 320.000 490.560 ;
    END
  END itasel[149]
  PIN itasel[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 224.000 4.000 224.560 ;
    END
  END itasel[14]
  PIN itasel[150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 492.800 320.000 493.360 ;
    END
  END itasel[150]
  PIN itasel[151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 495.600 320.000 496.160 ;
    END
  END itasel[151]
  PIN itasel[152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 498.400 320.000 498.960 ;
    END
  END itasel[152]
  PIN itasel[153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 501.200 320.000 501.760 ;
    END
  END itasel[153]
  PIN itasel[154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 504.000 320.000 504.560 ;
    END
  END itasel[154]
  PIN itasel[155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 506.800 320.000 507.360 ;
    END
  END itasel[155]
  PIN itasel[156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 509.600 320.000 510.160 ;
    END
  END itasel[156]
  PIN itasel[157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 512.400 320.000 512.960 ;
    END
  END itasel[157]
  PIN itasel[158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 515.200 320.000 515.760 ;
    END
  END itasel[158]
  PIN itasel[159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 518.000 320.000 518.560 ;
    END
  END itasel[159]
  PIN itasel[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 226.800 4.000 227.360 ;
    END
  END itasel[15]
  PIN itasel[160]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 520.800 320.000 521.360 ;
    END
  END itasel[160]
  PIN itasel[161]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 523.600 320.000 524.160 ;
    END
  END itasel[161]
  PIN itasel[162]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 526.400 320.000 526.960 ;
    END
  END itasel[162]
  PIN itasel[163]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 529.200 320.000 529.760 ;
    END
  END itasel[163]
  PIN itasel[164]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 532.000 320.000 532.560 ;
    END
  END itasel[164]
  PIN itasel[165]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 534.800 320.000 535.360 ;
    END
  END itasel[165]
  PIN itasel[166]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 537.600 320.000 538.160 ;
    END
  END itasel[166]
  PIN itasel[167]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 540.400 320.000 540.960 ;
    END
  END itasel[167]
  PIN itasel[168]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 543.200 320.000 543.760 ;
    END
  END itasel[168]
  PIN itasel[169]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 546.000 320.000 546.560 ;
    END
  END itasel[169]
  PIN itasel[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 229.600 4.000 230.160 ;
    END
  END itasel[16]
  PIN itasel[170]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 548.800 320.000 549.360 ;
    END
  END itasel[170]
  PIN itasel[171]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 551.600 320.000 552.160 ;
    END
  END itasel[171]
  PIN itasel[172]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 554.400 320.000 554.960 ;
    END
  END itasel[172]
  PIN itasel[173]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 557.200 320.000 557.760 ;
    END
  END itasel[173]
  PIN itasel[174]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 560.000 320.000 560.560 ;
    END
  END itasel[174]
  PIN itasel[175]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 562.800 320.000 563.360 ;
    END
  END itasel[175]
  PIN itasel[176]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 565.600 320.000 566.160 ;
    END
  END itasel[176]
  PIN itasel[177]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 568.400 320.000 568.960 ;
    END
  END itasel[177]
  PIN itasel[178]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 571.200 320.000 571.760 ;
    END
  END itasel[178]
  PIN itasel[179]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 574.000 320.000 574.560 ;
    END
  END itasel[179]
  PIN itasel[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 232.400 4.000 232.960 ;
    END
  END itasel[17]
  PIN itasel[180]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 576.800 320.000 577.360 ;
    END
  END itasel[180]
  PIN itasel[181]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 579.600 320.000 580.160 ;
    END
  END itasel[181]
  PIN itasel[182]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 582.400 320.000 582.960 ;
    END
  END itasel[182]
  PIN itasel[183]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 585.200 320.000 585.760 ;
    END
  END itasel[183]
  PIN itasel[184]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 588.000 320.000 588.560 ;
    END
  END itasel[184]
  PIN itasel[185]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 590.800 320.000 591.360 ;
    END
  END itasel[185]
  PIN itasel[186]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 593.600 320.000 594.160 ;
    END
  END itasel[186]
  PIN itasel[187]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 596.400 320.000 596.960 ;
    END
  END itasel[187]
  PIN itasel[188]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 599.200 320.000 599.760 ;
    END
  END itasel[188]
  PIN itasel[189]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 602.000 320.000 602.560 ;
    END
  END itasel[189]
  PIN itasel[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 235.200 4.000 235.760 ;
    END
  END itasel[18]
  PIN itasel[190]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 604.800 320.000 605.360 ;
    END
  END itasel[190]
  PIN itasel[191]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 607.600 320.000 608.160 ;
    END
  END itasel[191]
  PIN itasel[192]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 767.200 4.000 767.760 ;
    END
  END itasel[192]
  PIN itasel[193]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 770.000 4.000 770.560 ;
    END
  END itasel[193]
  PIN itasel[194]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 772.800 4.000 773.360 ;
    END
  END itasel[194]
  PIN itasel[195]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 775.600 4.000 776.160 ;
    END
  END itasel[195]
  PIN itasel[196]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 778.400 4.000 778.960 ;
    END
  END itasel[196]
  PIN itasel[197]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 781.200 4.000 781.760 ;
    END
  END itasel[197]
  PIN itasel[198]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 784.000 4.000 784.560 ;
    END
  END itasel[198]
  PIN itasel[199]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 786.800 4.000 787.360 ;
    END
  END itasel[199]
  PIN itasel[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 238.000 4.000 238.560 ;
    END
  END itasel[19]
  PIN itasel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 187.600 4.000 188.160 ;
    END
  END itasel[1]
  PIN itasel[200]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 789.600 4.000 790.160 ;
    END
  END itasel[200]
  PIN itasel[201]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 792.400 4.000 792.960 ;
    END
  END itasel[201]
  PIN itasel[202]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 795.200 4.000 795.760 ;
    END
  END itasel[202]
  PIN itasel[203]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 798.000 4.000 798.560 ;
    END
  END itasel[203]
  PIN itasel[204]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 800.800 4.000 801.360 ;
    END
  END itasel[204]
  PIN itasel[205]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 803.600 4.000 804.160 ;
    END
  END itasel[205]
  PIN itasel[206]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 806.400 4.000 806.960 ;
    END
  END itasel[206]
  PIN itasel[207]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 809.200 4.000 809.760 ;
    END
  END itasel[207]
  PIN itasel[208]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 812.000 4.000 812.560 ;
    END
  END itasel[208]
  PIN itasel[209]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 814.800 4.000 815.360 ;
    END
  END itasel[209]
  PIN itasel[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 240.800 4.000 241.360 ;
    END
  END itasel[20]
  PIN itasel[210]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 817.600 4.000 818.160 ;
    END
  END itasel[210]
  PIN itasel[211]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 820.400 4.000 820.960 ;
    END
  END itasel[211]
  PIN itasel[212]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 823.200 4.000 823.760 ;
    END
  END itasel[212]
  PIN itasel[213]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 826.000 4.000 826.560 ;
    END
  END itasel[213]
  PIN itasel[214]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 828.800 4.000 829.360 ;
    END
  END itasel[214]
  PIN itasel[215]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 831.600 4.000 832.160 ;
    END
  END itasel[215]
  PIN itasel[216]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 834.400 4.000 834.960 ;
    END
  END itasel[216]
  PIN itasel[217]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 837.200 4.000 837.760 ;
    END
  END itasel[217]
  PIN itasel[218]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 840.000 4.000 840.560 ;
    END
  END itasel[218]
  PIN itasel[219]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 842.800 4.000 843.360 ;
    END
  END itasel[219]
  PIN itasel[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 243.600 4.000 244.160 ;
    END
  END itasel[21]
  PIN itasel[220]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 845.600 4.000 846.160 ;
    END
  END itasel[220]
  PIN itasel[221]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 848.400 4.000 848.960 ;
    END
  END itasel[221]
  PIN itasel[222]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 851.200 4.000 851.760 ;
    END
  END itasel[222]
  PIN itasel[223]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 854.000 4.000 854.560 ;
    END
  END itasel[223]
  PIN itasel[224]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 856.800 4.000 857.360 ;
    END
  END itasel[224]
  PIN itasel[225]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 859.600 4.000 860.160 ;
    END
  END itasel[225]
  PIN itasel[226]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 862.400 4.000 862.960 ;
    END
  END itasel[226]
  PIN itasel[227]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 865.200 4.000 865.760 ;
    END
  END itasel[227]
  PIN itasel[228]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 868.000 4.000 868.560 ;
    END
  END itasel[228]
  PIN itasel[229]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 870.800 4.000 871.360 ;
    END
  END itasel[229]
  PIN itasel[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 246.400 4.000 246.960 ;
    END
  END itasel[22]
  PIN itasel[230]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 873.600 4.000 874.160 ;
    END
  END itasel[230]
  PIN itasel[231]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 876.400 4.000 876.960 ;
    END
  END itasel[231]
  PIN itasel[232]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 879.200 4.000 879.760 ;
    END
  END itasel[232]
  PIN itasel[233]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 882.000 4.000 882.560 ;
    END
  END itasel[233]
  PIN itasel[234]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 884.800 4.000 885.360 ;
    END
  END itasel[234]
  PIN itasel[235]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 887.600 4.000 888.160 ;
    END
  END itasel[235]
  PIN itasel[236]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 890.400 4.000 890.960 ;
    END
  END itasel[236]
  PIN itasel[237]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 893.200 4.000 893.760 ;
    END
  END itasel[237]
  PIN itasel[238]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 896.000 4.000 896.560 ;
    END
  END itasel[238]
  PIN itasel[239]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 898.800 4.000 899.360 ;
    END
  END itasel[239]
  PIN itasel[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 249.200 4.000 249.760 ;
    END
  END itasel[23]
  PIN itasel[240]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 767.200 320.000 767.760 ;
    END
  END itasel[240]
  PIN itasel[241]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 770.000 320.000 770.560 ;
    END
  END itasel[241]
  PIN itasel[242]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 772.800 320.000 773.360 ;
    END
  END itasel[242]
  PIN itasel[243]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 775.600 320.000 776.160 ;
    END
  END itasel[243]
  PIN itasel[244]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 778.400 320.000 778.960 ;
    END
  END itasel[244]
  PIN itasel[245]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 781.200 320.000 781.760 ;
    END
  END itasel[245]
  PIN itasel[246]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 784.000 320.000 784.560 ;
    END
  END itasel[246]
  PIN itasel[247]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 786.800 320.000 787.360 ;
    END
  END itasel[247]
  PIN itasel[248]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 789.600 320.000 790.160 ;
    END
  END itasel[248]
  PIN itasel[249]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 792.400 320.000 792.960 ;
    END
  END itasel[249]
  PIN itasel[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 252.000 4.000 252.560 ;
    END
  END itasel[24]
  PIN itasel[250]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 795.200 320.000 795.760 ;
    END
  END itasel[250]
  PIN itasel[251]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 798.000 320.000 798.560 ;
    END
  END itasel[251]
  PIN itasel[252]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 800.800 320.000 801.360 ;
    END
  END itasel[252]
  PIN itasel[253]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 803.600 320.000 804.160 ;
    END
  END itasel[253]
  PIN itasel[254]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 806.400 320.000 806.960 ;
    END
  END itasel[254]
  PIN itasel[255]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 809.200 320.000 809.760 ;
    END
  END itasel[255]
  PIN itasel[256]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 812.000 320.000 812.560 ;
    END
  END itasel[256]
  PIN itasel[257]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 814.800 320.000 815.360 ;
    END
  END itasel[257]
  PIN itasel[258]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 817.600 320.000 818.160 ;
    END
  END itasel[258]
  PIN itasel[259]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 820.400 320.000 820.960 ;
    END
  END itasel[259]
  PIN itasel[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 254.800 4.000 255.360 ;
    END
  END itasel[25]
  PIN itasel[260]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 823.200 320.000 823.760 ;
    END
  END itasel[260]
  PIN itasel[261]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 826.000 320.000 826.560 ;
    END
  END itasel[261]
  PIN itasel[262]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 828.800 320.000 829.360 ;
    END
  END itasel[262]
  PIN itasel[263]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 831.600 320.000 832.160 ;
    END
  END itasel[263]
  PIN itasel[264]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 834.400 320.000 834.960 ;
    END
  END itasel[264]
  PIN itasel[265]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 837.200 320.000 837.760 ;
    END
  END itasel[265]
  PIN itasel[266]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 840.000 320.000 840.560 ;
    END
  END itasel[266]
  PIN itasel[267]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 842.800 320.000 843.360 ;
    END
  END itasel[267]
  PIN itasel[268]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 845.600 320.000 846.160 ;
    END
  END itasel[268]
  PIN itasel[269]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 848.400 320.000 848.960 ;
    END
  END itasel[269]
  PIN itasel[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 257.600 4.000 258.160 ;
    END
  END itasel[26]
  PIN itasel[270]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 851.200 320.000 851.760 ;
    END
  END itasel[270]
  PIN itasel[271]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 854.000 320.000 854.560 ;
    END
  END itasel[271]
  PIN itasel[272]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 856.800 320.000 857.360 ;
    END
  END itasel[272]
  PIN itasel[273]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 859.600 320.000 860.160 ;
    END
  END itasel[273]
  PIN itasel[274]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 862.400 320.000 862.960 ;
    END
  END itasel[274]
  PIN itasel[275]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 865.200 320.000 865.760 ;
    END
  END itasel[275]
  PIN itasel[276]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 868.000 320.000 868.560 ;
    END
  END itasel[276]
  PIN itasel[277]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 870.800 320.000 871.360 ;
    END
  END itasel[277]
  PIN itasel[278]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 873.600 320.000 874.160 ;
    END
  END itasel[278]
  PIN itasel[279]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 876.400 320.000 876.960 ;
    END
  END itasel[279]
  PIN itasel[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 260.400 4.000 260.960 ;
    END
  END itasel[27]
  PIN itasel[280]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 879.200 320.000 879.760 ;
    END
  END itasel[280]
  PIN itasel[281]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 882.000 320.000 882.560 ;
    END
  END itasel[281]
  PIN itasel[282]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 884.800 320.000 885.360 ;
    END
  END itasel[282]
  PIN itasel[283]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 887.600 320.000 888.160 ;
    END
  END itasel[283]
  PIN itasel[284]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 890.400 320.000 890.960 ;
    END
  END itasel[284]
  PIN itasel[285]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 893.200 320.000 893.760 ;
    END
  END itasel[285]
  PIN itasel[286]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 896.000 320.000 896.560 ;
    END
  END itasel[286]
  PIN itasel[287]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 898.800 320.000 899.360 ;
    END
  END itasel[287]
  PIN itasel[288]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1058.400 4.000 1058.960 ;
    END
  END itasel[288]
  PIN itasel[289]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1061.200 4.000 1061.760 ;
    END
  END itasel[289]
  PIN itasel[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 263.200 4.000 263.760 ;
    END
  END itasel[28]
  PIN itasel[290]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1064.000 4.000 1064.560 ;
    END
  END itasel[290]
  PIN itasel[291]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1066.800 4.000 1067.360 ;
    END
  END itasel[291]
  PIN itasel[292]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1069.600 4.000 1070.160 ;
    END
  END itasel[292]
  PIN itasel[293]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1072.400 4.000 1072.960 ;
    END
  END itasel[293]
  PIN itasel[294]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1075.200 4.000 1075.760 ;
    END
  END itasel[294]
  PIN itasel[295]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1078.000 4.000 1078.560 ;
    END
  END itasel[295]
  PIN itasel[296]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1080.800 4.000 1081.360 ;
    END
  END itasel[296]
  PIN itasel[297]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1083.600 4.000 1084.160 ;
    END
  END itasel[297]
  PIN itasel[298]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1086.400 4.000 1086.960 ;
    END
  END itasel[298]
  PIN itasel[299]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1089.200 4.000 1089.760 ;
    END
  END itasel[299]
  PIN itasel[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 266.000 4.000 266.560 ;
    END
  END itasel[29]
  PIN itasel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 190.400 4.000 190.960 ;
    END
  END itasel[2]
  PIN itasel[300]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1092.000 4.000 1092.560 ;
    END
  END itasel[300]
  PIN itasel[301]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1094.800 4.000 1095.360 ;
    END
  END itasel[301]
  PIN itasel[302]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1097.600 4.000 1098.160 ;
    END
  END itasel[302]
  PIN itasel[303]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1100.400 4.000 1100.960 ;
    END
  END itasel[303]
  PIN itasel[304]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1103.200 4.000 1103.760 ;
    END
  END itasel[304]
  PIN itasel[305]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1106.000 4.000 1106.560 ;
    END
  END itasel[305]
  PIN itasel[306]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1108.800 4.000 1109.360 ;
    END
  END itasel[306]
  PIN itasel[307]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1111.600 4.000 1112.160 ;
    END
  END itasel[307]
  PIN itasel[308]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1114.400 4.000 1114.960 ;
    END
  END itasel[308]
  PIN itasel[309]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1117.200 4.000 1117.760 ;
    END
  END itasel[309]
  PIN itasel[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 268.800 4.000 269.360 ;
    END
  END itasel[30]
  PIN itasel[310]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1120.000 4.000 1120.560 ;
    END
  END itasel[310]
  PIN itasel[311]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1122.800 4.000 1123.360 ;
    END
  END itasel[311]
  PIN itasel[312]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1125.600 4.000 1126.160 ;
    END
  END itasel[312]
  PIN itasel[313]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1128.400 4.000 1128.960 ;
    END
  END itasel[313]
  PIN itasel[314]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1131.200 4.000 1131.760 ;
    END
  END itasel[314]
  PIN itasel[315]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1134.000 4.000 1134.560 ;
    END
  END itasel[315]
  PIN itasel[316]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1136.800 4.000 1137.360 ;
    END
  END itasel[316]
  PIN itasel[317]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1139.600 4.000 1140.160 ;
    END
  END itasel[317]
  PIN itasel[318]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1142.400 4.000 1142.960 ;
    END
  END itasel[318]
  PIN itasel[319]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1145.200 4.000 1145.760 ;
    END
  END itasel[319]
  PIN itasel[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 271.600 4.000 272.160 ;
    END
  END itasel[31]
  PIN itasel[320]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1148.000 4.000 1148.560 ;
    END
  END itasel[320]
  PIN itasel[321]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1150.800 4.000 1151.360 ;
    END
  END itasel[321]
  PIN itasel[322]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1153.600 4.000 1154.160 ;
    END
  END itasel[322]
  PIN itasel[323]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1156.400 4.000 1156.960 ;
    END
  END itasel[323]
  PIN itasel[324]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1159.200 4.000 1159.760 ;
    END
  END itasel[324]
  PIN itasel[325]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1162.000 4.000 1162.560 ;
    END
  END itasel[325]
  PIN itasel[326]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1164.800 4.000 1165.360 ;
    END
  END itasel[326]
  PIN itasel[327]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1167.600 4.000 1168.160 ;
    END
  END itasel[327]
  PIN itasel[328]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1170.400 4.000 1170.960 ;
    END
  END itasel[328]
  PIN itasel[329]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1173.200 4.000 1173.760 ;
    END
  END itasel[329]
  PIN itasel[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 274.400 4.000 274.960 ;
    END
  END itasel[32]
  PIN itasel[330]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1176.000 4.000 1176.560 ;
    END
  END itasel[330]
  PIN itasel[331]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1178.800 4.000 1179.360 ;
    END
  END itasel[331]
  PIN itasel[332]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1181.600 4.000 1182.160 ;
    END
  END itasel[332]
  PIN itasel[333]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1184.400 4.000 1184.960 ;
    END
  END itasel[333]
  PIN itasel[334]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1187.200 4.000 1187.760 ;
    END
  END itasel[334]
  PIN itasel[335]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1190.000 4.000 1190.560 ;
    END
  END itasel[335]
  PIN itasel[336]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1058.400 320.000 1058.960 ;
    END
  END itasel[336]
  PIN itasel[337]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1061.200 320.000 1061.760 ;
    END
  END itasel[337]
  PIN itasel[338]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1064.000 320.000 1064.560 ;
    END
  END itasel[338]
  PIN itasel[339]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1066.800 320.000 1067.360 ;
    END
  END itasel[339]
  PIN itasel[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 277.200 4.000 277.760 ;
    END
  END itasel[33]
  PIN itasel[340]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1069.600 320.000 1070.160 ;
    END
  END itasel[340]
  PIN itasel[341]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1072.400 320.000 1072.960 ;
    END
  END itasel[341]
  PIN itasel[342]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1075.200 320.000 1075.760 ;
    END
  END itasel[342]
  PIN itasel[343]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1078.000 320.000 1078.560 ;
    END
  END itasel[343]
  PIN itasel[344]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1080.800 320.000 1081.360 ;
    END
  END itasel[344]
  PIN itasel[345]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1083.600 320.000 1084.160 ;
    END
  END itasel[345]
  PIN itasel[346]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1086.400 320.000 1086.960 ;
    END
  END itasel[346]
  PIN itasel[347]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1089.200 320.000 1089.760 ;
    END
  END itasel[347]
  PIN itasel[348]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1092.000 320.000 1092.560 ;
    END
  END itasel[348]
  PIN itasel[349]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1094.800 320.000 1095.360 ;
    END
  END itasel[349]
  PIN itasel[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 280.000 4.000 280.560 ;
    END
  END itasel[34]
  PIN itasel[350]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1097.600 320.000 1098.160 ;
    END
  END itasel[350]
  PIN itasel[351]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1100.400 320.000 1100.960 ;
    END
  END itasel[351]
  PIN itasel[352]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1103.200 320.000 1103.760 ;
    END
  END itasel[352]
  PIN itasel[353]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1106.000 320.000 1106.560 ;
    END
  END itasel[353]
  PIN itasel[354]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1108.800 320.000 1109.360 ;
    END
  END itasel[354]
  PIN itasel[355]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1111.600 320.000 1112.160 ;
    END
  END itasel[355]
  PIN itasel[356]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1114.400 320.000 1114.960 ;
    END
  END itasel[356]
  PIN itasel[357]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1117.200 320.000 1117.760 ;
    END
  END itasel[357]
  PIN itasel[358]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1120.000 320.000 1120.560 ;
    END
  END itasel[358]
  PIN itasel[359]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1122.800 320.000 1123.360 ;
    END
  END itasel[359]
  PIN itasel[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 282.800 4.000 283.360 ;
    END
  END itasel[35]
  PIN itasel[360]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1125.600 320.000 1126.160 ;
    END
  END itasel[360]
  PIN itasel[361]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1128.400 320.000 1128.960 ;
    END
  END itasel[361]
  PIN itasel[362]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1131.200 320.000 1131.760 ;
    END
  END itasel[362]
  PIN itasel[363]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1134.000 320.000 1134.560 ;
    END
  END itasel[363]
  PIN itasel[364]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1136.800 320.000 1137.360 ;
    END
  END itasel[364]
  PIN itasel[365]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1139.600 320.000 1140.160 ;
    END
  END itasel[365]
  PIN itasel[366]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1142.400 320.000 1142.960 ;
    END
  END itasel[366]
  PIN itasel[367]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1145.200 320.000 1145.760 ;
    END
  END itasel[367]
  PIN itasel[368]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1148.000 320.000 1148.560 ;
    END
  END itasel[368]
  PIN itasel[369]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1150.800 320.000 1151.360 ;
    END
  END itasel[369]
  PIN itasel[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 285.600 4.000 286.160 ;
    END
  END itasel[36]
  PIN itasel[370]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1153.600 320.000 1154.160 ;
    END
  END itasel[370]
  PIN itasel[371]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1156.400 320.000 1156.960 ;
    END
  END itasel[371]
  PIN itasel[372]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1159.200 320.000 1159.760 ;
    END
  END itasel[372]
  PIN itasel[373]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1162.000 320.000 1162.560 ;
    END
  END itasel[373]
  PIN itasel[374]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1164.800 320.000 1165.360 ;
    END
  END itasel[374]
  PIN itasel[375]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1167.600 320.000 1168.160 ;
    END
  END itasel[375]
  PIN itasel[376]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1170.400 320.000 1170.960 ;
    END
  END itasel[376]
  PIN itasel[377]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1173.200 320.000 1173.760 ;
    END
  END itasel[377]
  PIN itasel[378]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1176.000 320.000 1176.560 ;
    END
  END itasel[378]
  PIN itasel[379]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1178.800 320.000 1179.360 ;
    END
  END itasel[379]
  PIN itasel[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 288.400 4.000 288.960 ;
    END
  END itasel[37]
  PIN itasel[380]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1181.600 320.000 1182.160 ;
    END
  END itasel[380]
  PIN itasel[381]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1184.400 320.000 1184.960 ;
    END
  END itasel[381]
  PIN itasel[382]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1187.200 320.000 1187.760 ;
    END
  END itasel[382]
  PIN itasel[383]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1190.000 320.000 1190.560 ;
    END
  END itasel[383]
  PIN itasel[384]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1349.600 4.000 1350.160 ;
    END
  END itasel[384]
  PIN itasel[385]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1352.400 4.000 1352.960 ;
    END
  END itasel[385]
  PIN itasel[386]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1355.200 4.000 1355.760 ;
    END
  END itasel[386]
  PIN itasel[387]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1358.000 4.000 1358.560 ;
    END
  END itasel[387]
  PIN itasel[388]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1360.800 4.000 1361.360 ;
    END
  END itasel[388]
  PIN itasel[389]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1363.600 4.000 1364.160 ;
    END
  END itasel[389]
  PIN itasel[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 291.200 4.000 291.760 ;
    END
  END itasel[38]
  PIN itasel[390]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1366.400 4.000 1366.960 ;
    END
  END itasel[390]
  PIN itasel[391]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1369.200 4.000 1369.760 ;
    END
  END itasel[391]
  PIN itasel[392]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1372.000 4.000 1372.560 ;
    END
  END itasel[392]
  PIN itasel[393]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1374.800 4.000 1375.360 ;
    END
  END itasel[393]
  PIN itasel[394]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1377.600 4.000 1378.160 ;
    END
  END itasel[394]
  PIN itasel[395]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1380.400 4.000 1380.960 ;
    END
  END itasel[395]
  PIN itasel[396]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1383.200 4.000 1383.760 ;
    END
  END itasel[396]
  PIN itasel[397]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1386.000 4.000 1386.560 ;
    END
  END itasel[397]
  PIN itasel[398]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1388.800 4.000 1389.360 ;
    END
  END itasel[398]
  PIN itasel[399]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1391.600 4.000 1392.160 ;
    END
  END itasel[399]
  PIN itasel[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 294.000 4.000 294.560 ;
    END
  END itasel[39]
  PIN itasel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 193.200 4.000 193.760 ;
    END
  END itasel[3]
  PIN itasel[400]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1394.400 4.000 1394.960 ;
    END
  END itasel[400]
  PIN itasel[401]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1397.200 4.000 1397.760 ;
    END
  END itasel[401]
  PIN itasel[402]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1400.000 4.000 1400.560 ;
    END
  END itasel[402]
  PIN itasel[403]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1402.800 4.000 1403.360 ;
    END
  END itasel[403]
  PIN itasel[404]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1405.600 4.000 1406.160 ;
    END
  END itasel[404]
  PIN itasel[405]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1408.400 4.000 1408.960 ;
    END
  END itasel[405]
  PIN itasel[406]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1411.200 4.000 1411.760 ;
    END
  END itasel[406]
  PIN itasel[407]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1414.000 4.000 1414.560 ;
    END
  END itasel[407]
  PIN itasel[408]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1416.800 4.000 1417.360 ;
    END
  END itasel[408]
  PIN itasel[409]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1419.600 4.000 1420.160 ;
    END
  END itasel[409]
  PIN itasel[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 296.800 4.000 297.360 ;
    END
  END itasel[40]
  PIN itasel[410]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1422.400 4.000 1422.960 ;
    END
  END itasel[410]
  PIN itasel[411]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1425.200 4.000 1425.760 ;
    END
  END itasel[411]
  PIN itasel[412]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1428.000 4.000 1428.560 ;
    END
  END itasel[412]
  PIN itasel[413]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1430.800 4.000 1431.360 ;
    END
  END itasel[413]
  PIN itasel[414]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1433.600 4.000 1434.160 ;
    END
  END itasel[414]
  PIN itasel[415]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1436.400 4.000 1436.960 ;
    END
  END itasel[415]
  PIN itasel[416]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1439.200 4.000 1439.760 ;
    END
  END itasel[416]
  PIN itasel[417]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1442.000 4.000 1442.560 ;
    END
  END itasel[417]
  PIN itasel[418]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1444.800 4.000 1445.360 ;
    END
  END itasel[418]
  PIN itasel[419]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1447.600 4.000 1448.160 ;
    END
  END itasel[419]
  PIN itasel[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 299.600 4.000 300.160 ;
    END
  END itasel[41]
  PIN itasel[420]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1450.400 4.000 1450.960 ;
    END
  END itasel[420]
  PIN itasel[421]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1453.200 4.000 1453.760 ;
    END
  END itasel[421]
  PIN itasel[422]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1456.000 4.000 1456.560 ;
    END
  END itasel[422]
  PIN itasel[423]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1458.800 4.000 1459.360 ;
    END
  END itasel[423]
  PIN itasel[424]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1461.600 4.000 1462.160 ;
    END
  END itasel[424]
  PIN itasel[425]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1464.400 4.000 1464.960 ;
    END
  END itasel[425]
  PIN itasel[426]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1467.200 4.000 1467.760 ;
    END
  END itasel[426]
  PIN itasel[427]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1470.000 4.000 1470.560 ;
    END
  END itasel[427]
  PIN itasel[428]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1472.800 4.000 1473.360 ;
    END
  END itasel[428]
  PIN itasel[429]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1475.600 4.000 1476.160 ;
    END
  END itasel[429]
  PIN itasel[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 302.400 4.000 302.960 ;
    END
  END itasel[42]
  PIN itasel[430]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1478.400 4.000 1478.960 ;
    END
  END itasel[430]
  PIN itasel[431]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1481.200 4.000 1481.760 ;
    END
  END itasel[431]
  PIN itasel[432]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1349.600 320.000 1350.160 ;
    END
  END itasel[432]
  PIN itasel[433]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1352.400 320.000 1352.960 ;
    END
  END itasel[433]
  PIN itasel[434]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1355.200 320.000 1355.760 ;
    END
  END itasel[434]
  PIN itasel[435]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1358.000 320.000 1358.560 ;
    END
  END itasel[435]
  PIN itasel[436]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1360.800 320.000 1361.360 ;
    END
  END itasel[436]
  PIN itasel[437]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1363.600 320.000 1364.160 ;
    END
  END itasel[437]
  PIN itasel[438]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1366.400 320.000 1366.960 ;
    END
  END itasel[438]
  PIN itasel[439]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1369.200 320.000 1369.760 ;
    END
  END itasel[439]
  PIN itasel[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 305.200 4.000 305.760 ;
    END
  END itasel[43]
  PIN itasel[440]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1372.000 320.000 1372.560 ;
    END
  END itasel[440]
  PIN itasel[441]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1374.800 320.000 1375.360 ;
    END
  END itasel[441]
  PIN itasel[442]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1377.600 320.000 1378.160 ;
    END
  END itasel[442]
  PIN itasel[443]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1380.400 320.000 1380.960 ;
    END
  END itasel[443]
  PIN itasel[444]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1383.200 320.000 1383.760 ;
    END
  END itasel[444]
  PIN itasel[445]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1386.000 320.000 1386.560 ;
    END
  END itasel[445]
  PIN itasel[446]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1388.800 320.000 1389.360 ;
    END
  END itasel[446]
  PIN itasel[447]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1391.600 320.000 1392.160 ;
    END
  END itasel[447]
  PIN itasel[448]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1394.400 320.000 1394.960 ;
    END
  END itasel[448]
  PIN itasel[449]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1397.200 320.000 1397.760 ;
    END
  END itasel[449]
  PIN itasel[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 308.000 4.000 308.560 ;
    END
  END itasel[44]
  PIN itasel[450]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1400.000 320.000 1400.560 ;
    END
  END itasel[450]
  PIN itasel[451]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1402.800 320.000 1403.360 ;
    END
  END itasel[451]
  PIN itasel[452]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1405.600 320.000 1406.160 ;
    END
  END itasel[452]
  PIN itasel[453]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1408.400 320.000 1408.960 ;
    END
  END itasel[453]
  PIN itasel[454]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1411.200 320.000 1411.760 ;
    END
  END itasel[454]
  PIN itasel[455]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1414.000 320.000 1414.560 ;
    END
  END itasel[455]
  PIN itasel[456]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1416.800 320.000 1417.360 ;
    END
  END itasel[456]
  PIN itasel[457]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1419.600 320.000 1420.160 ;
    END
  END itasel[457]
  PIN itasel[458]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1422.400 320.000 1422.960 ;
    END
  END itasel[458]
  PIN itasel[459]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1425.200 320.000 1425.760 ;
    END
  END itasel[459]
  PIN itasel[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 310.800 4.000 311.360 ;
    END
  END itasel[45]
  PIN itasel[460]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1428.000 320.000 1428.560 ;
    END
  END itasel[460]
  PIN itasel[461]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1430.800 320.000 1431.360 ;
    END
  END itasel[461]
  PIN itasel[462]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1433.600 320.000 1434.160 ;
    END
  END itasel[462]
  PIN itasel[463]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1436.400 320.000 1436.960 ;
    END
  END itasel[463]
  PIN itasel[464]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1439.200 320.000 1439.760 ;
    END
  END itasel[464]
  PIN itasel[465]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1442.000 320.000 1442.560 ;
    END
  END itasel[465]
  PIN itasel[466]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1444.800 320.000 1445.360 ;
    END
  END itasel[466]
  PIN itasel[467]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1447.600 320.000 1448.160 ;
    END
  END itasel[467]
  PIN itasel[468]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1450.400 320.000 1450.960 ;
    END
  END itasel[468]
  PIN itasel[469]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1453.200 320.000 1453.760 ;
    END
  END itasel[469]
  PIN itasel[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 313.600 4.000 314.160 ;
    END
  END itasel[46]
  PIN itasel[470]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1456.000 320.000 1456.560 ;
    END
  END itasel[470]
  PIN itasel[471]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1458.800 320.000 1459.360 ;
    END
  END itasel[471]
  PIN itasel[472]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1461.600 320.000 1462.160 ;
    END
  END itasel[472]
  PIN itasel[473]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1464.400 320.000 1464.960 ;
    END
  END itasel[473]
  PIN itasel[474]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1467.200 320.000 1467.760 ;
    END
  END itasel[474]
  PIN itasel[475]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1470.000 320.000 1470.560 ;
    END
  END itasel[475]
  PIN itasel[476]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1472.800 320.000 1473.360 ;
    END
  END itasel[476]
  PIN itasel[477]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1475.600 320.000 1476.160 ;
    END
  END itasel[477]
  PIN itasel[478]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1478.400 320.000 1478.960 ;
    END
  END itasel[478]
  PIN itasel[479]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1481.200 320.000 1481.760 ;
    END
  END itasel[479]
  PIN itasel[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 316.400 4.000 316.960 ;
    END
  END itasel[47]
  PIN itasel[480]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1640.800 4.000 1641.360 ;
    END
  END itasel[480]
  PIN itasel[481]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1643.600 4.000 1644.160 ;
    END
  END itasel[481]
  PIN itasel[482]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1646.400 4.000 1646.960 ;
    END
  END itasel[482]
  PIN itasel[483]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1649.200 4.000 1649.760 ;
    END
  END itasel[483]
  PIN itasel[484]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1652.000 4.000 1652.560 ;
    END
  END itasel[484]
  PIN itasel[485]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1654.800 4.000 1655.360 ;
    END
  END itasel[485]
  PIN itasel[486]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1657.600 4.000 1658.160 ;
    END
  END itasel[486]
  PIN itasel[487]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1660.400 4.000 1660.960 ;
    END
  END itasel[487]
  PIN itasel[488]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1663.200 4.000 1663.760 ;
    END
  END itasel[488]
  PIN itasel[489]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1666.000 4.000 1666.560 ;
    END
  END itasel[489]
  PIN itasel[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 184.800 320.000 185.360 ;
    END
  END itasel[48]
  PIN itasel[490]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1668.800 4.000 1669.360 ;
    END
  END itasel[490]
  PIN itasel[491]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1671.600 4.000 1672.160 ;
    END
  END itasel[491]
  PIN itasel[492]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1674.400 4.000 1674.960 ;
    END
  END itasel[492]
  PIN itasel[493]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1677.200 4.000 1677.760 ;
    END
  END itasel[493]
  PIN itasel[494]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1680.000 4.000 1680.560 ;
    END
  END itasel[494]
  PIN itasel[495]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1682.800 4.000 1683.360 ;
    END
  END itasel[495]
  PIN itasel[496]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1685.600 4.000 1686.160 ;
    END
  END itasel[496]
  PIN itasel[497]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1688.400 4.000 1688.960 ;
    END
  END itasel[497]
  PIN itasel[498]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1691.200 4.000 1691.760 ;
    END
  END itasel[498]
  PIN itasel[499]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1694.000 4.000 1694.560 ;
    END
  END itasel[499]
  PIN itasel[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 187.600 320.000 188.160 ;
    END
  END itasel[49]
  PIN itasel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 196.000 4.000 196.560 ;
    END
  END itasel[4]
  PIN itasel[500]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1696.800 4.000 1697.360 ;
    END
  END itasel[500]
  PIN itasel[501]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1699.600 4.000 1700.160 ;
    END
  END itasel[501]
  PIN itasel[502]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1702.400 4.000 1702.960 ;
    END
  END itasel[502]
  PIN itasel[503]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1705.200 4.000 1705.760 ;
    END
  END itasel[503]
  PIN itasel[504]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1708.000 4.000 1708.560 ;
    END
  END itasel[504]
  PIN itasel[505]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1710.800 4.000 1711.360 ;
    END
  END itasel[505]
  PIN itasel[506]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1713.600 4.000 1714.160 ;
    END
  END itasel[506]
  PIN itasel[507]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1716.400 4.000 1716.960 ;
    END
  END itasel[507]
  PIN itasel[508]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1719.200 4.000 1719.760 ;
    END
  END itasel[508]
  PIN itasel[509]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1722.000 4.000 1722.560 ;
    END
  END itasel[509]
  PIN itasel[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 190.400 320.000 190.960 ;
    END
  END itasel[50]
  PIN itasel[510]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1724.800 4.000 1725.360 ;
    END
  END itasel[510]
  PIN itasel[511]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1727.600 4.000 1728.160 ;
    END
  END itasel[511]
  PIN itasel[512]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1730.400 4.000 1730.960 ;
    END
  END itasel[512]
  PIN itasel[513]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1733.200 4.000 1733.760 ;
    END
  END itasel[513]
  PIN itasel[514]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1736.000 4.000 1736.560 ;
    END
  END itasel[514]
  PIN itasel[515]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1738.800 4.000 1739.360 ;
    END
  END itasel[515]
  PIN itasel[516]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1741.600 4.000 1742.160 ;
    END
  END itasel[516]
  PIN itasel[517]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1744.400 4.000 1744.960 ;
    END
  END itasel[517]
  PIN itasel[518]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1747.200 4.000 1747.760 ;
    END
  END itasel[518]
  PIN itasel[519]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1750.000 4.000 1750.560 ;
    END
  END itasel[519]
  PIN itasel[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 193.200 320.000 193.760 ;
    END
  END itasel[51]
  PIN itasel[520]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1752.800 4.000 1753.360 ;
    END
  END itasel[520]
  PIN itasel[521]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1755.600 4.000 1756.160 ;
    END
  END itasel[521]
  PIN itasel[522]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1758.400 4.000 1758.960 ;
    END
  END itasel[522]
  PIN itasel[523]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1761.200 4.000 1761.760 ;
    END
  END itasel[523]
  PIN itasel[524]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1764.000 4.000 1764.560 ;
    END
  END itasel[524]
  PIN itasel[525]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1766.800 4.000 1767.360 ;
    END
  END itasel[525]
  PIN itasel[526]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1769.600 4.000 1770.160 ;
    END
  END itasel[526]
  PIN itasel[527]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1772.400 4.000 1772.960 ;
    END
  END itasel[527]
  PIN itasel[528]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1640.800 320.000 1641.360 ;
    END
  END itasel[528]
  PIN itasel[529]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1643.600 320.000 1644.160 ;
    END
  END itasel[529]
  PIN itasel[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 196.000 320.000 196.560 ;
    END
  END itasel[52]
  PIN itasel[530]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1646.400 320.000 1646.960 ;
    END
  END itasel[530]
  PIN itasel[531]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1649.200 320.000 1649.760 ;
    END
  END itasel[531]
  PIN itasel[532]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1652.000 320.000 1652.560 ;
    END
  END itasel[532]
  PIN itasel[533]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1654.800 320.000 1655.360 ;
    END
  END itasel[533]
  PIN itasel[534]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1657.600 320.000 1658.160 ;
    END
  END itasel[534]
  PIN itasel[535]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1660.400 320.000 1660.960 ;
    END
  END itasel[535]
  PIN itasel[536]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1663.200 320.000 1663.760 ;
    END
  END itasel[536]
  PIN itasel[537]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1666.000 320.000 1666.560 ;
    END
  END itasel[537]
  PIN itasel[538]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1668.800 320.000 1669.360 ;
    END
  END itasel[538]
  PIN itasel[539]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1671.600 320.000 1672.160 ;
    END
  END itasel[539]
  PIN itasel[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 198.800 320.000 199.360 ;
    END
  END itasel[53]
  PIN itasel[540]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1674.400 320.000 1674.960 ;
    END
  END itasel[540]
  PIN itasel[541]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1677.200 320.000 1677.760 ;
    END
  END itasel[541]
  PIN itasel[542]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1680.000 320.000 1680.560 ;
    END
  END itasel[542]
  PIN itasel[543]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1682.800 320.000 1683.360 ;
    END
  END itasel[543]
  PIN itasel[544]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1685.600 320.000 1686.160 ;
    END
  END itasel[544]
  PIN itasel[545]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1688.400 320.000 1688.960 ;
    END
  END itasel[545]
  PIN itasel[546]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1691.200 320.000 1691.760 ;
    END
  END itasel[546]
  PIN itasel[547]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1694.000 320.000 1694.560 ;
    END
  END itasel[547]
  PIN itasel[548]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1696.800 320.000 1697.360 ;
    END
  END itasel[548]
  PIN itasel[549]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1699.600 320.000 1700.160 ;
    END
  END itasel[549]
  PIN itasel[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 201.600 320.000 202.160 ;
    END
  END itasel[54]
  PIN itasel[550]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1702.400 320.000 1702.960 ;
    END
  END itasel[550]
  PIN itasel[551]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1705.200 320.000 1705.760 ;
    END
  END itasel[551]
  PIN itasel[552]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1708.000 320.000 1708.560 ;
    END
  END itasel[552]
  PIN itasel[553]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1710.800 320.000 1711.360 ;
    END
  END itasel[553]
  PIN itasel[554]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1713.600 320.000 1714.160 ;
    END
  END itasel[554]
  PIN itasel[555]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1716.400 320.000 1716.960 ;
    END
  END itasel[555]
  PIN itasel[556]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1719.200 320.000 1719.760 ;
    END
  END itasel[556]
  PIN itasel[557]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1722.000 320.000 1722.560 ;
    END
  END itasel[557]
  PIN itasel[558]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1724.800 320.000 1725.360 ;
    END
  END itasel[558]
  PIN itasel[559]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1727.600 320.000 1728.160 ;
    END
  END itasel[559]
  PIN itasel[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 204.400 320.000 204.960 ;
    END
  END itasel[55]
  PIN itasel[560]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1730.400 320.000 1730.960 ;
    END
  END itasel[560]
  PIN itasel[561]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1733.200 320.000 1733.760 ;
    END
  END itasel[561]
  PIN itasel[562]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1736.000 320.000 1736.560 ;
    END
  END itasel[562]
  PIN itasel[563]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1738.800 320.000 1739.360 ;
    END
  END itasel[563]
  PIN itasel[564]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1741.600 320.000 1742.160 ;
    END
  END itasel[564]
  PIN itasel[565]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1744.400 320.000 1744.960 ;
    END
  END itasel[565]
  PIN itasel[566]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1747.200 320.000 1747.760 ;
    END
  END itasel[566]
  PIN itasel[567]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1750.000 320.000 1750.560 ;
    END
  END itasel[567]
  PIN itasel[568]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1752.800 320.000 1753.360 ;
    END
  END itasel[568]
  PIN itasel[569]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1755.600 320.000 1756.160 ;
    END
  END itasel[569]
  PIN itasel[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 207.200 320.000 207.760 ;
    END
  END itasel[56]
  PIN itasel[570]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1758.400 320.000 1758.960 ;
    END
  END itasel[570]
  PIN itasel[571]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1761.200 320.000 1761.760 ;
    END
  END itasel[571]
  PIN itasel[572]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1764.000 320.000 1764.560 ;
    END
  END itasel[572]
  PIN itasel[573]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1766.800 320.000 1767.360 ;
    END
  END itasel[573]
  PIN itasel[574]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1769.600 320.000 1770.160 ;
    END
  END itasel[574]
  PIN itasel[575]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1772.400 320.000 1772.960 ;
    END
  END itasel[575]
  PIN itasel[576]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1932.000 4.000 1932.560 ;
    END
  END itasel[576]
  PIN itasel[577]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1934.800 4.000 1935.360 ;
    END
  END itasel[577]
  PIN itasel[578]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1937.600 4.000 1938.160 ;
    END
  END itasel[578]
  PIN itasel[579]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1940.400 4.000 1940.960 ;
    END
  END itasel[579]
  PIN itasel[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 210.000 320.000 210.560 ;
    END
  END itasel[57]
  PIN itasel[580]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1943.200 4.000 1943.760 ;
    END
  END itasel[580]
  PIN itasel[581]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1946.000 4.000 1946.560 ;
    END
  END itasel[581]
  PIN itasel[582]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1948.800 4.000 1949.360 ;
    END
  END itasel[582]
  PIN itasel[583]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1951.600 4.000 1952.160 ;
    END
  END itasel[583]
  PIN itasel[584]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1954.400 4.000 1954.960 ;
    END
  END itasel[584]
  PIN itasel[585]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1957.200 4.000 1957.760 ;
    END
  END itasel[585]
  PIN itasel[586]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1960.000 4.000 1960.560 ;
    END
  END itasel[586]
  PIN itasel[587]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1962.800 4.000 1963.360 ;
    END
  END itasel[587]
  PIN itasel[588]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1965.600 4.000 1966.160 ;
    END
  END itasel[588]
  PIN itasel[589]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1968.400 4.000 1968.960 ;
    END
  END itasel[589]
  PIN itasel[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 212.800 320.000 213.360 ;
    END
  END itasel[58]
  PIN itasel[590]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1971.200 4.000 1971.760 ;
    END
  END itasel[590]
  PIN itasel[591]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1974.000 4.000 1974.560 ;
    END
  END itasel[591]
  PIN itasel[592]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1976.800 4.000 1977.360 ;
    END
  END itasel[592]
  PIN itasel[593]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1979.600 4.000 1980.160 ;
    END
  END itasel[593]
  PIN itasel[594]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1982.400 4.000 1982.960 ;
    END
  END itasel[594]
  PIN itasel[595]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1985.200 4.000 1985.760 ;
    END
  END itasel[595]
  PIN itasel[596]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1988.000 4.000 1988.560 ;
    END
  END itasel[596]
  PIN itasel[597]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1990.800 4.000 1991.360 ;
    END
  END itasel[597]
  PIN itasel[598]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1993.600 4.000 1994.160 ;
    END
  END itasel[598]
  PIN itasel[599]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1996.400 4.000 1996.960 ;
    END
  END itasel[599]
  PIN itasel[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 215.600 320.000 216.160 ;
    END
  END itasel[59]
  PIN itasel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 198.800 4.000 199.360 ;
    END
  END itasel[5]
  PIN itasel[600]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1999.200 4.000 1999.760 ;
    END
  END itasel[600]
  PIN itasel[601]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2002.000 4.000 2002.560 ;
    END
  END itasel[601]
  PIN itasel[602]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2004.800 4.000 2005.360 ;
    END
  END itasel[602]
  PIN itasel[603]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2007.600 4.000 2008.160 ;
    END
  END itasel[603]
  PIN itasel[604]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2010.400 4.000 2010.960 ;
    END
  END itasel[604]
  PIN itasel[605]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2013.200 4.000 2013.760 ;
    END
  END itasel[605]
  PIN itasel[606]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2016.000 4.000 2016.560 ;
    END
  END itasel[606]
  PIN itasel[607]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2018.800 4.000 2019.360 ;
    END
  END itasel[607]
  PIN itasel[608]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2021.600 4.000 2022.160 ;
    END
  END itasel[608]
  PIN itasel[609]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2024.400 4.000 2024.960 ;
    END
  END itasel[609]
  PIN itasel[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 218.400 320.000 218.960 ;
    END
  END itasel[60]
  PIN itasel[610]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2027.200 4.000 2027.760 ;
    END
  END itasel[610]
  PIN itasel[611]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2030.000 4.000 2030.560 ;
    END
  END itasel[611]
  PIN itasel[612]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2032.800 4.000 2033.360 ;
    END
  END itasel[612]
  PIN itasel[613]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2035.600 4.000 2036.160 ;
    END
  END itasel[613]
  PIN itasel[614]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2038.400 4.000 2038.960 ;
    END
  END itasel[614]
  PIN itasel[615]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2041.200 4.000 2041.760 ;
    END
  END itasel[615]
  PIN itasel[616]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2044.000 4.000 2044.560 ;
    END
  END itasel[616]
  PIN itasel[617]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2046.800 4.000 2047.360 ;
    END
  END itasel[617]
  PIN itasel[618]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2049.600 4.000 2050.160 ;
    END
  END itasel[618]
  PIN itasel[619]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2052.400 4.000 2052.960 ;
    END
  END itasel[619]
  PIN itasel[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 221.200 320.000 221.760 ;
    END
  END itasel[61]
  PIN itasel[620]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2055.200 4.000 2055.760 ;
    END
  END itasel[620]
  PIN itasel[621]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2058.000 4.000 2058.560 ;
    END
  END itasel[621]
  PIN itasel[622]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2060.800 4.000 2061.360 ;
    END
  END itasel[622]
  PIN itasel[623]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2063.600 4.000 2064.160 ;
    END
  END itasel[623]
  PIN itasel[624]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1932.000 320.000 1932.560 ;
    END
  END itasel[624]
  PIN itasel[625]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1934.800 320.000 1935.360 ;
    END
  END itasel[625]
  PIN itasel[626]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1937.600 320.000 1938.160 ;
    END
  END itasel[626]
  PIN itasel[627]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1940.400 320.000 1940.960 ;
    END
  END itasel[627]
  PIN itasel[628]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1943.200 320.000 1943.760 ;
    END
  END itasel[628]
  PIN itasel[629]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1946.000 320.000 1946.560 ;
    END
  END itasel[629]
  PIN itasel[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 224.000 320.000 224.560 ;
    END
  END itasel[62]
  PIN itasel[630]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1948.800 320.000 1949.360 ;
    END
  END itasel[630]
  PIN itasel[631]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1951.600 320.000 1952.160 ;
    END
  END itasel[631]
  PIN itasel[632]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1954.400 320.000 1954.960 ;
    END
  END itasel[632]
  PIN itasel[633]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1957.200 320.000 1957.760 ;
    END
  END itasel[633]
  PIN itasel[634]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1960.000 320.000 1960.560 ;
    END
  END itasel[634]
  PIN itasel[635]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1962.800 320.000 1963.360 ;
    END
  END itasel[635]
  PIN itasel[636]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1965.600 320.000 1966.160 ;
    END
  END itasel[636]
  PIN itasel[637]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1968.400 320.000 1968.960 ;
    END
  END itasel[637]
  PIN itasel[638]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1971.200 320.000 1971.760 ;
    END
  END itasel[638]
  PIN itasel[639]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1974.000 320.000 1974.560 ;
    END
  END itasel[639]
  PIN itasel[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 226.800 320.000 227.360 ;
    END
  END itasel[63]
  PIN itasel[640]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1976.800 320.000 1977.360 ;
    END
  END itasel[640]
  PIN itasel[641]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1979.600 320.000 1980.160 ;
    END
  END itasel[641]
  PIN itasel[642]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1982.400 320.000 1982.960 ;
    END
  END itasel[642]
  PIN itasel[643]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1985.200 320.000 1985.760 ;
    END
  END itasel[643]
  PIN itasel[644]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1988.000 320.000 1988.560 ;
    END
  END itasel[644]
  PIN itasel[645]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1990.800 320.000 1991.360 ;
    END
  END itasel[645]
  PIN itasel[646]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1993.600 320.000 1994.160 ;
    END
  END itasel[646]
  PIN itasel[647]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1996.400 320.000 1996.960 ;
    END
  END itasel[647]
  PIN itasel[648]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 1999.200 320.000 1999.760 ;
    END
  END itasel[648]
  PIN itasel[649]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2002.000 320.000 2002.560 ;
    END
  END itasel[649]
  PIN itasel[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 229.600 320.000 230.160 ;
    END
  END itasel[64]
  PIN itasel[650]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2004.800 320.000 2005.360 ;
    END
  END itasel[650]
  PIN itasel[651]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2007.600 320.000 2008.160 ;
    END
  END itasel[651]
  PIN itasel[652]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2010.400 320.000 2010.960 ;
    END
  END itasel[652]
  PIN itasel[653]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2013.200 320.000 2013.760 ;
    END
  END itasel[653]
  PIN itasel[654]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2016.000 320.000 2016.560 ;
    END
  END itasel[654]
  PIN itasel[655]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2018.800 320.000 2019.360 ;
    END
  END itasel[655]
  PIN itasel[656]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2021.600 320.000 2022.160 ;
    END
  END itasel[656]
  PIN itasel[657]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2024.400 320.000 2024.960 ;
    END
  END itasel[657]
  PIN itasel[658]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2027.200 320.000 2027.760 ;
    END
  END itasel[658]
  PIN itasel[659]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2030.000 320.000 2030.560 ;
    END
  END itasel[659]
  PIN itasel[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 232.400 320.000 232.960 ;
    END
  END itasel[65]
  PIN itasel[660]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2032.800 320.000 2033.360 ;
    END
  END itasel[660]
  PIN itasel[661]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2035.600 320.000 2036.160 ;
    END
  END itasel[661]
  PIN itasel[662]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2038.400 320.000 2038.960 ;
    END
  END itasel[662]
  PIN itasel[663]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2041.200 320.000 2041.760 ;
    END
  END itasel[663]
  PIN itasel[664]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2044.000 320.000 2044.560 ;
    END
  END itasel[664]
  PIN itasel[665]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2046.800 320.000 2047.360 ;
    END
  END itasel[665]
  PIN itasel[666]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2049.600 320.000 2050.160 ;
    END
  END itasel[666]
  PIN itasel[667]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2052.400 320.000 2052.960 ;
    END
  END itasel[667]
  PIN itasel[668]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.408000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2055.200 320.000 2055.760 ;
    END
  END itasel[668]
  PIN itasel[669]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.408000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2058.000 320.000 2058.560 ;
    END
  END itasel[669]
  PIN itasel[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 235.200 320.000 235.760 ;
    END
  END itasel[66]
  PIN itasel[670]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2060.800 320.000 2061.360 ;
    END
  END itasel[670]
  PIN itasel[671]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2063.600 320.000 2064.160 ;
    END
  END itasel[671]
  PIN itasel[672]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2223.200 4.000 2223.760 ;
    END
  END itasel[672]
  PIN itasel[673]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2226.000 4.000 2226.560 ;
    END
  END itasel[673]
  PIN itasel[674]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2228.800 4.000 2229.360 ;
    END
  END itasel[674]
  PIN itasel[675]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2231.600 4.000 2232.160 ;
    END
  END itasel[675]
  PIN itasel[676]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2234.400 4.000 2234.960 ;
    END
  END itasel[676]
  PIN itasel[677]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2237.200 4.000 2237.760 ;
    END
  END itasel[677]
  PIN itasel[678]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2240.000 4.000 2240.560 ;
    END
  END itasel[678]
  PIN itasel[679]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2242.800 4.000 2243.360 ;
    END
  END itasel[679]
  PIN itasel[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 238.000 320.000 238.560 ;
    END
  END itasel[67]
  PIN itasel[680]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2245.600 4.000 2246.160 ;
    END
  END itasel[680]
  PIN itasel[681]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2248.400 4.000 2248.960 ;
    END
  END itasel[681]
  PIN itasel[682]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2251.200 4.000 2251.760 ;
    END
  END itasel[682]
  PIN itasel[683]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2254.000 4.000 2254.560 ;
    END
  END itasel[683]
  PIN itasel[684]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2256.800 4.000 2257.360 ;
    END
  END itasel[684]
  PIN itasel[685]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2259.600 4.000 2260.160 ;
    END
  END itasel[685]
  PIN itasel[686]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2262.400 4.000 2262.960 ;
    END
  END itasel[686]
  PIN itasel[687]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2265.200 4.000 2265.760 ;
    END
  END itasel[687]
  PIN itasel[688]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2268.000 4.000 2268.560 ;
    END
  END itasel[688]
  PIN itasel[689]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2270.800 4.000 2271.360 ;
    END
  END itasel[689]
  PIN itasel[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 240.800 320.000 241.360 ;
    END
  END itasel[68]
  PIN itasel[690]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2273.600 4.000 2274.160 ;
    END
  END itasel[690]
  PIN itasel[691]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2276.400 4.000 2276.960 ;
    END
  END itasel[691]
  PIN itasel[692]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2279.200 4.000 2279.760 ;
    END
  END itasel[692]
  PIN itasel[693]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2282.000 4.000 2282.560 ;
    END
  END itasel[693]
  PIN itasel[694]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2284.800 4.000 2285.360 ;
    END
  END itasel[694]
  PIN itasel[695]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2287.600 4.000 2288.160 ;
    END
  END itasel[695]
  PIN itasel[696]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2290.400 4.000 2290.960 ;
    END
  END itasel[696]
  PIN itasel[697]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2293.200 4.000 2293.760 ;
    END
  END itasel[697]
  PIN itasel[698]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2296.000 4.000 2296.560 ;
    END
  END itasel[698]
  PIN itasel[699]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2298.800 4.000 2299.360 ;
    END
  END itasel[699]
  PIN itasel[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 243.600 320.000 244.160 ;
    END
  END itasel[69]
  PIN itasel[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 201.600 4.000 202.160 ;
    END
  END itasel[6]
  PIN itasel[700]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2301.600 4.000 2302.160 ;
    END
  END itasel[700]
  PIN itasel[701]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2304.400 4.000 2304.960 ;
    END
  END itasel[701]
  PIN itasel[702]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2307.200 4.000 2307.760 ;
    END
  END itasel[702]
  PIN itasel[703]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2310.000 4.000 2310.560 ;
    END
  END itasel[703]
  PIN itasel[704]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2312.800 4.000 2313.360 ;
    END
  END itasel[704]
  PIN itasel[705]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2315.600 4.000 2316.160 ;
    END
  END itasel[705]
  PIN itasel[706]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2318.400 4.000 2318.960 ;
    END
  END itasel[706]
  PIN itasel[707]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2321.200 4.000 2321.760 ;
    END
  END itasel[707]
  PIN itasel[708]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2324.000 4.000 2324.560 ;
    END
  END itasel[708]
  PIN itasel[709]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2326.800 4.000 2327.360 ;
    END
  END itasel[709]
  PIN itasel[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 246.400 320.000 246.960 ;
    END
  END itasel[70]
  PIN itasel[710]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2329.600 4.000 2330.160 ;
    END
  END itasel[710]
  PIN itasel[711]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2332.400 4.000 2332.960 ;
    END
  END itasel[711]
  PIN itasel[712]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2335.200 4.000 2335.760 ;
    END
  END itasel[712]
  PIN itasel[713]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2338.000 4.000 2338.560 ;
    END
  END itasel[713]
  PIN itasel[714]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2340.800 4.000 2341.360 ;
    END
  END itasel[714]
  PIN itasel[715]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2343.600 4.000 2344.160 ;
    END
  END itasel[715]
  PIN itasel[716]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2346.400 4.000 2346.960 ;
    END
  END itasel[716]
  PIN itasel[717]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2349.200 4.000 2349.760 ;
    END
  END itasel[717]
  PIN itasel[718]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2352.000 4.000 2352.560 ;
    END
  END itasel[718]
  PIN itasel[719]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2354.800 4.000 2355.360 ;
    END
  END itasel[719]
  PIN itasel[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 249.200 320.000 249.760 ;
    END
  END itasel[71]
  PIN itasel[720]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2223.200 320.000 2223.760 ;
    END
  END itasel[720]
  PIN itasel[721]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2226.000 320.000 2226.560 ;
    END
  END itasel[721]
  PIN itasel[722]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2228.800 320.000 2229.360 ;
    END
  END itasel[722]
  PIN itasel[723]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2231.600 320.000 2232.160 ;
    END
  END itasel[723]
  PIN itasel[724]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2234.400 320.000 2234.960 ;
    END
  END itasel[724]
  PIN itasel[725]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2237.200 320.000 2237.760 ;
    END
  END itasel[725]
  PIN itasel[726]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2240.000 320.000 2240.560 ;
    END
  END itasel[726]
  PIN itasel[727]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2242.800 320.000 2243.360 ;
    END
  END itasel[727]
  PIN itasel[728]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2245.600 320.000 2246.160 ;
    END
  END itasel[728]
  PIN itasel[729]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2248.400 320.000 2248.960 ;
    END
  END itasel[729]
  PIN itasel[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 252.000 320.000 252.560 ;
    END
  END itasel[72]
  PIN itasel[730]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2251.200 320.000 2251.760 ;
    END
  END itasel[730]
  PIN itasel[731]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2254.000 320.000 2254.560 ;
    END
  END itasel[731]
  PIN itasel[732]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2256.800 320.000 2257.360 ;
    END
  END itasel[732]
  PIN itasel[733]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2259.600 320.000 2260.160 ;
    END
  END itasel[733]
  PIN itasel[734]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2262.400 320.000 2262.960 ;
    END
  END itasel[734]
  PIN itasel[735]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2265.200 320.000 2265.760 ;
    END
  END itasel[735]
  PIN itasel[736]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2268.000 320.000 2268.560 ;
    END
  END itasel[736]
  PIN itasel[737]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2270.800 320.000 2271.360 ;
    END
  END itasel[737]
  PIN itasel[738]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2273.600 320.000 2274.160 ;
    END
  END itasel[738]
  PIN itasel[739]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2276.400 320.000 2276.960 ;
    END
  END itasel[739]
  PIN itasel[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 254.800 320.000 255.360 ;
    END
  END itasel[73]
  PIN itasel[740]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2279.200 320.000 2279.760 ;
    END
  END itasel[740]
  PIN itasel[741]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2282.000 320.000 2282.560 ;
    END
  END itasel[741]
  PIN itasel[742]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2284.800 320.000 2285.360 ;
    END
  END itasel[742]
  PIN itasel[743]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2287.600 320.000 2288.160 ;
    END
  END itasel[743]
  PIN itasel[744]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2290.400 320.000 2290.960 ;
    END
  END itasel[744]
  PIN itasel[745]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2293.200 320.000 2293.760 ;
    END
  END itasel[745]
  PIN itasel[746]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2296.000 320.000 2296.560 ;
    END
  END itasel[746]
  PIN itasel[747]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2298.800 320.000 2299.360 ;
    END
  END itasel[747]
  PIN itasel[748]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2301.600 320.000 2302.160 ;
    END
  END itasel[748]
  PIN itasel[749]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2304.400 320.000 2304.960 ;
    END
  END itasel[749]
  PIN itasel[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 257.600 320.000 258.160 ;
    END
  END itasel[74]
  PIN itasel[750]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2307.200 320.000 2307.760 ;
    END
  END itasel[750]
  PIN itasel[751]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2310.000 320.000 2310.560 ;
    END
  END itasel[751]
  PIN itasel[752]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2312.800 320.000 2313.360 ;
    END
  END itasel[752]
  PIN itasel[753]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2315.600 320.000 2316.160 ;
    END
  END itasel[753]
  PIN itasel[754]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2318.400 320.000 2318.960 ;
    END
  END itasel[754]
  PIN itasel[755]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2321.200 320.000 2321.760 ;
    END
  END itasel[755]
  PIN itasel[756]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2324.000 320.000 2324.560 ;
    END
  END itasel[756]
  PIN itasel[757]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2326.800 320.000 2327.360 ;
    END
  END itasel[757]
  PIN itasel[758]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2329.600 320.000 2330.160 ;
    END
  END itasel[758]
  PIN itasel[759]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2332.400 320.000 2332.960 ;
    END
  END itasel[759]
  PIN itasel[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 260.400 320.000 260.960 ;
    END
  END itasel[75]
  PIN itasel[760]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2335.200 320.000 2335.760 ;
    END
  END itasel[760]
  PIN itasel[761]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2338.000 320.000 2338.560 ;
    END
  END itasel[761]
  PIN itasel[762]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2340.800 320.000 2341.360 ;
    END
  END itasel[762]
  PIN itasel[763]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2343.600 320.000 2344.160 ;
    END
  END itasel[763]
  PIN itasel[764]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2346.400 320.000 2346.960 ;
    END
  END itasel[764]
  PIN itasel[765]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2349.200 320.000 2349.760 ;
    END
  END itasel[765]
  PIN itasel[766]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2352.000 320.000 2352.560 ;
    END
  END itasel[766]
  PIN itasel[767]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 2354.800 320.000 2355.360 ;
    END
  END itasel[767]
  PIN itasel[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 263.200 320.000 263.760 ;
    END
  END itasel[76]
  PIN itasel[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 266.000 320.000 266.560 ;
    END
  END itasel[77]
  PIN itasel[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 268.800 320.000 269.360 ;
    END
  END itasel[78]
  PIN itasel[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 271.600 320.000 272.160 ;
    END
  END itasel[79]
  PIN itasel[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 204.400 4.000 204.960 ;
    END
  END itasel[7]
  PIN itasel[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 274.400 320.000 274.960 ;
    END
  END itasel[80]
  PIN itasel[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 277.200 320.000 277.760 ;
    END
  END itasel[81]
  PIN itasel[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 280.000 320.000 280.560 ;
    END
  END itasel[82]
  PIN itasel[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 282.800 320.000 283.360 ;
    END
  END itasel[83]
  PIN itasel[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 285.600 320.000 286.160 ;
    END
  END itasel[84]
  PIN itasel[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 288.400 320.000 288.960 ;
    END
  END itasel[85]
  PIN itasel[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 291.200 320.000 291.760 ;
    END
  END itasel[86]
  PIN itasel[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 294.000 320.000 294.560 ;
    END
  END itasel[87]
  PIN itasel[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 296.800 320.000 297.360 ;
    END
  END itasel[88]
  PIN itasel[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 299.600 320.000 300.160 ;
    END
  END itasel[89]
  PIN itasel[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 207.200 4.000 207.760 ;
    END
  END itasel[8]
  PIN itasel[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 302.400 320.000 302.960 ;
    END
  END itasel[90]
  PIN itasel[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 305.200 320.000 305.760 ;
    END
  END itasel[91]
  PIN itasel[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 308.000 320.000 308.560 ;
    END
  END itasel[92]
  PIN itasel[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 310.800 320.000 311.360 ;
    END
  END itasel[93]
  PIN itasel[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 313.600 320.000 314.160 ;
    END
  END itasel[94]
  PIN itasel[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 316.400 320.000 316.960 ;
    END
  END itasel[95]
  PIN itasel[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 476.000 4.000 476.560 ;
    END
  END itasel[96]
  PIN itasel[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 478.800 4.000 479.360 ;
    END
  END itasel[97]
  PIN itasel[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 481.600 4.000 482.160 ;
    END
  END itasel[98]
  PIN itasel[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 484.400 4.000 484.960 ;
    END
  END itasel[99]
  PIN itasel[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 210.000 4.000 210.560 ;
    END
  END itasel[9]
  PIN nsel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 5.600 2698.000 6.160 2702.000 ;
    END
  END nsel[0]
  PIN nsel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 11.200 2698.000 11.760 2702.000 ;
    END
  END nsel[1]
  PIN nsel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 16.800 2698.000 17.360 2702.000 ;
    END
  END nsel[2]
  PIN nsel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 22.400 2698.000 22.960 2702.000 ;
    END
  END nsel[3]
  PIN nsel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 28.000 2698.000 28.560 2702.000 ;
    END
  END nsel[4]
  PIN nsel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 33.600 2698.000 34.160 2702.000 ;
    END
  END nsel[5]
  PIN segm[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 31.360 0.000 31.920 4.000 ;
    END
  END segm[0]
  PIN segm[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 244.160 0.000 244.720 4.000 ;
    END
  END segm[10]
  PIN segm[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 265.440 0.000 266.000 4.000 ;
    END
  END segm[11]
  PIN segm[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 286.720 0.000 287.280 4.000 ;
    END
  END segm[12]
  PIN segm[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 308.000 0.000 308.560 4.000 ;
    END
  END segm[13]
  PIN segm[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 52.640 0.000 53.200 4.000 ;
    END
  END segm[1]
  PIN segm[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 73.920 0.000 74.480 4.000 ;
    END
  END segm[2]
  PIN segm[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 95.200 0.000 95.760 4.000 ;
    END
  END segm[3]
  PIN segm[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 116.480 0.000 117.040 4.000 ;
    END
  END segm[4]
  PIN segm[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 137.760 0.000 138.320 4.000 ;
    END
  END segm[5]
  PIN segm[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 159.040 0.000 159.600 4.000 ;
    END
  END segm[6]
  PIN segm[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 180.320 0.000 180.880 4.000 ;
    END
  END segm[7]
  PIN segm[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 201.600 0.000 202.160 4.000 ;
    END
  END segm[8]
  PIN segm[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 222.880 0.000 223.440 4.000 ;
    END
  END segm[9]
  PIN sel[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 39.200 2698.000 39.760 2702.000 ;
    END
  END sel[0]
  PIN sel[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 95.200 2698.000 95.760 2702.000 ;
    END
  END sel[10]
  PIN sel[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 100.800 2698.000 101.360 2702.000 ;
    END
  END sel[11]
  PIN sel[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 44.800 2698.000 45.360 2702.000 ;
    END
  END sel[1]
  PIN sel[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 50.400 2698.000 50.960 2702.000 ;
    END
  END sel[2]
  PIN sel[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 56.000 2698.000 56.560 2702.000 ;
    END
  END sel[3]
  PIN sel[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 61.600 2698.000 62.160 2702.000 ;
    END
  END sel[4]
  PIN sel[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 67.200 2698.000 67.760 2702.000 ;
    END
  END sel[5]
  PIN sel[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 72.800 2698.000 73.360 2702.000 ;
    END
  END sel[6]
  PIN sel[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 78.400 2698.000 78.960 2702.000 ;
    END
  END sel[7]
  PIN sel[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 84.000 2698.000 84.560 2702.000 ;
    END
  END sel[8]
  PIN sel[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 89.600 2698.000 90.160 2702.000 ;
    END
  END sel[9]
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 2685.500 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 2685.500 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 2685.500 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 2685.500 ;
    END
  END vss
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 313.040 2686.170 ;
      LAYER Metal2 ;
        RECT 2.380 2697.700 5.300 2698.500 ;
        RECT 6.460 2697.700 10.900 2698.500 ;
        RECT 12.060 2697.700 16.500 2698.500 ;
        RECT 17.660 2697.700 22.100 2698.500 ;
        RECT 23.260 2697.700 27.700 2698.500 ;
        RECT 28.860 2697.700 33.300 2698.500 ;
        RECT 34.460 2697.700 38.900 2698.500 ;
        RECT 40.060 2697.700 44.500 2698.500 ;
        RECT 45.660 2697.700 50.100 2698.500 ;
        RECT 51.260 2697.700 55.700 2698.500 ;
        RECT 56.860 2697.700 61.300 2698.500 ;
        RECT 62.460 2697.700 66.900 2698.500 ;
        RECT 68.060 2697.700 72.500 2698.500 ;
        RECT 73.660 2697.700 78.100 2698.500 ;
        RECT 79.260 2697.700 83.700 2698.500 ;
        RECT 84.860 2697.700 89.300 2698.500 ;
        RECT 90.460 2697.700 94.900 2698.500 ;
        RECT 96.060 2697.700 100.500 2698.500 ;
        RECT 101.660 2697.700 106.100 2698.500 ;
        RECT 107.260 2697.700 111.700 2698.500 ;
        RECT 112.860 2697.700 117.300 2698.500 ;
        RECT 118.460 2697.700 122.900 2698.500 ;
        RECT 124.060 2697.700 128.500 2698.500 ;
        RECT 129.660 2697.700 134.100 2698.500 ;
        RECT 135.260 2697.700 139.700 2698.500 ;
        RECT 140.860 2697.700 145.300 2698.500 ;
        RECT 146.460 2697.700 150.900 2698.500 ;
        RECT 152.060 2697.700 156.500 2698.500 ;
        RECT 157.660 2697.700 162.100 2698.500 ;
        RECT 163.260 2697.700 167.700 2698.500 ;
        RECT 168.860 2697.700 173.300 2698.500 ;
        RECT 174.460 2697.700 178.900 2698.500 ;
        RECT 180.060 2697.700 184.500 2698.500 ;
        RECT 185.660 2697.700 190.100 2698.500 ;
        RECT 191.260 2697.700 195.700 2698.500 ;
        RECT 196.860 2697.700 201.300 2698.500 ;
        RECT 202.460 2697.700 206.900 2698.500 ;
        RECT 208.060 2697.700 212.500 2698.500 ;
        RECT 213.660 2697.700 218.100 2698.500 ;
        RECT 219.260 2697.700 223.700 2698.500 ;
        RECT 224.860 2697.700 229.300 2698.500 ;
        RECT 230.460 2697.700 234.900 2698.500 ;
        RECT 236.060 2697.700 240.500 2698.500 ;
        RECT 241.660 2697.700 246.100 2698.500 ;
        RECT 247.260 2697.700 251.700 2698.500 ;
        RECT 252.860 2697.700 257.300 2698.500 ;
        RECT 258.460 2697.700 262.900 2698.500 ;
        RECT 264.060 2697.700 268.500 2698.500 ;
        RECT 269.660 2697.700 274.100 2698.500 ;
        RECT 275.260 2697.700 279.700 2698.500 ;
        RECT 280.860 2697.700 285.300 2698.500 ;
        RECT 286.460 2697.700 290.900 2698.500 ;
        RECT 292.060 2697.700 296.500 2698.500 ;
        RECT 297.660 2697.700 302.100 2698.500 ;
        RECT 303.260 2697.700 307.700 2698.500 ;
        RECT 308.860 2697.700 313.300 2698.500 ;
        RECT 314.460 2697.700 317.940 2698.500 ;
        RECT 2.380 4.300 317.940 2697.700 ;
        RECT 2.380 3.500 9.780 4.300 ;
        RECT 10.940 3.500 31.060 4.300 ;
        RECT 32.220 3.500 52.340 4.300 ;
        RECT 53.500 3.500 73.620 4.300 ;
        RECT 74.780 3.500 94.900 4.300 ;
        RECT 96.060 3.500 116.180 4.300 ;
        RECT 117.340 3.500 137.460 4.300 ;
        RECT 138.620 3.500 158.740 4.300 ;
        RECT 159.900 3.500 180.020 4.300 ;
        RECT 181.180 3.500 201.300 4.300 ;
        RECT 202.460 3.500 222.580 4.300 ;
        RECT 223.740 3.500 243.860 4.300 ;
        RECT 245.020 3.500 265.140 4.300 ;
        RECT 266.300 3.500 286.420 4.300 ;
        RECT 287.580 3.500 307.700 4.300 ;
        RECT 308.860 3.500 317.940 4.300 ;
      LAYER Metal3 ;
        RECT 2.330 2512.460 317.990 2685.340 ;
        RECT 4.300 2511.300 315.700 2512.460 ;
        RECT 2.330 2509.660 317.990 2511.300 ;
        RECT 4.300 2508.500 315.700 2509.660 ;
        RECT 2.330 2506.860 317.990 2508.500 ;
        RECT 4.300 2505.700 315.700 2506.860 ;
        RECT 2.330 2504.060 317.990 2505.700 ;
        RECT 4.300 2502.900 315.700 2504.060 ;
        RECT 2.330 2501.260 317.990 2502.900 ;
        RECT 4.300 2500.100 315.700 2501.260 ;
        RECT 2.330 2498.460 317.990 2500.100 ;
        RECT 4.300 2497.300 315.700 2498.460 ;
        RECT 2.330 2495.660 317.990 2497.300 ;
        RECT 4.300 2494.500 315.700 2495.660 ;
        RECT 2.330 2492.860 317.990 2494.500 ;
        RECT 4.300 2491.700 315.700 2492.860 ;
        RECT 2.330 2490.060 317.990 2491.700 ;
        RECT 4.300 2488.900 315.700 2490.060 ;
        RECT 2.330 2487.260 317.990 2488.900 ;
        RECT 4.300 2486.100 315.700 2487.260 ;
        RECT 2.330 2484.460 317.990 2486.100 ;
        RECT 4.300 2483.300 315.700 2484.460 ;
        RECT 2.330 2481.660 317.990 2483.300 ;
        RECT 4.300 2480.500 315.700 2481.660 ;
        RECT 2.330 2478.860 317.990 2480.500 ;
        RECT 4.300 2477.700 315.700 2478.860 ;
        RECT 2.330 2476.060 317.990 2477.700 ;
        RECT 4.300 2474.900 315.700 2476.060 ;
        RECT 2.330 2473.260 317.990 2474.900 ;
        RECT 4.300 2472.100 315.700 2473.260 ;
        RECT 2.330 2470.460 317.990 2472.100 ;
        RECT 4.300 2469.300 315.700 2470.460 ;
        RECT 2.330 2467.660 317.990 2469.300 ;
        RECT 4.300 2466.500 315.700 2467.660 ;
        RECT 2.330 2464.860 317.990 2466.500 ;
        RECT 4.300 2463.700 315.700 2464.860 ;
        RECT 2.330 2462.060 317.990 2463.700 ;
        RECT 4.300 2460.900 315.700 2462.060 ;
        RECT 2.330 2459.260 317.990 2460.900 ;
        RECT 4.300 2458.100 315.700 2459.260 ;
        RECT 2.330 2456.460 317.990 2458.100 ;
        RECT 4.300 2455.300 315.700 2456.460 ;
        RECT 2.330 2453.660 317.990 2455.300 ;
        RECT 4.300 2452.500 315.700 2453.660 ;
        RECT 2.330 2450.860 317.990 2452.500 ;
        RECT 4.300 2449.700 315.700 2450.860 ;
        RECT 2.330 2448.060 317.990 2449.700 ;
        RECT 4.300 2446.900 315.700 2448.060 ;
        RECT 2.330 2445.260 317.990 2446.900 ;
        RECT 4.300 2444.100 315.700 2445.260 ;
        RECT 2.330 2442.460 317.990 2444.100 ;
        RECT 4.300 2441.300 315.700 2442.460 ;
        RECT 2.330 2439.660 317.990 2441.300 ;
        RECT 4.300 2438.500 315.700 2439.660 ;
        RECT 2.330 2436.860 317.990 2438.500 ;
        RECT 4.300 2435.700 315.700 2436.860 ;
        RECT 2.330 2434.060 317.990 2435.700 ;
        RECT 4.300 2432.900 315.700 2434.060 ;
        RECT 2.330 2431.260 317.990 2432.900 ;
        RECT 4.300 2430.100 315.700 2431.260 ;
        RECT 2.330 2428.460 317.990 2430.100 ;
        RECT 4.300 2427.300 315.700 2428.460 ;
        RECT 2.330 2425.660 317.990 2427.300 ;
        RECT 4.300 2424.500 315.700 2425.660 ;
        RECT 2.330 2422.860 317.990 2424.500 ;
        RECT 4.300 2421.700 315.700 2422.860 ;
        RECT 2.330 2420.060 317.990 2421.700 ;
        RECT 4.300 2418.900 315.700 2420.060 ;
        RECT 2.330 2417.260 317.990 2418.900 ;
        RECT 4.300 2416.100 315.700 2417.260 ;
        RECT 2.330 2414.460 317.990 2416.100 ;
        RECT 4.300 2413.300 315.700 2414.460 ;
        RECT 2.330 2411.660 317.990 2413.300 ;
        RECT 4.300 2410.500 315.700 2411.660 ;
        RECT 2.330 2408.860 317.990 2410.500 ;
        RECT 4.300 2407.700 315.700 2408.860 ;
        RECT 2.330 2406.060 317.990 2407.700 ;
        RECT 4.300 2404.900 315.700 2406.060 ;
        RECT 2.330 2403.260 317.990 2404.900 ;
        RECT 4.300 2402.100 315.700 2403.260 ;
        RECT 2.330 2400.460 317.990 2402.100 ;
        RECT 4.300 2399.300 315.700 2400.460 ;
        RECT 2.330 2397.660 317.990 2399.300 ;
        RECT 4.300 2396.500 315.700 2397.660 ;
        RECT 2.330 2394.860 317.990 2396.500 ;
        RECT 4.300 2393.700 315.700 2394.860 ;
        RECT 2.330 2392.060 317.990 2393.700 ;
        RECT 4.300 2390.900 315.700 2392.060 ;
        RECT 2.330 2389.260 317.990 2390.900 ;
        RECT 4.300 2388.100 315.700 2389.260 ;
        RECT 2.330 2386.460 317.990 2388.100 ;
        RECT 4.300 2385.300 315.700 2386.460 ;
        RECT 2.330 2383.660 317.990 2385.300 ;
        RECT 4.300 2382.500 315.700 2383.660 ;
        RECT 2.330 2380.860 317.990 2382.500 ;
        RECT 4.300 2379.700 315.700 2380.860 ;
        RECT 2.330 2378.060 317.990 2379.700 ;
        RECT 4.300 2376.900 315.700 2378.060 ;
        RECT 2.330 2375.260 317.990 2376.900 ;
        RECT 4.300 2374.100 315.700 2375.260 ;
        RECT 2.330 2372.460 317.990 2374.100 ;
        RECT 4.300 2371.300 315.700 2372.460 ;
        RECT 2.330 2369.660 317.990 2371.300 ;
        RECT 4.300 2368.500 315.700 2369.660 ;
        RECT 2.330 2366.860 317.990 2368.500 ;
        RECT 4.300 2365.700 315.700 2366.860 ;
        RECT 2.330 2364.060 317.990 2365.700 ;
        RECT 4.300 2362.900 315.700 2364.060 ;
        RECT 2.330 2361.260 317.990 2362.900 ;
        RECT 4.300 2360.100 315.700 2361.260 ;
        RECT 2.330 2358.460 317.990 2360.100 ;
        RECT 4.300 2357.300 315.700 2358.460 ;
        RECT 2.330 2355.660 317.990 2357.300 ;
        RECT 4.300 2354.500 315.700 2355.660 ;
        RECT 2.330 2352.860 317.990 2354.500 ;
        RECT 4.300 2351.700 315.700 2352.860 ;
        RECT 2.330 2350.060 317.990 2351.700 ;
        RECT 4.300 2348.900 315.700 2350.060 ;
        RECT 2.330 2347.260 317.990 2348.900 ;
        RECT 4.300 2346.100 315.700 2347.260 ;
        RECT 2.330 2344.460 317.990 2346.100 ;
        RECT 4.300 2343.300 315.700 2344.460 ;
        RECT 2.330 2341.660 317.990 2343.300 ;
        RECT 4.300 2340.500 315.700 2341.660 ;
        RECT 2.330 2338.860 317.990 2340.500 ;
        RECT 4.300 2337.700 315.700 2338.860 ;
        RECT 2.330 2336.060 317.990 2337.700 ;
        RECT 4.300 2334.900 315.700 2336.060 ;
        RECT 2.330 2333.260 317.990 2334.900 ;
        RECT 4.300 2332.100 315.700 2333.260 ;
        RECT 2.330 2330.460 317.990 2332.100 ;
        RECT 4.300 2329.300 315.700 2330.460 ;
        RECT 2.330 2327.660 317.990 2329.300 ;
        RECT 4.300 2326.500 315.700 2327.660 ;
        RECT 2.330 2324.860 317.990 2326.500 ;
        RECT 4.300 2323.700 315.700 2324.860 ;
        RECT 2.330 2322.060 317.990 2323.700 ;
        RECT 4.300 2320.900 315.700 2322.060 ;
        RECT 2.330 2319.260 317.990 2320.900 ;
        RECT 4.300 2318.100 315.700 2319.260 ;
        RECT 2.330 2316.460 317.990 2318.100 ;
        RECT 4.300 2315.300 315.700 2316.460 ;
        RECT 2.330 2313.660 317.990 2315.300 ;
        RECT 4.300 2312.500 315.700 2313.660 ;
        RECT 2.330 2310.860 317.990 2312.500 ;
        RECT 4.300 2309.700 315.700 2310.860 ;
        RECT 2.330 2308.060 317.990 2309.700 ;
        RECT 4.300 2306.900 315.700 2308.060 ;
        RECT 2.330 2305.260 317.990 2306.900 ;
        RECT 4.300 2304.100 315.700 2305.260 ;
        RECT 2.330 2302.460 317.990 2304.100 ;
        RECT 4.300 2301.300 315.700 2302.460 ;
        RECT 2.330 2299.660 317.990 2301.300 ;
        RECT 4.300 2298.500 315.700 2299.660 ;
        RECT 2.330 2296.860 317.990 2298.500 ;
        RECT 4.300 2295.700 315.700 2296.860 ;
        RECT 2.330 2294.060 317.990 2295.700 ;
        RECT 4.300 2292.900 315.700 2294.060 ;
        RECT 2.330 2291.260 317.990 2292.900 ;
        RECT 4.300 2290.100 315.700 2291.260 ;
        RECT 2.330 2288.460 317.990 2290.100 ;
        RECT 4.300 2287.300 315.700 2288.460 ;
        RECT 2.330 2285.660 317.990 2287.300 ;
        RECT 4.300 2284.500 315.700 2285.660 ;
        RECT 2.330 2282.860 317.990 2284.500 ;
        RECT 4.300 2281.700 315.700 2282.860 ;
        RECT 2.330 2280.060 317.990 2281.700 ;
        RECT 4.300 2278.900 315.700 2280.060 ;
        RECT 2.330 2277.260 317.990 2278.900 ;
        RECT 4.300 2276.100 315.700 2277.260 ;
        RECT 2.330 2274.460 317.990 2276.100 ;
        RECT 4.300 2273.300 315.700 2274.460 ;
        RECT 2.330 2271.660 317.990 2273.300 ;
        RECT 4.300 2270.500 315.700 2271.660 ;
        RECT 2.330 2268.860 317.990 2270.500 ;
        RECT 4.300 2267.700 315.700 2268.860 ;
        RECT 2.330 2266.060 317.990 2267.700 ;
        RECT 4.300 2264.900 315.700 2266.060 ;
        RECT 2.330 2263.260 317.990 2264.900 ;
        RECT 4.300 2262.100 315.700 2263.260 ;
        RECT 2.330 2260.460 317.990 2262.100 ;
        RECT 4.300 2259.300 315.700 2260.460 ;
        RECT 2.330 2257.660 317.990 2259.300 ;
        RECT 4.300 2256.500 315.700 2257.660 ;
        RECT 2.330 2254.860 317.990 2256.500 ;
        RECT 4.300 2253.700 315.700 2254.860 ;
        RECT 2.330 2252.060 317.990 2253.700 ;
        RECT 4.300 2250.900 315.700 2252.060 ;
        RECT 2.330 2249.260 317.990 2250.900 ;
        RECT 4.300 2248.100 315.700 2249.260 ;
        RECT 2.330 2246.460 317.990 2248.100 ;
        RECT 4.300 2245.300 315.700 2246.460 ;
        RECT 2.330 2243.660 317.990 2245.300 ;
        RECT 4.300 2242.500 315.700 2243.660 ;
        RECT 2.330 2240.860 317.990 2242.500 ;
        RECT 4.300 2239.700 315.700 2240.860 ;
        RECT 2.330 2238.060 317.990 2239.700 ;
        RECT 4.300 2236.900 315.700 2238.060 ;
        RECT 2.330 2235.260 317.990 2236.900 ;
        RECT 4.300 2234.100 315.700 2235.260 ;
        RECT 2.330 2232.460 317.990 2234.100 ;
        RECT 4.300 2231.300 315.700 2232.460 ;
        RECT 2.330 2229.660 317.990 2231.300 ;
        RECT 4.300 2228.500 315.700 2229.660 ;
        RECT 2.330 2226.860 317.990 2228.500 ;
        RECT 4.300 2225.700 315.700 2226.860 ;
        RECT 2.330 2224.060 317.990 2225.700 ;
        RECT 4.300 2222.900 315.700 2224.060 ;
        RECT 2.330 2221.260 317.990 2222.900 ;
        RECT 4.300 2220.100 315.700 2221.260 ;
        RECT 2.330 2218.460 317.990 2220.100 ;
        RECT 4.300 2217.300 315.700 2218.460 ;
        RECT 2.330 2215.660 317.990 2217.300 ;
        RECT 4.300 2214.500 315.700 2215.660 ;
        RECT 2.330 2212.860 317.990 2214.500 ;
        RECT 4.300 2211.700 315.700 2212.860 ;
        RECT 2.330 2210.060 317.990 2211.700 ;
        RECT 4.300 2208.900 315.700 2210.060 ;
        RECT 2.330 2207.260 317.990 2208.900 ;
        RECT 4.300 2206.100 315.700 2207.260 ;
        RECT 2.330 2204.460 317.990 2206.100 ;
        RECT 4.300 2203.300 315.700 2204.460 ;
        RECT 2.330 2201.660 317.990 2203.300 ;
        RECT 4.300 2200.500 315.700 2201.660 ;
        RECT 2.330 2198.860 317.990 2200.500 ;
        RECT 4.300 2197.700 315.700 2198.860 ;
        RECT 2.330 2196.060 317.990 2197.700 ;
        RECT 4.300 2194.900 315.700 2196.060 ;
        RECT 2.330 2193.260 317.990 2194.900 ;
        RECT 4.300 2192.100 315.700 2193.260 ;
        RECT 2.330 2190.460 317.990 2192.100 ;
        RECT 4.300 2189.300 315.700 2190.460 ;
        RECT 2.330 2187.660 317.990 2189.300 ;
        RECT 4.300 2186.500 315.700 2187.660 ;
        RECT 2.330 2184.860 317.990 2186.500 ;
        RECT 4.300 2183.700 315.700 2184.860 ;
        RECT 2.330 2182.060 317.990 2183.700 ;
        RECT 4.300 2180.900 315.700 2182.060 ;
        RECT 2.330 2179.260 317.990 2180.900 ;
        RECT 4.300 2178.100 315.700 2179.260 ;
        RECT 2.330 2176.460 317.990 2178.100 ;
        RECT 4.300 2175.300 315.700 2176.460 ;
        RECT 2.330 2173.660 317.990 2175.300 ;
        RECT 4.300 2172.500 315.700 2173.660 ;
        RECT 2.330 2170.860 317.990 2172.500 ;
        RECT 4.300 2169.700 315.700 2170.860 ;
        RECT 2.330 2168.060 317.990 2169.700 ;
        RECT 4.300 2166.900 315.700 2168.060 ;
        RECT 2.330 2165.260 317.990 2166.900 ;
        RECT 4.300 2164.100 315.700 2165.260 ;
        RECT 2.330 2162.460 317.990 2164.100 ;
        RECT 4.300 2161.300 315.700 2162.460 ;
        RECT 2.330 2159.660 317.990 2161.300 ;
        RECT 4.300 2158.500 315.700 2159.660 ;
        RECT 2.330 2156.860 317.990 2158.500 ;
        RECT 4.300 2155.700 315.700 2156.860 ;
        RECT 2.330 2154.060 317.990 2155.700 ;
        RECT 4.300 2152.900 315.700 2154.060 ;
        RECT 2.330 2151.260 317.990 2152.900 ;
        RECT 4.300 2150.100 315.700 2151.260 ;
        RECT 2.330 2148.460 317.990 2150.100 ;
        RECT 4.300 2147.300 315.700 2148.460 ;
        RECT 2.330 2145.660 317.990 2147.300 ;
        RECT 4.300 2144.500 315.700 2145.660 ;
        RECT 2.330 2142.860 317.990 2144.500 ;
        RECT 4.300 2141.700 315.700 2142.860 ;
        RECT 2.330 2140.060 317.990 2141.700 ;
        RECT 4.300 2138.900 315.700 2140.060 ;
        RECT 2.330 2137.260 317.990 2138.900 ;
        RECT 4.300 2136.100 315.700 2137.260 ;
        RECT 2.330 2134.460 317.990 2136.100 ;
        RECT 4.300 2133.300 315.700 2134.460 ;
        RECT 2.330 2131.660 317.990 2133.300 ;
        RECT 4.300 2130.500 315.700 2131.660 ;
        RECT 2.330 2128.860 317.990 2130.500 ;
        RECT 4.300 2127.700 315.700 2128.860 ;
        RECT 2.330 2126.060 317.990 2127.700 ;
        RECT 4.300 2124.900 315.700 2126.060 ;
        RECT 2.330 2123.260 317.990 2124.900 ;
        RECT 4.300 2122.100 315.700 2123.260 ;
        RECT 2.330 2120.460 317.990 2122.100 ;
        RECT 4.300 2119.300 315.700 2120.460 ;
        RECT 2.330 2117.660 317.990 2119.300 ;
        RECT 4.300 2116.500 315.700 2117.660 ;
        RECT 2.330 2114.860 317.990 2116.500 ;
        RECT 4.300 2113.700 315.700 2114.860 ;
        RECT 2.330 2112.060 317.990 2113.700 ;
        RECT 4.300 2110.900 315.700 2112.060 ;
        RECT 2.330 2109.260 317.990 2110.900 ;
        RECT 4.300 2108.100 315.700 2109.260 ;
        RECT 2.330 2106.460 317.990 2108.100 ;
        RECT 4.300 2105.300 315.700 2106.460 ;
        RECT 2.330 2103.660 317.990 2105.300 ;
        RECT 4.300 2102.500 315.700 2103.660 ;
        RECT 2.330 2100.860 317.990 2102.500 ;
        RECT 4.300 2099.700 315.700 2100.860 ;
        RECT 2.330 2098.060 317.990 2099.700 ;
        RECT 4.300 2096.900 315.700 2098.060 ;
        RECT 2.330 2095.260 317.990 2096.900 ;
        RECT 4.300 2094.100 315.700 2095.260 ;
        RECT 2.330 2092.460 317.990 2094.100 ;
        RECT 4.300 2091.300 315.700 2092.460 ;
        RECT 2.330 2089.660 317.990 2091.300 ;
        RECT 4.300 2088.500 315.700 2089.660 ;
        RECT 2.330 2086.860 317.990 2088.500 ;
        RECT 4.300 2085.700 315.700 2086.860 ;
        RECT 2.330 2084.060 317.990 2085.700 ;
        RECT 4.300 2082.900 315.700 2084.060 ;
        RECT 2.330 2081.260 317.990 2082.900 ;
        RECT 4.300 2080.100 315.700 2081.260 ;
        RECT 2.330 2078.460 317.990 2080.100 ;
        RECT 4.300 2077.300 315.700 2078.460 ;
        RECT 2.330 2075.660 317.990 2077.300 ;
        RECT 4.300 2074.500 315.700 2075.660 ;
        RECT 2.330 2072.860 317.990 2074.500 ;
        RECT 4.300 2071.700 315.700 2072.860 ;
        RECT 2.330 2070.060 317.990 2071.700 ;
        RECT 4.300 2068.900 315.700 2070.060 ;
        RECT 2.330 2067.260 317.990 2068.900 ;
        RECT 4.300 2066.100 315.700 2067.260 ;
        RECT 2.330 2064.460 317.990 2066.100 ;
        RECT 4.300 2063.300 315.700 2064.460 ;
        RECT 2.330 2061.660 317.990 2063.300 ;
        RECT 4.300 2060.500 315.700 2061.660 ;
        RECT 2.330 2058.860 317.990 2060.500 ;
        RECT 4.300 2057.700 315.700 2058.860 ;
        RECT 2.330 2056.060 317.990 2057.700 ;
        RECT 4.300 2054.900 315.700 2056.060 ;
        RECT 2.330 2053.260 317.990 2054.900 ;
        RECT 4.300 2052.100 315.700 2053.260 ;
        RECT 2.330 2050.460 317.990 2052.100 ;
        RECT 4.300 2049.300 315.700 2050.460 ;
        RECT 2.330 2047.660 317.990 2049.300 ;
        RECT 4.300 2046.500 315.700 2047.660 ;
        RECT 2.330 2044.860 317.990 2046.500 ;
        RECT 4.300 2043.700 315.700 2044.860 ;
        RECT 2.330 2042.060 317.990 2043.700 ;
        RECT 4.300 2040.900 315.700 2042.060 ;
        RECT 2.330 2039.260 317.990 2040.900 ;
        RECT 4.300 2038.100 315.700 2039.260 ;
        RECT 2.330 2036.460 317.990 2038.100 ;
        RECT 4.300 2035.300 315.700 2036.460 ;
        RECT 2.330 2033.660 317.990 2035.300 ;
        RECT 4.300 2032.500 315.700 2033.660 ;
        RECT 2.330 2030.860 317.990 2032.500 ;
        RECT 4.300 2029.700 315.700 2030.860 ;
        RECT 2.330 2028.060 317.990 2029.700 ;
        RECT 4.300 2026.900 315.700 2028.060 ;
        RECT 2.330 2025.260 317.990 2026.900 ;
        RECT 4.300 2024.100 315.700 2025.260 ;
        RECT 2.330 2022.460 317.990 2024.100 ;
        RECT 4.300 2021.300 315.700 2022.460 ;
        RECT 2.330 2019.660 317.990 2021.300 ;
        RECT 4.300 2018.500 315.700 2019.660 ;
        RECT 2.330 2016.860 317.990 2018.500 ;
        RECT 4.300 2015.700 315.700 2016.860 ;
        RECT 2.330 2014.060 317.990 2015.700 ;
        RECT 4.300 2012.900 315.700 2014.060 ;
        RECT 2.330 2011.260 317.990 2012.900 ;
        RECT 4.300 2010.100 315.700 2011.260 ;
        RECT 2.330 2008.460 317.990 2010.100 ;
        RECT 4.300 2007.300 315.700 2008.460 ;
        RECT 2.330 2005.660 317.990 2007.300 ;
        RECT 4.300 2004.500 315.700 2005.660 ;
        RECT 2.330 2002.860 317.990 2004.500 ;
        RECT 4.300 2001.700 315.700 2002.860 ;
        RECT 2.330 2000.060 317.990 2001.700 ;
        RECT 4.300 1998.900 315.700 2000.060 ;
        RECT 2.330 1997.260 317.990 1998.900 ;
        RECT 4.300 1996.100 315.700 1997.260 ;
        RECT 2.330 1994.460 317.990 1996.100 ;
        RECT 4.300 1993.300 315.700 1994.460 ;
        RECT 2.330 1991.660 317.990 1993.300 ;
        RECT 4.300 1990.500 315.700 1991.660 ;
        RECT 2.330 1988.860 317.990 1990.500 ;
        RECT 4.300 1987.700 315.700 1988.860 ;
        RECT 2.330 1986.060 317.990 1987.700 ;
        RECT 4.300 1984.900 315.700 1986.060 ;
        RECT 2.330 1983.260 317.990 1984.900 ;
        RECT 4.300 1982.100 315.700 1983.260 ;
        RECT 2.330 1980.460 317.990 1982.100 ;
        RECT 4.300 1979.300 315.700 1980.460 ;
        RECT 2.330 1977.660 317.990 1979.300 ;
        RECT 4.300 1976.500 315.700 1977.660 ;
        RECT 2.330 1974.860 317.990 1976.500 ;
        RECT 4.300 1973.700 315.700 1974.860 ;
        RECT 2.330 1972.060 317.990 1973.700 ;
        RECT 4.300 1970.900 315.700 1972.060 ;
        RECT 2.330 1969.260 317.990 1970.900 ;
        RECT 4.300 1968.100 315.700 1969.260 ;
        RECT 2.330 1966.460 317.990 1968.100 ;
        RECT 4.300 1965.300 315.700 1966.460 ;
        RECT 2.330 1963.660 317.990 1965.300 ;
        RECT 4.300 1962.500 315.700 1963.660 ;
        RECT 2.330 1960.860 317.990 1962.500 ;
        RECT 4.300 1959.700 315.700 1960.860 ;
        RECT 2.330 1958.060 317.990 1959.700 ;
        RECT 4.300 1956.900 315.700 1958.060 ;
        RECT 2.330 1955.260 317.990 1956.900 ;
        RECT 4.300 1954.100 315.700 1955.260 ;
        RECT 2.330 1952.460 317.990 1954.100 ;
        RECT 4.300 1951.300 315.700 1952.460 ;
        RECT 2.330 1949.660 317.990 1951.300 ;
        RECT 4.300 1948.500 315.700 1949.660 ;
        RECT 2.330 1946.860 317.990 1948.500 ;
        RECT 4.300 1945.700 315.700 1946.860 ;
        RECT 2.330 1944.060 317.990 1945.700 ;
        RECT 4.300 1942.900 315.700 1944.060 ;
        RECT 2.330 1941.260 317.990 1942.900 ;
        RECT 4.300 1940.100 315.700 1941.260 ;
        RECT 2.330 1938.460 317.990 1940.100 ;
        RECT 4.300 1937.300 315.700 1938.460 ;
        RECT 2.330 1935.660 317.990 1937.300 ;
        RECT 4.300 1934.500 315.700 1935.660 ;
        RECT 2.330 1932.860 317.990 1934.500 ;
        RECT 4.300 1931.700 315.700 1932.860 ;
        RECT 2.330 1930.060 317.990 1931.700 ;
        RECT 4.300 1928.900 315.700 1930.060 ;
        RECT 2.330 1927.260 317.990 1928.900 ;
        RECT 4.300 1926.100 315.700 1927.260 ;
        RECT 2.330 1924.460 317.990 1926.100 ;
        RECT 4.300 1923.300 315.700 1924.460 ;
        RECT 2.330 1921.660 317.990 1923.300 ;
        RECT 4.300 1920.500 315.700 1921.660 ;
        RECT 2.330 1918.860 317.990 1920.500 ;
        RECT 4.300 1917.700 315.700 1918.860 ;
        RECT 2.330 1916.060 317.990 1917.700 ;
        RECT 4.300 1914.900 315.700 1916.060 ;
        RECT 2.330 1913.260 317.990 1914.900 ;
        RECT 4.300 1912.100 315.700 1913.260 ;
        RECT 2.330 1910.460 317.990 1912.100 ;
        RECT 4.300 1909.300 315.700 1910.460 ;
        RECT 2.330 1907.660 317.990 1909.300 ;
        RECT 4.300 1906.500 315.700 1907.660 ;
        RECT 2.330 1904.860 317.990 1906.500 ;
        RECT 4.300 1903.700 315.700 1904.860 ;
        RECT 2.330 1902.060 317.990 1903.700 ;
        RECT 4.300 1900.900 315.700 1902.060 ;
        RECT 2.330 1899.260 317.990 1900.900 ;
        RECT 4.300 1898.100 315.700 1899.260 ;
        RECT 2.330 1896.460 317.990 1898.100 ;
        RECT 4.300 1895.300 315.700 1896.460 ;
        RECT 2.330 1893.660 317.990 1895.300 ;
        RECT 4.300 1892.500 315.700 1893.660 ;
        RECT 2.330 1890.860 317.990 1892.500 ;
        RECT 4.300 1889.700 315.700 1890.860 ;
        RECT 2.330 1888.060 317.990 1889.700 ;
        RECT 4.300 1886.900 315.700 1888.060 ;
        RECT 2.330 1885.260 317.990 1886.900 ;
        RECT 4.300 1884.100 315.700 1885.260 ;
        RECT 2.330 1882.460 317.990 1884.100 ;
        RECT 4.300 1881.300 315.700 1882.460 ;
        RECT 2.330 1879.660 317.990 1881.300 ;
        RECT 4.300 1878.500 315.700 1879.660 ;
        RECT 2.330 1876.860 317.990 1878.500 ;
        RECT 4.300 1875.700 315.700 1876.860 ;
        RECT 2.330 1874.060 317.990 1875.700 ;
        RECT 4.300 1872.900 315.700 1874.060 ;
        RECT 2.330 1871.260 317.990 1872.900 ;
        RECT 4.300 1870.100 315.700 1871.260 ;
        RECT 2.330 1868.460 317.990 1870.100 ;
        RECT 4.300 1867.300 315.700 1868.460 ;
        RECT 2.330 1865.660 317.990 1867.300 ;
        RECT 4.300 1864.500 315.700 1865.660 ;
        RECT 2.330 1862.860 317.990 1864.500 ;
        RECT 4.300 1861.700 315.700 1862.860 ;
        RECT 2.330 1860.060 317.990 1861.700 ;
        RECT 4.300 1858.900 315.700 1860.060 ;
        RECT 2.330 1857.260 317.990 1858.900 ;
        RECT 4.300 1856.100 315.700 1857.260 ;
        RECT 2.330 1854.460 317.990 1856.100 ;
        RECT 4.300 1853.300 315.700 1854.460 ;
        RECT 2.330 1851.660 317.990 1853.300 ;
        RECT 4.300 1850.500 315.700 1851.660 ;
        RECT 2.330 1848.860 317.990 1850.500 ;
        RECT 4.300 1847.700 315.700 1848.860 ;
        RECT 2.330 1846.060 317.990 1847.700 ;
        RECT 4.300 1844.900 315.700 1846.060 ;
        RECT 2.330 1843.260 317.990 1844.900 ;
        RECT 4.300 1842.100 315.700 1843.260 ;
        RECT 2.330 1840.460 317.990 1842.100 ;
        RECT 4.300 1839.300 315.700 1840.460 ;
        RECT 2.330 1837.660 317.990 1839.300 ;
        RECT 4.300 1836.500 315.700 1837.660 ;
        RECT 2.330 1834.860 317.990 1836.500 ;
        RECT 4.300 1833.700 315.700 1834.860 ;
        RECT 2.330 1832.060 317.990 1833.700 ;
        RECT 4.300 1830.900 315.700 1832.060 ;
        RECT 2.330 1829.260 317.990 1830.900 ;
        RECT 4.300 1828.100 315.700 1829.260 ;
        RECT 2.330 1826.460 317.990 1828.100 ;
        RECT 4.300 1825.300 315.700 1826.460 ;
        RECT 2.330 1823.660 317.990 1825.300 ;
        RECT 4.300 1822.500 315.700 1823.660 ;
        RECT 2.330 1820.860 317.990 1822.500 ;
        RECT 4.300 1819.700 315.700 1820.860 ;
        RECT 2.330 1818.060 317.990 1819.700 ;
        RECT 4.300 1816.900 315.700 1818.060 ;
        RECT 2.330 1815.260 317.990 1816.900 ;
        RECT 4.300 1814.100 315.700 1815.260 ;
        RECT 2.330 1812.460 317.990 1814.100 ;
        RECT 4.300 1811.300 315.700 1812.460 ;
        RECT 2.330 1809.660 317.990 1811.300 ;
        RECT 4.300 1808.500 315.700 1809.660 ;
        RECT 2.330 1806.860 317.990 1808.500 ;
        RECT 4.300 1805.700 315.700 1806.860 ;
        RECT 2.330 1804.060 317.990 1805.700 ;
        RECT 4.300 1802.900 315.700 1804.060 ;
        RECT 2.330 1801.260 317.990 1802.900 ;
        RECT 4.300 1800.100 315.700 1801.260 ;
        RECT 2.330 1798.460 317.990 1800.100 ;
        RECT 4.300 1797.300 315.700 1798.460 ;
        RECT 2.330 1795.660 317.990 1797.300 ;
        RECT 4.300 1794.500 315.700 1795.660 ;
        RECT 2.330 1792.860 317.990 1794.500 ;
        RECT 4.300 1791.700 315.700 1792.860 ;
        RECT 2.330 1790.060 317.990 1791.700 ;
        RECT 4.300 1788.900 315.700 1790.060 ;
        RECT 2.330 1787.260 317.990 1788.900 ;
        RECT 4.300 1786.100 315.700 1787.260 ;
        RECT 2.330 1784.460 317.990 1786.100 ;
        RECT 4.300 1783.300 315.700 1784.460 ;
        RECT 2.330 1781.660 317.990 1783.300 ;
        RECT 4.300 1780.500 315.700 1781.660 ;
        RECT 2.330 1778.860 317.990 1780.500 ;
        RECT 4.300 1777.700 315.700 1778.860 ;
        RECT 2.330 1776.060 317.990 1777.700 ;
        RECT 4.300 1774.900 315.700 1776.060 ;
        RECT 2.330 1773.260 317.990 1774.900 ;
        RECT 4.300 1772.100 315.700 1773.260 ;
        RECT 2.330 1770.460 317.990 1772.100 ;
        RECT 4.300 1769.300 315.700 1770.460 ;
        RECT 2.330 1767.660 317.990 1769.300 ;
        RECT 4.300 1766.500 315.700 1767.660 ;
        RECT 2.330 1764.860 317.990 1766.500 ;
        RECT 4.300 1763.700 315.700 1764.860 ;
        RECT 2.330 1762.060 317.990 1763.700 ;
        RECT 4.300 1760.900 315.700 1762.060 ;
        RECT 2.330 1759.260 317.990 1760.900 ;
        RECT 4.300 1758.100 315.700 1759.260 ;
        RECT 2.330 1756.460 317.990 1758.100 ;
        RECT 4.300 1755.300 315.700 1756.460 ;
        RECT 2.330 1753.660 317.990 1755.300 ;
        RECT 4.300 1752.500 315.700 1753.660 ;
        RECT 2.330 1750.860 317.990 1752.500 ;
        RECT 4.300 1749.700 315.700 1750.860 ;
        RECT 2.330 1748.060 317.990 1749.700 ;
        RECT 4.300 1746.900 315.700 1748.060 ;
        RECT 2.330 1745.260 317.990 1746.900 ;
        RECT 4.300 1744.100 315.700 1745.260 ;
        RECT 2.330 1742.460 317.990 1744.100 ;
        RECT 4.300 1741.300 315.700 1742.460 ;
        RECT 2.330 1739.660 317.990 1741.300 ;
        RECT 4.300 1738.500 315.700 1739.660 ;
        RECT 2.330 1736.860 317.990 1738.500 ;
        RECT 4.300 1735.700 315.700 1736.860 ;
        RECT 2.330 1734.060 317.990 1735.700 ;
        RECT 4.300 1732.900 315.700 1734.060 ;
        RECT 2.330 1731.260 317.990 1732.900 ;
        RECT 4.300 1730.100 315.700 1731.260 ;
        RECT 2.330 1728.460 317.990 1730.100 ;
        RECT 4.300 1727.300 315.700 1728.460 ;
        RECT 2.330 1725.660 317.990 1727.300 ;
        RECT 4.300 1724.500 315.700 1725.660 ;
        RECT 2.330 1722.860 317.990 1724.500 ;
        RECT 4.300 1721.700 315.700 1722.860 ;
        RECT 2.330 1720.060 317.990 1721.700 ;
        RECT 4.300 1718.900 315.700 1720.060 ;
        RECT 2.330 1717.260 317.990 1718.900 ;
        RECT 4.300 1716.100 315.700 1717.260 ;
        RECT 2.330 1714.460 317.990 1716.100 ;
        RECT 4.300 1713.300 315.700 1714.460 ;
        RECT 2.330 1711.660 317.990 1713.300 ;
        RECT 4.300 1710.500 315.700 1711.660 ;
        RECT 2.330 1708.860 317.990 1710.500 ;
        RECT 4.300 1707.700 315.700 1708.860 ;
        RECT 2.330 1706.060 317.990 1707.700 ;
        RECT 4.300 1704.900 315.700 1706.060 ;
        RECT 2.330 1703.260 317.990 1704.900 ;
        RECT 4.300 1702.100 315.700 1703.260 ;
        RECT 2.330 1700.460 317.990 1702.100 ;
        RECT 4.300 1699.300 315.700 1700.460 ;
        RECT 2.330 1697.660 317.990 1699.300 ;
        RECT 4.300 1696.500 315.700 1697.660 ;
        RECT 2.330 1694.860 317.990 1696.500 ;
        RECT 4.300 1693.700 315.700 1694.860 ;
        RECT 2.330 1692.060 317.990 1693.700 ;
        RECT 4.300 1690.900 315.700 1692.060 ;
        RECT 2.330 1689.260 317.990 1690.900 ;
        RECT 4.300 1688.100 315.700 1689.260 ;
        RECT 2.330 1686.460 317.990 1688.100 ;
        RECT 4.300 1685.300 315.700 1686.460 ;
        RECT 2.330 1683.660 317.990 1685.300 ;
        RECT 4.300 1682.500 315.700 1683.660 ;
        RECT 2.330 1680.860 317.990 1682.500 ;
        RECT 4.300 1679.700 315.700 1680.860 ;
        RECT 2.330 1678.060 317.990 1679.700 ;
        RECT 4.300 1676.900 315.700 1678.060 ;
        RECT 2.330 1675.260 317.990 1676.900 ;
        RECT 4.300 1674.100 315.700 1675.260 ;
        RECT 2.330 1672.460 317.990 1674.100 ;
        RECT 4.300 1671.300 315.700 1672.460 ;
        RECT 2.330 1669.660 317.990 1671.300 ;
        RECT 4.300 1668.500 315.700 1669.660 ;
        RECT 2.330 1666.860 317.990 1668.500 ;
        RECT 4.300 1665.700 315.700 1666.860 ;
        RECT 2.330 1664.060 317.990 1665.700 ;
        RECT 4.300 1662.900 315.700 1664.060 ;
        RECT 2.330 1661.260 317.990 1662.900 ;
        RECT 4.300 1660.100 315.700 1661.260 ;
        RECT 2.330 1658.460 317.990 1660.100 ;
        RECT 4.300 1657.300 315.700 1658.460 ;
        RECT 2.330 1655.660 317.990 1657.300 ;
        RECT 4.300 1654.500 315.700 1655.660 ;
        RECT 2.330 1652.860 317.990 1654.500 ;
        RECT 4.300 1651.700 315.700 1652.860 ;
        RECT 2.330 1650.060 317.990 1651.700 ;
        RECT 4.300 1648.900 315.700 1650.060 ;
        RECT 2.330 1647.260 317.990 1648.900 ;
        RECT 4.300 1646.100 315.700 1647.260 ;
        RECT 2.330 1644.460 317.990 1646.100 ;
        RECT 4.300 1643.300 315.700 1644.460 ;
        RECT 2.330 1641.660 317.990 1643.300 ;
        RECT 4.300 1640.500 315.700 1641.660 ;
        RECT 2.330 1638.860 317.990 1640.500 ;
        RECT 4.300 1637.700 315.700 1638.860 ;
        RECT 2.330 1636.060 317.990 1637.700 ;
        RECT 4.300 1634.900 315.700 1636.060 ;
        RECT 2.330 1633.260 317.990 1634.900 ;
        RECT 4.300 1632.100 315.700 1633.260 ;
        RECT 2.330 1630.460 317.990 1632.100 ;
        RECT 4.300 1629.300 315.700 1630.460 ;
        RECT 2.330 1627.660 317.990 1629.300 ;
        RECT 4.300 1626.500 315.700 1627.660 ;
        RECT 2.330 1624.860 317.990 1626.500 ;
        RECT 4.300 1623.700 315.700 1624.860 ;
        RECT 2.330 1622.060 317.990 1623.700 ;
        RECT 4.300 1620.900 315.700 1622.060 ;
        RECT 2.330 1619.260 317.990 1620.900 ;
        RECT 4.300 1618.100 315.700 1619.260 ;
        RECT 2.330 1616.460 317.990 1618.100 ;
        RECT 4.300 1615.300 315.700 1616.460 ;
        RECT 2.330 1613.660 317.990 1615.300 ;
        RECT 4.300 1612.500 315.700 1613.660 ;
        RECT 2.330 1610.860 317.990 1612.500 ;
        RECT 4.300 1609.700 315.700 1610.860 ;
        RECT 2.330 1608.060 317.990 1609.700 ;
        RECT 4.300 1606.900 315.700 1608.060 ;
        RECT 2.330 1605.260 317.990 1606.900 ;
        RECT 4.300 1604.100 315.700 1605.260 ;
        RECT 2.330 1602.460 317.990 1604.100 ;
        RECT 4.300 1601.300 315.700 1602.460 ;
        RECT 2.330 1599.660 317.990 1601.300 ;
        RECT 4.300 1598.500 315.700 1599.660 ;
        RECT 2.330 1596.860 317.990 1598.500 ;
        RECT 4.300 1595.700 315.700 1596.860 ;
        RECT 2.330 1594.060 317.990 1595.700 ;
        RECT 4.300 1592.900 315.700 1594.060 ;
        RECT 2.330 1591.260 317.990 1592.900 ;
        RECT 4.300 1590.100 315.700 1591.260 ;
        RECT 2.330 1588.460 317.990 1590.100 ;
        RECT 4.300 1587.300 315.700 1588.460 ;
        RECT 2.330 1585.660 317.990 1587.300 ;
        RECT 4.300 1584.500 315.700 1585.660 ;
        RECT 2.330 1582.860 317.990 1584.500 ;
        RECT 4.300 1581.700 315.700 1582.860 ;
        RECT 2.330 1580.060 317.990 1581.700 ;
        RECT 4.300 1578.900 315.700 1580.060 ;
        RECT 2.330 1577.260 317.990 1578.900 ;
        RECT 4.300 1576.100 315.700 1577.260 ;
        RECT 2.330 1574.460 317.990 1576.100 ;
        RECT 4.300 1573.300 315.700 1574.460 ;
        RECT 2.330 1571.660 317.990 1573.300 ;
        RECT 4.300 1570.500 315.700 1571.660 ;
        RECT 2.330 1568.860 317.990 1570.500 ;
        RECT 4.300 1567.700 315.700 1568.860 ;
        RECT 2.330 1566.060 317.990 1567.700 ;
        RECT 4.300 1564.900 315.700 1566.060 ;
        RECT 2.330 1563.260 317.990 1564.900 ;
        RECT 4.300 1562.100 315.700 1563.260 ;
        RECT 2.330 1560.460 317.990 1562.100 ;
        RECT 4.300 1559.300 315.700 1560.460 ;
        RECT 2.330 1557.660 317.990 1559.300 ;
        RECT 4.300 1556.500 315.700 1557.660 ;
        RECT 2.330 1554.860 317.990 1556.500 ;
        RECT 4.300 1553.700 315.700 1554.860 ;
        RECT 2.330 1552.060 317.990 1553.700 ;
        RECT 4.300 1550.900 315.700 1552.060 ;
        RECT 2.330 1549.260 317.990 1550.900 ;
        RECT 4.300 1548.100 315.700 1549.260 ;
        RECT 2.330 1546.460 317.990 1548.100 ;
        RECT 4.300 1545.300 315.700 1546.460 ;
        RECT 2.330 1543.660 317.990 1545.300 ;
        RECT 4.300 1542.500 315.700 1543.660 ;
        RECT 2.330 1540.860 317.990 1542.500 ;
        RECT 4.300 1539.700 315.700 1540.860 ;
        RECT 2.330 1538.060 317.990 1539.700 ;
        RECT 4.300 1536.900 315.700 1538.060 ;
        RECT 2.330 1535.260 317.990 1536.900 ;
        RECT 4.300 1534.100 315.700 1535.260 ;
        RECT 2.330 1532.460 317.990 1534.100 ;
        RECT 4.300 1531.300 315.700 1532.460 ;
        RECT 2.330 1529.660 317.990 1531.300 ;
        RECT 4.300 1528.500 315.700 1529.660 ;
        RECT 2.330 1526.860 317.990 1528.500 ;
        RECT 4.300 1525.700 315.700 1526.860 ;
        RECT 2.330 1524.060 317.990 1525.700 ;
        RECT 4.300 1522.900 315.700 1524.060 ;
        RECT 2.330 1521.260 317.990 1522.900 ;
        RECT 4.300 1520.100 315.700 1521.260 ;
        RECT 2.330 1518.460 317.990 1520.100 ;
        RECT 4.300 1517.300 315.700 1518.460 ;
        RECT 2.330 1515.660 317.990 1517.300 ;
        RECT 4.300 1514.500 315.700 1515.660 ;
        RECT 2.330 1512.860 317.990 1514.500 ;
        RECT 4.300 1511.700 315.700 1512.860 ;
        RECT 2.330 1510.060 317.990 1511.700 ;
        RECT 4.300 1508.900 315.700 1510.060 ;
        RECT 2.330 1507.260 317.990 1508.900 ;
        RECT 4.300 1506.100 315.700 1507.260 ;
        RECT 2.330 1504.460 317.990 1506.100 ;
        RECT 4.300 1503.300 315.700 1504.460 ;
        RECT 2.330 1501.660 317.990 1503.300 ;
        RECT 4.300 1500.500 315.700 1501.660 ;
        RECT 2.330 1498.860 317.990 1500.500 ;
        RECT 4.300 1497.700 315.700 1498.860 ;
        RECT 2.330 1496.060 317.990 1497.700 ;
        RECT 4.300 1494.900 315.700 1496.060 ;
        RECT 2.330 1493.260 317.990 1494.900 ;
        RECT 4.300 1492.100 315.700 1493.260 ;
        RECT 2.330 1490.460 317.990 1492.100 ;
        RECT 4.300 1489.300 315.700 1490.460 ;
        RECT 2.330 1487.660 317.990 1489.300 ;
        RECT 4.300 1486.500 315.700 1487.660 ;
        RECT 2.330 1484.860 317.990 1486.500 ;
        RECT 4.300 1483.700 315.700 1484.860 ;
        RECT 2.330 1482.060 317.990 1483.700 ;
        RECT 4.300 1480.900 315.700 1482.060 ;
        RECT 2.330 1479.260 317.990 1480.900 ;
        RECT 4.300 1478.100 315.700 1479.260 ;
        RECT 2.330 1476.460 317.990 1478.100 ;
        RECT 4.300 1475.300 315.700 1476.460 ;
        RECT 2.330 1473.660 317.990 1475.300 ;
        RECT 4.300 1472.500 315.700 1473.660 ;
        RECT 2.330 1470.860 317.990 1472.500 ;
        RECT 4.300 1469.700 315.700 1470.860 ;
        RECT 2.330 1468.060 317.990 1469.700 ;
        RECT 4.300 1466.900 315.700 1468.060 ;
        RECT 2.330 1465.260 317.990 1466.900 ;
        RECT 4.300 1464.100 315.700 1465.260 ;
        RECT 2.330 1462.460 317.990 1464.100 ;
        RECT 4.300 1461.300 315.700 1462.460 ;
        RECT 2.330 1459.660 317.990 1461.300 ;
        RECT 4.300 1458.500 315.700 1459.660 ;
        RECT 2.330 1456.860 317.990 1458.500 ;
        RECT 4.300 1455.700 315.700 1456.860 ;
        RECT 2.330 1454.060 317.990 1455.700 ;
        RECT 4.300 1452.900 315.700 1454.060 ;
        RECT 2.330 1451.260 317.990 1452.900 ;
        RECT 4.300 1450.100 315.700 1451.260 ;
        RECT 2.330 1448.460 317.990 1450.100 ;
        RECT 4.300 1447.300 315.700 1448.460 ;
        RECT 2.330 1445.660 317.990 1447.300 ;
        RECT 4.300 1444.500 315.700 1445.660 ;
        RECT 2.330 1442.860 317.990 1444.500 ;
        RECT 4.300 1441.700 315.700 1442.860 ;
        RECT 2.330 1440.060 317.990 1441.700 ;
        RECT 4.300 1438.900 315.700 1440.060 ;
        RECT 2.330 1437.260 317.990 1438.900 ;
        RECT 4.300 1436.100 315.700 1437.260 ;
        RECT 2.330 1434.460 317.990 1436.100 ;
        RECT 4.300 1433.300 315.700 1434.460 ;
        RECT 2.330 1431.660 317.990 1433.300 ;
        RECT 4.300 1430.500 315.700 1431.660 ;
        RECT 2.330 1428.860 317.990 1430.500 ;
        RECT 4.300 1427.700 315.700 1428.860 ;
        RECT 2.330 1426.060 317.990 1427.700 ;
        RECT 4.300 1424.900 315.700 1426.060 ;
        RECT 2.330 1423.260 317.990 1424.900 ;
        RECT 4.300 1422.100 315.700 1423.260 ;
        RECT 2.330 1420.460 317.990 1422.100 ;
        RECT 4.300 1419.300 315.700 1420.460 ;
        RECT 2.330 1417.660 317.990 1419.300 ;
        RECT 4.300 1416.500 315.700 1417.660 ;
        RECT 2.330 1414.860 317.990 1416.500 ;
        RECT 4.300 1413.700 315.700 1414.860 ;
        RECT 2.330 1412.060 317.990 1413.700 ;
        RECT 4.300 1410.900 315.700 1412.060 ;
        RECT 2.330 1409.260 317.990 1410.900 ;
        RECT 4.300 1408.100 315.700 1409.260 ;
        RECT 2.330 1406.460 317.990 1408.100 ;
        RECT 4.300 1405.300 315.700 1406.460 ;
        RECT 2.330 1403.660 317.990 1405.300 ;
        RECT 4.300 1402.500 315.700 1403.660 ;
        RECT 2.330 1400.860 317.990 1402.500 ;
        RECT 4.300 1399.700 315.700 1400.860 ;
        RECT 2.330 1398.060 317.990 1399.700 ;
        RECT 4.300 1396.900 315.700 1398.060 ;
        RECT 2.330 1395.260 317.990 1396.900 ;
        RECT 4.300 1394.100 315.700 1395.260 ;
        RECT 2.330 1392.460 317.990 1394.100 ;
        RECT 4.300 1391.300 315.700 1392.460 ;
        RECT 2.330 1389.660 317.990 1391.300 ;
        RECT 4.300 1388.500 315.700 1389.660 ;
        RECT 2.330 1386.860 317.990 1388.500 ;
        RECT 4.300 1385.700 315.700 1386.860 ;
        RECT 2.330 1384.060 317.990 1385.700 ;
        RECT 4.300 1382.900 315.700 1384.060 ;
        RECT 2.330 1381.260 317.990 1382.900 ;
        RECT 4.300 1380.100 315.700 1381.260 ;
        RECT 2.330 1378.460 317.990 1380.100 ;
        RECT 4.300 1377.300 315.700 1378.460 ;
        RECT 2.330 1375.660 317.990 1377.300 ;
        RECT 4.300 1374.500 315.700 1375.660 ;
        RECT 2.330 1372.860 317.990 1374.500 ;
        RECT 4.300 1371.700 315.700 1372.860 ;
        RECT 2.330 1370.060 317.990 1371.700 ;
        RECT 4.300 1368.900 315.700 1370.060 ;
        RECT 2.330 1367.260 317.990 1368.900 ;
        RECT 4.300 1366.100 315.700 1367.260 ;
        RECT 2.330 1364.460 317.990 1366.100 ;
        RECT 4.300 1363.300 315.700 1364.460 ;
        RECT 2.330 1361.660 317.990 1363.300 ;
        RECT 4.300 1360.500 315.700 1361.660 ;
        RECT 2.330 1358.860 317.990 1360.500 ;
        RECT 4.300 1357.700 315.700 1358.860 ;
        RECT 2.330 1356.060 317.990 1357.700 ;
        RECT 4.300 1354.900 315.700 1356.060 ;
        RECT 2.330 1353.260 317.990 1354.900 ;
        RECT 4.300 1352.100 315.700 1353.260 ;
        RECT 2.330 1350.460 317.990 1352.100 ;
        RECT 4.300 1349.300 315.700 1350.460 ;
        RECT 2.330 1347.660 317.990 1349.300 ;
        RECT 4.300 1346.500 315.700 1347.660 ;
        RECT 2.330 1344.860 317.990 1346.500 ;
        RECT 4.300 1343.700 315.700 1344.860 ;
        RECT 2.330 1342.060 317.990 1343.700 ;
        RECT 4.300 1340.900 315.700 1342.060 ;
        RECT 2.330 1339.260 317.990 1340.900 ;
        RECT 4.300 1338.100 315.700 1339.260 ;
        RECT 2.330 1336.460 317.990 1338.100 ;
        RECT 4.300 1335.300 315.700 1336.460 ;
        RECT 2.330 1333.660 317.990 1335.300 ;
        RECT 4.300 1332.500 315.700 1333.660 ;
        RECT 2.330 1330.860 317.990 1332.500 ;
        RECT 4.300 1329.700 315.700 1330.860 ;
        RECT 2.330 1328.060 317.990 1329.700 ;
        RECT 4.300 1326.900 315.700 1328.060 ;
        RECT 2.330 1325.260 317.990 1326.900 ;
        RECT 4.300 1324.100 315.700 1325.260 ;
        RECT 2.330 1322.460 317.990 1324.100 ;
        RECT 4.300 1321.300 315.700 1322.460 ;
        RECT 2.330 1319.660 317.990 1321.300 ;
        RECT 4.300 1318.500 315.700 1319.660 ;
        RECT 2.330 1316.860 317.990 1318.500 ;
        RECT 4.300 1315.700 315.700 1316.860 ;
        RECT 2.330 1314.060 317.990 1315.700 ;
        RECT 4.300 1312.900 315.700 1314.060 ;
        RECT 2.330 1311.260 317.990 1312.900 ;
        RECT 4.300 1310.100 315.700 1311.260 ;
        RECT 2.330 1308.460 317.990 1310.100 ;
        RECT 4.300 1307.300 315.700 1308.460 ;
        RECT 2.330 1305.660 317.990 1307.300 ;
        RECT 4.300 1304.500 315.700 1305.660 ;
        RECT 2.330 1302.860 317.990 1304.500 ;
        RECT 4.300 1301.700 315.700 1302.860 ;
        RECT 2.330 1300.060 317.990 1301.700 ;
        RECT 4.300 1298.900 315.700 1300.060 ;
        RECT 2.330 1297.260 317.990 1298.900 ;
        RECT 4.300 1296.100 315.700 1297.260 ;
        RECT 2.330 1294.460 317.990 1296.100 ;
        RECT 4.300 1293.300 315.700 1294.460 ;
        RECT 2.330 1291.660 317.990 1293.300 ;
        RECT 4.300 1290.500 315.700 1291.660 ;
        RECT 2.330 1288.860 317.990 1290.500 ;
        RECT 4.300 1287.700 315.700 1288.860 ;
        RECT 2.330 1286.060 317.990 1287.700 ;
        RECT 4.300 1284.900 315.700 1286.060 ;
        RECT 2.330 1283.260 317.990 1284.900 ;
        RECT 4.300 1282.100 315.700 1283.260 ;
        RECT 2.330 1280.460 317.990 1282.100 ;
        RECT 4.300 1279.300 315.700 1280.460 ;
        RECT 2.330 1277.660 317.990 1279.300 ;
        RECT 4.300 1276.500 315.700 1277.660 ;
        RECT 2.330 1274.860 317.990 1276.500 ;
        RECT 4.300 1273.700 315.700 1274.860 ;
        RECT 2.330 1272.060 317.990 1273.700 ;
        RECT 4.300 1270.900 315.700 1272.060 ;
        RECT 2.330 1269.260 317.990 1270.900 ;
        RECT 4.300 1268.100 315.700 1269.260 ;
        RECT 2.330 1266.460 317.990 1268.100 ;
        RECT 4.300 1265.300 315.700 1266.460 ;
        RECT 2.330 1263.660 317.990 1265.300 ;
        RECT 4.300 1262.500 315.700 1263.660 ;
        RECT 2.330 1260.860 317.990 1262.500 ;
        RECT 4.300 1259.700 315.700 1260.860 ;
        RECT 2.330 1258.060 317.990 1259.700 ;
        RECT 4.300 1256.900 315.700 1258.060 ;
        RECT 2.330 1255.260 317.990 1256.900 ;
        RECT 4.300 1254.100 315.700 1255.260 ;
        RECT 2.330 1252.460 317.990 1254.100 ;
        RECT 4.300 1251.300 315.700 1252.460 ;
        RECT 2.330 1249.660 317.990 1251.300 ;
        RECT 4.300 1248.500 315.700 1249.660 ;
        RECT 2.330 1246.860 317.990 1248.500 ;
        RECT 4.300 1245.700 315.700 1246.860 ;
        RECT 2.330 1244.060 317.990 1245.700 ;
        RECT 4.300 1242.900 315.700 1244.060 ;
        RECT 2.330 1241.260 317.990 1242.900 ;
        RECT 4.300 1240.100 315.700 1241.260 ;
        RECT 2.330 1238.460 317.990 1240.100 ;
        RECT 4.300 1237.300 315.700 1238.460 ;
        RECT 2.330 1235.660 317.990 1237.300 ;
        RECT 4.300 1234.500 315.700 1235.660 ;
        RECT 2.330 1232.860 317.990 1234.500 ;
        RECT 4.300 1231.700 315.700 1232.860 ;
        RECT 2.330 1230.060 317.990 1231.700 ;
        RECT 4.300 1228.900 315.700 1230.060 ;
        RECT 2.330 1227.260 317.990 1228.900 ;
        RECT 4.300 1226.100 315.700 1227.260 ;
        RECT 2.330 1224.460 317.990 1226.100 ;
        RECT 4.300 1223.300 315.700 1224.460 ;
        RECT 2.330 1221.660 317.990 1223.300 ;
        RECT 4.300 1220.500 315.700 1221.660 ;
        RECT 2.330 1218.860 317.990 1220.500 ;
        RECT 4.300 1217.700 315.700 1218.860 ;
        RECT 2.330 1216.060 317.990 1217.700 ;
        RECT 4.300 1214.900 315.700 1216.060 ;
        RECT 2.330 1213.260 317.990 1214.900 ;
        RECT 4.300 1212.100 315.700 1213.260 ;
        RECT 2.330 1210.460 317.990 1212.100 ;
        RECT 4.300 1209.300 315.700 1210.460 ;
        RECT 2.330 1207.660 317.990 1209.300 ;
        RECT 4.300 1206.500 315.700 1207.660 ;
        RECT 2.330 1204.860 317.990 1206.500 ;
        RECT 4.300 1203.700 315.700 1204.860 ;
        RECT 2.330 1202.060 317.990 1203.700 ;
        RECT 4.300 1200.900 315.700 1202.060 ;
        RECT 2.330 1199.260 317.990 1200.900 ;
        RECT 4.300 1198.100 315.700 1199.260 ;
        RECT 2.330 1196.460 317.990 1198.100 ;
        RECT 4.300 1195.300 315.700 1196.460 ;
        RECT 2.330 1193.660 317.990 1195.300 ;
        RECT 4.300 1192.500 315.700 1193.660 ;
        RECT 2.330 1190.860 317.990 1192.500 ;
        RECT 4.300 1189.700 315.700 1190.860 ;
        RECT 2.330 1188.060 317.990 1189.700 ;
        RECT 4.300 1186.900 315.700 1188.060 ;
        RECT 2.330 1185.260 317.990 1186.900 ;
        RECT 4.300 1184.100 315.700 1185.260 ;
        RECT 2.330 1182.460 317.990 1184.100 ;
        RECT 4.300 1181.300 315.700 1182.460 ;
        RECT 2.330 1179.660 317.990 1181.300 ;
        RECT 4.300 1178.500 315.700 1179.660 ;
        RECT 2.330 1176.860 317.990 1178.500 ;
        RECT 4.300 1175.700 315.700 1176.860 ;
        RECT 2.330 1174.060 317.990 1175.700 ;
        RECT 4.300 1172.900 315.700 1174.060 ;
        RECT 2.330 1171.260 317.990 1172.900 ;
        RECT 4.300 1170.100 315.700 1171.260 ;
        RECT 2.330 1168.460 317.990 1170.100 ;
        RECT 4.300 1167.300 315.700 1168.460 ;
        RECT 2.330 1165.660 317.990 1167.300 ;
        RECT 4.300 1164.500 315.700 1165.660 ;
        RECT 2.330 1162.860 317.990 1164.500 ;
        RECT 4.300 1161.700 315.700 1162.860 ;
        RECT 2.330 1160.060 317.990 1161.700 ;
        RECT 4.300 1158.900 315.700 1160.060 ;
        RECT 2.330 1157.260 317.990 1158.900 ;
        RECT 4.300 1156.100 315.700 1157.260 ;
        RECT 2.330 1154.460 317.990 1156.100 ;
        RECT 4.300 1153.300 315.700 1154.460 ;
        RECT 2.330 1151.660 317.990 1153.300 ;
        RECT 4.300 1150.500 315.700 1151.660 ;
        RECT 2.330 1148.860 317.990 1150.500 ;
        RECT 4.300 1147.700 315.700 1148.860 ;
        RECT 2.330 1146.060 317.990 1147.700 ;
        RECT 4.300 1144.900 315.700 1146.060 ;
        RECT 2.330 1143.260 317.990 1144.900 ;
        RECT 4.300 1142.100 315.700 1143.260 ;
        RECT 2.330 1140.460 317.990 1142.100 ;
        RECT 4.300 1139.300 315.700 1140.460 ;
        RECT 2.330 1137.660 317.990 1139.300 ;
        RECT 4.300 1136.500 315.700 1137.660 ;
        RECT 2.330 1134.860 317.990 1136.500 ;
        RECT 4.300 1133.700 315.700 1134.860 ;
        RECT 2.330 1132.060 317.990 1133.700 ;
        RECT 4.300 1130.900 315.700 1132.060 ;
        RECT 2.330 1129.260 317.990 1130.900 ;
        RECT 4.300 1128.100 315.700 1129.260 ;
        RECT 2.330 1126.460 317.990 1128.100 ;
        RECT 4.300 1125.300 315.700 1126.460 ;
        RECT 2.330 1123.660 317.990 1125.300 ;
        RECT 4.300 1122.500 315.700 1123.660 ;
        RECT 2.330 1120.860 317.990 1122.500 ;
        RECT 4.300 1119.700 315.700 1120.860 ;
        RECT 2.330 1118.060 317.990 1119.700 ;
        RECT 4.300 1116.900 315.700 1118.060 ;
        RECT 2.330 1115.260 317.990 1116.900 ;
        RECT 4.300 1114.100 315.700 1115.260 ;
        RECT 2.330 1112.460 317.990 1114.100 ;
        RECT 4.300 1111.300 315.700 1112.460 ;
        RECT 2.330 1109.660 317.990 1111.300 ;
        RECT 4.300 1108.500 315.700 1109.660 ;
        RECT 2.330 1106.860 317.990 1108.500 ;
        RECT 4.300 1105.700 315.700 1106.860 ;
        RECT 2.330 1104.060 317.990 1105.700 ;
        RECT 4.300 1102.900 315.700 1104.060 ;
        RECT 2.330 1101.260 317.990 1102.900 ;
        RECT 4.300 1100.100 315.700 1101.260 ;
        RECT 2.330 1098.460 317.990 1100.100 ;
        RECT 4.300 1097.300 315.700 1098.460 ;
        RECT 2.330 1095.660 317.990 1097.300 ;
        RECT 4.300 1094.500 315.700 1095.660 ;
        RECT 2.330 1092.860 317.990 1094.500 ;
        RECT 4.300 1091.700 315.700 1092.860 ;
        RECT 2.330 1090.060 317.990 1091.700 ;
        RECT 4.300 1088.900 315.700 1090.060 ;
        RECT 2.330 1087.260 317.990 1088.900 ;
        RECT 4.300 1086.100 315.700 1087.260 ;
        RECT 2.330 1084.460 317.990 1086.100 ;
        RECT 4.300 1083.300 315.700 1084.460 ;
        RECT 2.330 1081.660 317.990 1083.300 ;
        RECT 4.300 1080.500 315.700 1081.660 ;
        RECT 2.330 1078.860 317.990 1080.500 ;
        RECT 4.300 1077.700 315.700 1078.860 ;
        RECT 2.330 1076.060 317.990 1077.700 ;
        RECT 4.300 1074.900 315.700 1076.060 ;
        RECT 2.330 1073.260 317.990 1074.900 ;
        RECT 4.300 1072.100 315.700 1073.260 ;
        RECT 2.330 1070.460 317.990 1072.100 ;
        RECT 4.300 1069.300 315.700 1070.460 ;
        RECT 2.330 1067.660 317.990 1069.300 ;
        RECT 4.300 1066.500 315.700 1067.660 ;
        RECT 2.330 1064.860 317.990 1066.500 ;
        RECT 4.300 1063.700 315.700 1064.860 ;
        RECT 2.330 1062.060 317.990 1063.700 ;
        RECT 4.300 1060.900 315.700 1062.060 ;
        RECT 2.330 1059.260 317.990 1060.900 ;
        RECT 4.300 1058.100 315.700 1059.260 ;
        RECT 2.330 1056.460 317.990 1058.100 ;
        RECT 4.300 1055.300 315.700 1056.460 ;
        RECT 2.330 1053.660 317.990 1055.300 ;
        RECT 4.300 1052.500 315.700 1053.660 ;
        RECT 2.330 1050.860 317.990 1052.500 ;
        RECT 4.300 1049.700 315.700 1050.860 ;
        RECT 2.330 1048.060 317.990 1049.700 ;
        RECT 4.300 1046.900 315.700 1048.060 ;
        RECT 2.330 1045.260 317.990 1046.900 ;
        RECT 4.300 1044.100 315.700 1045.260 ;
        RECT 2.330 1042.460 317.990 1044.100 ;
        RECT 4.300 1041.300 315.700 1042.460 ;
        RECT 2.330 1039.660 317.990 1041.300 ;
        RECT 4.300 1038.500 315.700 1039.660 ;
        RECT 2.330 1036.860 317.990 1038.500 ;
        RECT 4.300 1035.700 315.700 1036.860 ;
        RECT 2.330 1034.060 317.990 1035.700 ;
        RECT 4.300 1032.900 315.700 1034.060 ;
        RECT 2.330 1031.260 317.990 1032.900 ;
        RECT 4.300 1030.100 315.700 1031.260 ;
        RECT 2.330 1028.460 317.990 1030.100 ;
        RECT 4.300 1027.300 315.700 1028.460 ;
        RECT 2.330 1025.660 317.990 1027.300 ;
        RECT 4.300 1024.500 315.700 1025.660 ;
        RECT 2.330 1022.860 317.990 1024.500 ;
        RECT 4.300 1021.700 315.700 1022.860 ;
        RECT 2.330 1020.060 317.990 1021.700 ;
        RECT 4.300 1018.900 315.700 1020.060 ;
        RECT 2.330 1017.260 317.990 1018.900 ;
        RECT 4.300 1016.100 315.700 1017.260 ;
        RECT 2.330 1014.460 317.990 1016.100 ;
        RECT 4.300 1013.300 315.700 1014.460 ;
        RECT 2.330 1011.660 317.990 1013.300 ;
        RECT 4.300 1010.500 315.700 1011.660 ;
        RECT 2.330 1008.860 317.990 1010.500 ;
        RECT 4.300 1007.700 315.700 1008.860 ;
        RECT 2.330 1006.060 317.990 1007.700 ;
        RECT 4.300 1004.900 315.700 1006.060 ;
        RECT 2.330 1003.260 317.990 1004.900 ;
        RECT 4.300 1002.100 315.700 1003.260 ;
        RECT 2.330 1000.460 317.990 1002.100 ;
        RECT 4.300 999.300 315.700 1000.460 ;
        RECT 2.330 997.660 317.990 999.300 ;
        RECT 4.300 996.500 315.700 997.660 ;
        RECT 2.330 994.860 317.990 996.500 ;
        RECT 4.300 993.700 315.700 994.860 ;
        RECT 2.330 992.060 317.990 993.700 ;
        RECT 4.300 990.900 315.700 992.060 ;
        RECT 2.330 989.260 317.990 990.900 ;
        RECT 4.300 988.100 315.700 989.260 ;
        RECT 2.330 986.460 317.990 988.100 ;
        RECT 4.300 985.300 315.700 986.460 ;
        RECT 2.330 983.660 317.990 985.300 ;
        RECT 4.300 982.500 315.700 983.660 ;
        RECT 2.330 980.860 317.990 982.500 ;
        RECT 4.300 979.700 315.700 980.860 ;
        RECT 2.330 978.060 317.990 979.700 ;
        RECT 4.300 976.900 315.700 978.060 ;
        RECT 2.330 975.260 317.990 976.900 ;
        RECT 4.300 974.100 315.700 975.260 ;
        RECT 2.330 972.460 317.990 974.100 ;
        RECT 4.300 971.300 315.700 972.460 ;
        RECT 2.330 969.660 317.990 971.300 ;
        RECT 4.300 968.500 315.700 969.660 ;
        RECT 2.330 966.860 317.990 968.500 ;
        RECT 4.300 965.700 315.700 966.860 ;
        RECT 2.330 964.060 317.990 965.700 ;
        RECT 4.300 962.900 315.700 964.060 ;
        RECT 2.330 961.260 317.990 962.900 ;
        RECT 4.300 960.100 315.700 961.260 ;
        RECT 2.330 958.460 317.990 960.100 ;
        RECT 4.300 957.300 315.700 958.460 ;
        RECT 2.330 955.660 317.990 957.300 ;
        RECT 4.300 954.500 315.700 955.660 ;
        RECT 2.330 952.860 317.990 954.500 ;
        RECT 4.300 951.700 315.700 952.860 ;
        RECT 2.330 950.060 317.990 951.700 ;
        RECT 4.300 948.900 315.700 950.060 ;
        RECT 2.330 947.260 317.990 948.900 ;
        RECT 4.300 946.100 315.700 947.260 ;
        RECT 2.330 944.460 317.990 946.100 ;
        RECT 4.300 943.300 315.700 944.460 ;
        RECT 2.330 941.660 317.990 943.300 ;
        RECT 4.300 940.500 315.700 941.660 ;
        RECT 2.330 938.860 317.990 940.500 ;
        RECT 4.300 937.700 315.700 938.860 ;
        RECT 2.330 936.060 317.990 937.700 ;
        RECT 4.300 934.900 315.700 936.060 ;
        RECT 2.330 933.260 317.990 934.900 ;
        RECT 4.300 932.100 315.700 933.260 ;
        RECT 2.330 930.460 317.990 932.100 ;
        RECT 4.300 929.300 315.700 930.460 ;
        RECT 2.330 927.660 317.990 929.300 ;
        RECT 4.300 926.500 315.700 927.660 ;
        RECT 2.330 924.860 317.990 926.500 ;
        RECT 4.300 923.700 315.700 924.860 ;
        RECT 2.330 922.060 317.990 923.700 ;
        RECT 4.300 920.900 315.700 922.060 ;
        RECT 2.330 919.260 317.990 920.900 ;
        RECT 4.300 918.100 315.700 919.260 ;
        RECT 2.330 916.460 317.990 918.100 ;
        RECT 4.300 915.300 315.700 916.460 ;
        RECT 2.330 913.660 317.990 915.300 ;
        RECT 4.300 912.500 315.700 913.660 ;
        RECT 2.330 910.860 317.990 912.500 ;
        RECT 4.300 909.700 315.700 910.860 ;
        RECT 2.330 908.060 317.990 909.700 ;
        RECT 4.300 906.900 315.700 908.060 ;
        RECT 2.330 905.260 317.990 906.900 ;
        RECT 4.300 904.100 315.700 905.260 ;
        RECT 2.330 902.460 317.990 904.100 ;
        RECT 4.300 901.300 315.700 902.460 ;
        RECT 2.330 899.660 317.990 901.300 ;
        RECT 4.300 898.500 315.700 899.660 ;
        RECT 2.330 896.860 317.990 898.500 ;
        RECT 4.300 895.700 315.700 896.860 ;
        RECT 2.330 894.060 317.990 895.700 ;
        RECT 4.300 892.900 315.700 894.060 ;
        RECT 2.330 891.260 317.990 892.900 ;
        RECT 4.300 890.100 315.700 891.260 ;
        RECT 2.330 888.460 317.990 890.100 ;
        RECT 4.300 887.300 315.700 888.460 ;
        RECT 2.330 885.660 317.990 887.300 ;
        RECT 4.300 884.500 315.700 885.660 ;
        RECT 2.330 882.860 317.990 884.500 ;
        RECT 4.300 881.700 315.700 882.860 ;
        RECT 2.330 880.060 317.990 881.700 ;
        RECT 4.300 878.900 315.700 880.060 ;
        RECT 2.330 877.260 317.990 878.900 ;
        RECT 4.300 876.100 315.700 877.260 ;
        RECT 2.330 874.460 317.990 876.100 ;
        RECT 4.300 873.300 315.700 874.460 ;
        RECT 2.330 871.660 317.990 873.300 ;
        RECT 4.300 870.500 315.700 871.660 ;
        RECT 2.330 868.860 317.990 870.500 ;
        RECT 4.300 867.700 315.700 868.860 ;
        RECT 2.330 866.060 317.990 867.700 ;
        RECT 4.300 864.900 315.700 866.060 ;
        RECT 2.330 863.260 317.990 864.900 ;
        RECT 4.300 862.100 315.700 863.260 ;
        RECT 2.330 860.460 317.990 862.100 ;
        RECT 4.300 859.300 315.700 860.460 ;
        RECT 2.330 857.660 317.990 859.300 ;
        RECT 4.300 856.500 315.700 857.660 ;
        RECT 2.330 854.860 317.990 856.500 ;
        RECT 4.300 853.700 315.700 854.860 ;
        RECT 2.330 852.060 317.990 853.700 ;
        RECT 4.300 850.900 315.700 852.060 ;
        RECT 2.330 849.260 317.990 850.900 ;
        RECT 4.300 848.100 315.700 849.260 ;
        RECT 2.330 846.460 317.990 848.100 ;
        RECT 4.300 845.300 315.700 846.460 ;
        RECT 2.330 843.660 317.990 845.300 ;
        RECT 4.300 842.500 315.700 843.660 ;
        RECT 2.330 840.860 317.990 842.500 ;
        RECT 4.300 839.700 315.700 840.860 ;
        RECT 2.330 838.060 317.990 839.700 ;
        RECT 4.300 836.900 315.700 838.060 ;
        RECT 2.330 835.260 317.990 836.900 ;
        RECT 4.300 834.100 315.700 835.260 ;
        RECT 2.330 832.460 317.990 834.100 ;
        RECT 4.300 831.300 315.700 832.460 ;
        RECT 2.330 829.660 317.990 831.300 ;
        RECT 4.300 828.500 315.700 829.660 ;
        RECT 2.330 826.860 317.990 828.500 ;
        RECT 4.300 825.700 315.700 826.860 ;
        RECT 2.330 824.060 317.990 825.700 ;
        RECT 4.300 822.900 315.700 824.060 ;
        RECT 2.330 821.260 317.990 822.900 ;
        RECT 4.300 820.100 315.700 821.260 ;
        RECT 2.330 818.460 317.990 820.100 ;
        RECT 4.300 817.300 315.700 818.460 ;
        RECT 2.330 815.660 317.990 817.300 ;
        RECT 4.300 814.500 315.700 815.660 ;
        RECT 2.330 812.860 317.990 814.500 ;
        RECT 4.300 811.700 315.700 812.860 ;
        RECT 2.330 810.060 317.990 811.700 ;
        RECT 4.300 808.900 315.700 810.060 ;
        RECT 2.330 807.260 317.990 808.900 ;
        RECT 4.300 806.100 315.700 807.260 ;
        RECT 2.330 804.460 317.990 806.100 ;
        RECT 4.300 803.300 315.700 804.460 ;
        RECT 2.330 801.660 317.990 803.300 ;
        RECT 4.300 800.500 315.700 801.660 ;
        RECT 2.330 798.860 317.990 800.500 ;
        RECT 4.300 797.700 315.700 798.860 ;
        RECT 2.330 796.060 317.990 797.700 ;
        RECT 4.300 794.900 315.700 796.060 ;
        RECT 2.330 793.260 317.990 794.900 ;
        RECT 4.300 792.100 315.700 793.260 ;
        RECT 2.330 790.460 317.990 792.100 ;
        RECT 4.300 789.300 315.700 790.460 ;
        RECT 2.330 787.660 317.990 789.300 ;
        RECT 4.300 786.500 315.700 787.660 ;
        RECT 2.330 784.860 317.990 786.500 ;
        RECT 4.300 783.700 315.700 784.860 ;
        RECT 2.330 782.060 317.990 783.700 ;
        RECT 4.300 780.900 315.700 782.060 ;
        RECT 2.330 779.260 317.990 780.900 ;
        RECT 4.300 778.100 315.700 779.260 ;
        RECT 2.330 776.460 317.990 778.100 ;
        RECT 4.300 775.300 315.700 776.460 ;
        RECT 2.330 773.660 317.990 775.300 ;
        RECT 4.300 772.500 315.700 773.660 ;
        RECT 2.330 770.860 317.990 772.500 ;
        RECT 4.300 769.700 315.700 770.860 ;
        RECT 2.330 768.060 317.990 769.700 ;
        RECT 4.300 766.900 315.700 768.060 ;
        RECT 2.330 765.260 317.990 766.900 ;
        RECT 4.300 764.100 315.700 765.260 ;
        RECT 2.330 762.460 317.990 764.100 ;
        RECT 4.300 761.300 315.700 762.460 ;
        RECT 2.330 759.660 317.990 761.300 ;
        RECT 4.300 758.500 315.700 759.660 ;
        RECT 2.330 756.860 317.990 758.500 ;
        RECT 4.300 755.700 315.700 756.860 ;
        RECT 2.330 754.060 317.990 755.700 ;
        RECT 4.300 752.900 315.700 754.060 ;
        RECT 2.330 751.260 317.990 752.900 ;
        RECT 4.300 750.100 315.700 751.260 ;
        RECT 2.330 748.460 317.990 750.100 ;
        RECT 4.300 747.300 315.700 748.460 ;
        RECT 2.330 745.660 317.990 747.300 ;
        RECT 4.300 744.500 315.700 745.660 ;
        RECT 2.330 742.860 317.990 744.500 ;
        RECT 4.300 741.700 315.700 742.860 ;
        RECT 2.330 740.060 317.990 741.700 ;
        RECT 4.300 738.900 315.700 740.060 ;
        RECT 2.330 737.260 317.990 738.900 ;
        RECT 4.300 736.100 315.700 737.260 ;
        RECT 2.330 734.460 317.990 736.100 ;
        RECT 4.300 733.300 315.700 734.460 ;
        RECT 2.330 731.660 317.990 733.300 ;
        RECT 4.300 730.500 315.700 731.660 ;
        RECT 2.330 728.860 317.990 730.500 ;
        RECT 4.300 727.700 315.700 728.860 ;
        RECT 2.330 726.060 317.990 727.700 ;
        RECT 4.300 724.900 315.700 726.060 ;
        RECT 2.330 723.260 317.990 724.900 ;
        RECT 4.300 722.100 315.700 723.260 ;
        RECT 2.330 720.460 317.990 722.100 ;
        RECT 4.300 719.300 315.700 720.460 ;
        RECT 2.330 717.660 317.990 719.300 ;
        RECT 4.300 716.500 315.700 717.660 ;
        RECT 2.330 714.860 317.990 716.500 ;
        RECT 4.300 713.700 315.700 714.860 ;
        RECT 2.330 712.060 317.990 713.700 ;
        RECT 4.300 710.900 315.700 712.060 ;
        RECT 2.330 709.260 317.990 710.900 ;
        RECT 4.300 708.100 315.700 709.260 ;
        RECT 2.330 706.460 317.990 708.100 ;
        RECT 4.300 705.300 315.700 706.460 ;
        RECT 2.330 703.660 317.990 705.300 ;
        RECT 4.300 702.500 315.700 703.660 ;
        RECT 2.330 700.860 317.990 702.500 ;
        RECT 4.300 699.700 315.700 700.860 ;
        RECT 2.330 698.060 317.990 699.700 ;
        RECT 4.300 696.900 315.700 698.060 ;
        RECT 2.330 695.260 317.990 696.900 ;
        RECT 4.300 694.100 315.700 695.260 ;
        RECT 2.330 692.460 317.990 694.100 ;
        RECT 4.300 691.300 315.700 692.460 ;
        RECT 2.330 689.660 317.990 691.300 ;
        RECT 4.300 688.500 315.700 689.660 ;
        RECT 2.330 686.860 317.990 688.500 ;
        RECT 4.300 685.700 315.700 686.860 ;
        RECT 2.330 684.060 317.990 685.700 ;
        RECT 4.300 682.900 315.700 684.060 ;
        RECT 2.330 681.260 317.990 682.900 ;
        RECT 4.300 680.100 315.700 681.260 ;
        RECT 2.330 678.460 317.990 680.100 ;
        RECT 4.300 677.300 315.700 678.460 ;
        RECT 2.330 675.660 317.990 677.300 ;
        RECT 4.300 674.500 315.700 675.660 ;
        RECT 2.330 672.860 317.990 674.500 ;
        RECT 4.300 671.700 315.700 672.860 ;
        RECT 2.330 670.060 317.990 671.700 ;
        RECT 4.300 668.900 315.700 670.060 ;
        RECT 2.330 667.260 317.990 668.900 ;
        RECT 4.300 666.100 315.700 667.260 ;
        RECT 2.330 664.460 317.990 666.100 ;
        RECT 4.300 663.300 315.700 664.460 ;
        RECT 2.330 661.660 317.990 663.300 ;
        RECT 4.300 660.500 315.700 661.660 ;
        RECT 2.330 658.860 317.990 660.500 ;
        RECT 4.300 657.700 315.700 658.860 ;
        RECT 2.330 656.060 317.990 657.700 ;
        RECT 4.300 654.900 315.700 656.060 ;
        RECT 2.330 653.260 317.990 654.900 ;
        RECT 4.300 652.100 315.700 653.260 ;
        RECT 2.330 650.460 317.990 652.100 ;
        RECT 4.300 649.300 315.700 650.460 ;
        RECT 2.330 647.660 317.990 649.300 ;
        RECT 4.300 646.500 315.700 647.660 ;
        RECT 2.330 644.860 317.990 646.500 ;
        RECT 4.300 643.700 315.700 644.860 ;
        RECT 2.330 642.060 317.990 643.700 ;
        RECT 4.300 640.900 315.700 642.060 ;
        RECT 2.330 639.260 317.990 640.900 ;
        RECT 4.300 638.100 315.700 639.260 ;
        RECT 2.330 636.460 317.990 638.100 ;
        RECT 4.300 635.300 315.700 636.460 ;
        RECT 2.330 633.660 317.990 635.300 ;
        RECT 4.300 632.500 315.700 633.660 ;
        RECT 2.330 630.860 317.990 632.500 ;
        RECT 4.300 629.700 315.700 630.860 ;
        RECT 2.330 628.060 317.990 629.700 ;
        RECT 4.300 626.900 315.700 628.060 ;
        RECT 2.330 625.260 317.990 626.900 ;
        RECT 4.300 624.100 315.700 625.260 ;
        RECT 2.330 622.460 317.990 624.100 ;
        RECT 4.300 621.300 315.700 622.460 ;
        RECT 2.330 619.660 317.990 621.300 ;
        RECT 4.300 618.500 315.700 619.660 ;
        RECT 2.330 616.860 317.990 618.500 ;
        RECT 4.300 615.700 315.700 616.860 ;
        RECT 2.330 614.060 317.990 615.700 ;
        RECT 4.300 612.900 315.700 614.060 ;
        RECT 2.330 611.260 317.990 612.900 ;
        RECT 4.300 610.100 315.700 611.260 ;
        RECT 2.330 608.460 317.990 610.100 ;
        RECT 4.300 607.300 315.700 608.460 ;
        RECT 2.330 605.660 317.990 607.300 ;
        RECT 4.300 604.500 315.700 605.660 ;
        RECT 2.330 602.860 317.990 604.500 ;
        RECT 4.300 601.700 315.700 602.860 ;
        RECT 2.330 600.060 317.990 601.700 ;
        RECT 4.300 598.900 315.700 600.060 ;
        RECT 2.330 597.260 317.990 598.900 ;
        RECT 4.300 596.100 315.700 597.260 ;
        RECT 2.330 594.460 317.990 596.100 ;
        RECT 4.300 593.300 315.700 594.460 ;
        RECT 2.330 591.660 317.990 593.300 ;
        RECT 4.300 590.500 315.700 591.660 ;
        RECT 2.330 588.860 317.990 590.500 ;
        RECT 4.300 587.700 315.700 588.860 ;
        RECT 2.330 586.060 317.990 587.700 ;
        RECT 4.300 584.900 315.700 586.060 ;
        RECT 2.330 583.260 317.990 584.900 ;
        RECT 4.300 582.100 315.700 583.260 ;
        RECT 2.330 580.460 317.990 582.100 ;
        RECT 4.300 579.300 315.700 580.460 ;
        RECT 2.330 577.660 317.990 579.300 ;
        RECT 4.300 576.500 315.700 577.660 ;
        RECT 2.330 574.860 317.990 576.500 ;
        RECT 4.300 573.700 315.700 574.860 ;
        RECT 2.330 572.060 317.990 573.700 ;
        RECT 4.300 570.900 315.700 572.060 ;
        RECT 2.330 569.260 317.990 570.900 ;
        RECT 4.300 568.100 315.700 569.260 ;
        RECT 2.330 566.460 317.990 568.100 ;
        RECT 4.300 565.300 315.700 566.460 ;
        RECT 2.330 563.660 317.990 565.300 ;
        RECT 4.300 562.500 315.700 563.660 ;
        RECT 2.330 560.860 317.990 562.500 ;
        RECT 4.300 559.700 315.700 560.860 ;
        RECT 2.330 558.060 317.990 559.700 ;
        RECT 4.300 556.900 315.700 558.060 ;
        RECT 2.330 555.260 317.990 556.900 ;
        RECT 4.300 554.100 315.700 555.260 ;
        RECT 2.330 552.460 317.990 554.100 ;
        RECT 4.300 551.300 315.700 552.460 ;
        RECT 2.330 549.660 317.990 551.300 ;
        RECT 4.300 548.500 315.700 549.660 ;
        RECT 2.330 546.860 317.990 548.500 ;
        RECT 4.300 545.700 315.700 546.860 ;
        RECT 2.330 544.060 317.990 545.700 ;
        RECT 4.300 542.900 315.700 544.060 ;
        RECT 2.330 541.260 317.990 542.900 ;
        RECT 4.300 540.100 315.700 541.260 ;
        RECT 2.330 538.460 317.990 540.100 ;
        RECT 4.300 537.300 315.700 538.460 ;
        RECT 2.330 535.660 317.990 537.300 ;
        RECT 4.300 534.500 315.700 535.660 ;
        RECT 2.330 532.860 317.990 534.500 ;
        RECT 4.300 531.700 315.700 532.860 ;
        RECT 2.330 530.060 317.990 531.700 ;
        RECT 4.300 528.900 315.700 530.060 ;
        RECT 2.330 527.260 317.990 528.900 ;
        RECT 4.300 526.100 315.700 527.260 ;
        RECT 2.330 524.460 317.990 526.100 ;
        RECT 4.300 523.300 315.700 524.460 ;
        RECT 2.330 521.660 317.990 523.300 ;
        RECT 4.300 520.500 315.700 521.660 ;
        RECT 2.330 518.860 317.990 520.500 ;
        RECT 4.300 517.700 315.700 518.860 ;
        RECT 2.330 516.060 317.990 517.700 ;
        RECT 4.300 514.900 315.700 516.060 ;
        RECT 2.330 513.260 317.990 514.900 ;
        RECT 4.300 512.100 315.700 513.260 ;
        RECT 2.330 510.460 317.990 512.100 ;
        RECT 4.300 509.300 315.700 510.460 ;
        RECT 2.330 507.660 317.990 509.300 ;
        RECT 4.300 506.500 315.700 507.660 ;
        RECT 2.330 504.860 317.990 506.500 ;
        RECT 4.300 503.700 315.700 504.860 ;
        RECT 2.330 502.060 317.990 503.700 ;
        RECT 4.300 500.900 315.700 502.060 ;
        RECT 2.330 499.260 317.990 500.900 ;
        RECT 4.300 498.100 315.700 499.260 ;
        RECT 2.330 496.460 317.990 498.100 ;
        RECT 4.300 495.300 315.700 496.460 ;
        RECT 2.330 493.660 317.990 495.300 ;
        RECT 4.300 492.500 315.700 493.660 ;
        RECT 2.330 490.860 317.990 492.500 ;
        RECT 4.300 489.700 315.700 490.860 ;
        RECT 2.330 488.060 317.990 489.700 ;
        RECT 4.300 486.900 315.700 488.060 ;
        RECT 2.330 485.260 317.990 486.900 ;
        RECT 4.300 484.100 315.700 485.260 ;
        RECT 2.330 482.460 317.990 484.100 ;
        RECT 4.300 481.300 315.700 482.460 ;
        RECT 2.330 479.660 317.990 481.300 ;
        RECT 4.300 478.500 315.700 479.660 ;
        RECT 2.330 476.860 317.990 478.500 ;
        RECT 4.300 475.700 315.700 476.860 ;
        RECT 2.330 474.060 317.990 475.700 ;
        RECT 4.300 472.900 315.700 474.060 ;
        RECT 2.330 471.260 317.990 472.900 ;
        RECT 4.300 470.100 315.700 471.260 ;
        RECT 2.330 468.460 317.990 470.100 ;
        RECT 4.300 467.300 315.700 468.460 ;
        RECT 2.330 465.660 317.990 467.300 ;
        RECT 4.300 464.500 315.700 465.660 ;
        RECT 2.330 462.860 317.990 464.500 ;
        RECT 4.300 461.700 315.700 462.860 ;
        RECT 2.330 460.060 317.990 461.700 ;
        RECT 4.300 458.900 315.700 460.060 ;
        RECT 2.330 457.260 317.990 458.900 ;
        RECT 4.300 456.100 315.700 457.260 ;
        RECT 2.330 454.460 317.990 456.100 ;
        RECT 4.300 453.300 315.700 454.460 ;
        RECT 2.330 451.660 317.990 453.300 ;
        RECT 4.300 450.500 315.700 451.660 ;
        RECT 2.330 448.860 317.990 450.500 ;
        RECT 4.300 447.700 315.700 448.860 ;
        RECT 2.330 446.060 317.990 447.700 ;
        RECT 4.300 444.900 315.700 446.060 ;
        RECT 2.330 443.260 317.990 444.900 ;
        RECT 4.300 442.100 315.700 443.260 ;
        RECT 2.330 440.460 317.990 442.100 ;
        RECT 4.300 439.300 315.700 440.460 ;
        RECT 2.330 437.660 317.990 439.300 ;
        RECT 4.300 436.500 315.700 437.660 ;
        RECT 2.330 434.860 317.990 436.500 ;
        RECT 4.300 433.700 315.700 434.860 ;
        RECT 2.330 432.060 317.990 433.700 ;
        RECT 4.300 430.900 315.700 432.060 ;
        RECT 2.330 429.260 317.990 430.900 ;
        RECT 4.300 428.100 315.700 429.260 ;
        RECT 2.330 426.460 317.990 428.100 ;
        RECT 4.300 425.300 315.700 426.460 ;
        RECT 2.330 423.660 317.990 425.300 ;
        RECT 4.300 422.500 315.700 423.660 ;
        RECT 2.330 420.860 317.990 422.500 ;
        RECT 4.300 419.700 315.700 420.860 ;
        RECT 2.330 418.060 317.990 419.700 ;
        RECT 4.300 416.900 315.700 418.060 ;
        RECT 2.330 415.260 317.990 416.900 ;
        RECT 4.300 414.100 315.700 415.260 ;
        RECT 2.330 412.460 317.990 414.100 ;
        RECT 4.300 411.300 315.700 412.460 ;
        RECT 2.330 409.660 317.990 411.300 ;
        RECT 4.300 408.500 315.700 409.660 ;
        RECT 2.330 406.860 317.990 408.500 ;
        RECT 4.300 405.700 315.700 406.860 ;
        RECT 2.330 404.060 317.990 405.700 ;
        RECT 4.300 402.900 315.700 404.060 ;
        RECT 2.330 401.260 317.990 402.900 ;
        RECT 4.300 400.100 315.700 401.260 ;
        RECT 2.330 398.460 317.990 400.100 ;
        RECT 4.300 397.300 315.700 398.460 ;
        RECT 2.330 395.660 317.990 397.300 ;
        RECT 4.300 394.500 315.700 395.660 ;
        RECT 2.330 392.860 317.990 394.500 ;
        RECT 4.300 391.700 315.700 392.860 ;
        RECT 2.330 390.060 317.990 391.700 ;
        RECT 4.300 388.900 315.700 390.060 ;
        RECT 2.330 387.260 317.990 388.900 ;
        RECT 4.300 386.100 315.700 387.260 ;
        RECT 2.330 384.460 317.990 386.100 ;
        RECT 4.300 383.300 315.700 384.460 ;
        RECT 2.330 381.660 317.990 383.300 ;
        RECT 4.300 380.500 315.700 381.660 ;
        RECT 2.330 378.860 317.990 380.500 ;
        RECT 4.300 377.700 315.700 378.860 ;
        RECT 2.330 376.060 317.990 377.700 ;
        RECT 4.300 374.900 315.700 376.060 ;
        RECT 2.330 373.260 317.990 374.900 ;
        RECT 4.300 372.100 315.700 373.260 ;
        RECT 2.330 370.460 317.990 372.100 ;
        RECT 4.300 369.300 315.700 370.460 ;
        RECT 2.330 367.660 317.990 369.300 ;
        RECT 4.300 366.500 315.700 367.660 ;
        RECT 2.330 364.860 317.990 366.500 ;
        RECT 4.300 363.700 315.700 364.860 ;
        RECT 2.330 362.060 317.990 363.700 ;
        RECT 4.300 360.900 315.700 362.060 ;
        RECT 2.330 359.260 317.990 360.900 ;
        RECT 4.300 358.100 315.700 359.260 ;
        RECT 2.330 356.460 317.990 358.100 ;
        RECT 4.300 355.300 315.700 356.460 ;
        RECT 2.330 353.660 317.990 355.300 ;
        RECT 4.300 352.500 315.700 353.660 ;
        RECT 2.330 350.860 317.990 352.500 ;
        RECT 4.300 349.700 315.700 350.860 ;
        RECT 2.330 348.060 317.990 349.700 ;
        RECT 4.300 346.900 315.700 348.060 ;
        RECT 2.330 345.260 317.990 346.900 ;
        RECT 4.300 344.100 315.700 345.260 ;
        RECT 2.330 342.460 317.990 344.100 ;
        RECT 4.300 341.300 315.700 342.460 ;
        RECT 2.330 339.660 317.990 341.300 ;
        RECT 4.300 338.500 315.700 339.660 ;
        RECT 2.330 336.860 317.990 338.500 ;
        RECT 4.300 335.700 315.700 336.860 ;
        RECT 2.330 334.060 317.990 335.700 ;
        RECT 4.300 332.900 315.700 334.060 ;
        RECT 2.330 331.260 317.990 332.900 ;
        RECT 4.300 330.100 315.700 331.260 ;
        RECT 2.330 328.460 317.990 330.100 ;
        RECT 4.300 327.300 315.700 328.460 ;
        RECT 2.330 325.660 317.990 327.300 ;
        RECT 4.300 324.500 315.700 325.660 ;
        RECT 2.330 322.860 317.990 324.500 ;
        RECT 4.300 321.700 315.700 322.860 ;
        RECT 2.330 320.060 317.990 321.700 ;
        RECT 4.300 318.900 315.700 320.060 ;
        RECT 2.330 317.260 317.990 318.900 ;
        RECT 4.300 316.100 315.700 317.260 ;
        RECT 2.330 314.460 317.990 316.100 ;
        RECT 4.300 313.300 315.700 314.460 ;
        RECT 2.330 311.660 317.990 313.300 ;
        RECT 4.300 310.500 315.700 311.660 ;
        RECT 2.330 308.860 317.990 310.500 ;
        RECT 4.300 307.700 315.700 308.860 ;
        RECT 2.330 306.060 317.990 307.700 ;
        RECT 4.300 304.900 315.700 306.060 ;
        RECT 2.330 303.260 317.990 304.900 ;
        RECT 4.300 302.100 315.700 303.260 ;
        RECT 2.330 300.460 317.990 302.100 ;
        RECT 4.300 299.300 315.700 300.460 ;
        RECT 2.330 297.660 317.990 299.300 ;
        RECT 4.300 296.500 315.700 297.660 ;
        RECT 2.330 294.860 317.990 296.500 ;
        RECT 4.300 293.700 315.700 294.860 ;
        RECT 2.330 292.060 317.990 293.700 ;
        RECT 4.300 290.900 315.700 292.060 ;
        RECT 2.330 289.260 317.990 290.900 ;
        RECT 4.300 288.100 315.700 289.260 ;
        RECT 2.330 286.460 317.990 288.100 ;
        RECT 4.300 285.300 315.700 286.460 ;
        RECT 2.330 283.660 317.990 285.300 ;
        RECT 4.300 282.500 315.700 283.660 ;
        RECT 2.330 280.860 317.990 282.500 ;
        RECT 4.300 279.700 315.700 280.860 ;
        RECT 2.330 278.060 317.990 279.700 ;
        RECT 4.300 276.900 315.700 278.060 ;
        RECT 2.330 275.260 317.990 276.900 ;
        RECT 4.300 274.100 315.700 275.260 ;
        RECT 2.330 272.460 317.990 274.100 ;
        RECT 4.300 271.300 315.700 272.460 ;
        RECT 2.330 269.660 317.990 271.300 ;
        RECT 4.300 268.500 315.700 269.660 ;
        RECT 2.330 266.860 317.990 268.500 ;
        RECT 4.300 265.700 315.700 266.860 ;
        RECT 2.330 264.060 317.990 265.700 ;
        RECT 4.300 262.900 315.700 264.060 ;
        RECT 2.330 261.260 317.990 262.900 ;
        RECT 4.300 260.100 315.700 261.260 ;
        RECT 2.330 258.460 317.990 260.100 ;
        RECT 4.300 257.300 315.700 258.460 ;
        RECT 2.330 255.660 317.990 257.300 ;
        RECT 4.300 254.500 315.700 255.660 ;
        RECT 2.330 252.860 317.990 254.500 ;
        RECT 4.300 251.700 315.700 252.860 ;
        RECT 2.330 250.060 317.990 251.700 ;
        RECT 4.300 248.900 315.700 250.060 ;
        RECT 2.330 247.260 317.990 248.900 ;
        RECT 4.300 246.100 315.700 247.260 ;
        RECT 2.330 244.460 317.990 246.100 ;
        RECT 4.300 243.300 315.700 244.460 ;
        RECT 2.330 241.660 317.990 243.300 ;
        RECT 4.300 240.500 315.700 241.660 ;
        RECT 2.330 238.860 317.990 240.500 ;
        RECT 4.300 237.700 315.700 238.860 ;
        RECT 2.330 236.060 317.990 237.700 ;
        RECT 4.300 234.900 315.700 236.060 ;
        RECT 2.330 233.260 317.990 234.900 ;
        RECT 4.300 232.100 315.700 233.260 ;
        RECT 2.330 230.460 317.990 232.100 ;
        RECT 4.300 229.300 315.700 230.460 ;
        RECT 2.330 227.660 317.990 229.300 ;
        RECT 4.300 226.500 315.700 227.660 ;
        RECT 2.330 224.860 317.990 226.500 ;
        RECT 4.300 223.700 315.700 224.860 ;
        RECT 2.330 222.060 317.990 223.700 ;
        RECT 4.300 220.900 315.700 222.060 ;
        RECT 2.330 219.260 317.990 220.900 ;
        RECT 4.300 218.100 315.700 219.260 ;
        RECT 2.330 216.460 317.990 218.100 ;
        RECT 4.300 215.300 315.700 216.460 ;
        RECT 2.330 213.660 317.990 215.300 ;
        RECT 4.300 212.500 315.700 213.660 ;
        RECT 2.330 210.860 317.990 212.500 ;
        RECT 4.300 209.700 315.700 210.860 ;
        RECT 2.330 208.060 317.990 209.700 ;
        RECT 4.300 206.900 315.700 208.060 ;
        RECT 2.330 205.260 317.990 206.900 ;
        RECT 4.300 204.100 315.700 205.260 ;
        RECT 2.330 202.460 317.990 204.100 ;
        RECT 4.300 201.300 315.700 202.460 ;
        RECT 2.330 199.660 317.990 201.300 ;
        RECT 4.300 198.500 315.700 199.660 ;
        RECT 2.330 196.860 317.990 198.500 ;
        RECT 4.300 195.700 315.700 196.860 ;
        RECT 2.330 194.060 317.990 195.700 ;
        RECT 4.300 192.900 315.700 194.060 ;
        RECT 2.330 191.260 317.990 192.900 ;
        RECT 4.300 190.100 315.700 191.260 ;
        RECT 2.330 188.460 317.990 190.100 ;
        RECT 4.300 187.300 315.700 188.460 ;
        RECT 2.330 185.660 317.990 187.300 ;
        RECT 4.300 184.500 315.700 185.660 ;
        RECT 2.330 15.540 317.990 184.500 ;
      LAYER Metal4 ;
        RECT 7.420 205.050 21.940 2679.510 ;
        RECT 24.140 205.050 98.740 2679.510 ;
        RECT 100.940 205.050 175.540 2679.510 ;
        RECT 177.740 205.050 252.340 2679.510 ;
        RECT 254.540 205.050 314.020 2679.510 ;
  END
END ita
END LIBRARY

