VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO ita27
  CLASS BLOCK ;
  FOREIGN ita27 ;
  ORIGIN 0.000 0.000 ;
  SIZE 210.000 BY 210.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 141.120 4.000 141.680 ;
    END
  END clk
  PIN segm[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 206.000 100.800 210.000 101.360 ;
    END
  END segm[0]
  PIN segm[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 206.000 80.640 210.000 81.200 ;
    END
  END segm[10]
  PIN segm[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 131.040 0.000 131.600 4.000 ;
    END
  END segm[11]
  PIN segm[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 206.000 104.160 210.000 104.720 ;
    END
  END segm[12]
  PIN segm[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 110.880 4.000 111.440 ;
    END
  END segm[13]
  PIN segm[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 87.360 4.000 87.920 ;
    END
  END segm[1]
  PIN segm[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 206.000 124.320 210.000 124.880 ;
    END
  END segm[2]
  PIN segm[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 90.720 0.000 91.280 4.000 ;
    END
  END segm[3]
  PIN segm[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 90.720 4.000 91.280 ;
    END
  END segm[4]
  PIN segm[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 124.320 206.000 124.880 210.000 ;
    END
  END segm[5]
  PIN segm[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 131.040 206.000 131.600 210.000 ;
    END
  END segm[6]
  PIN segm[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 127.680 206.000 128.240 210.000 ;
    END
  END segm[7]
  PIN segm[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 206.000 87.360 210.000 87.920 ;
    END
  END segm[8]
  PIN segm[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 107.520 0.000 108.080 4.000 ;
    END
  END segm[9]
  PIN sel[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 84.000 206.000 84.560 210.000 ;
    END
  END sel[0]
  PIN sel[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 104.160 4.000 104.720 ;
    END
  END sel[10]
  PIN sel[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 110.880 0.000 111.440 4.000 ;
    END
  END sel[11]
  PIN sel[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 100.800 206.000 101.360 210.000 ;
    END
  END sel[1]
  PIN sel[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 94.080 206.000 94.640 210.000 ;
    END
  END sel[2]
  PIN sel[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 114.240 206.000 114.800 210.000 ;
    END
  END sel[3]
  PIN sel[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 206.000 117.600 210.000 118.160 ;
    END
  END sel[4]
  PIN sel[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 127.680 4.000 128.240 ;
    END
  END sel[5]
  PIN sel[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 206.000 97.440 210.000 98.000 ;
    END
  END sel[6]
  PIN sel[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 117.600 4.000 118.160 ;
    END
  END sel[7]
  PIN sel[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 97.440 0.000 98.000 4.000 ;
    END
  END sel[8]
  PIN sel[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 206.000 127.680 210.000 128.240 ;
    END
  END sel[9]
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 192.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 192.380 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 192.380 ;
    END
  END vss
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 203.280 192.380 ;
      LAYER Metal2 ;
        RECT 9.660 205.700 83.700 206.000 ;
        RECT 84.860 205.700 93.780 206.000 ;
        RECT 94.940 205.700 100.500 206.000 ;
        RECT 101.660 205.700 113.940 206.000 ;
        RECT 115.100 205.700 124.020 206.000 ;
        RECT 125.180 205.700 127.380 206.000 ;
        RECT 128.540 205.700 130.740 206.000 ;
        RECT 131.900 205.700 201.460 206.000 ;
        RECT 9.660 4.300 201.460 205.700 ;
        RECT 9.660 4.000 90.420 4.300 ;
        RECT 91.580 4.000 97.140 4.300 ;
        RECT 98.300 4.000 107.220 4.300 ;
        RECT 108.380 4.000 110.580 4.300 ;
        RECT 111.740 4.000 130.740 4.300 ;
        RECT 131.900 4.000 201.460 4.300 ;
      LAYER Metal3 ;
        RECT 4.000 141.980 206.000 193.060 ;
        RECT 4.300 140.820 206.000 141.980 ;
        RECT 4.000 128.540 206.000 140.820 ;
        RECT 4.300 127.380 205.700 128.540 ;
        RECT 4.000 125.180 206.000 127.380 ;
        RECT 4.000 124.020 205.700 125.180 ;
        RECT 4.000 118.460 206.000 124.020 ;
        RECT 4.300 117.300 205.700 118.460 ;
        RECT 4.000 111.740 206.000 117.300 ;
        RECT 4.300 110.580 206.000 111.740 ;
        RECT 4.000 105.020 206.000 110.580 ;
        RECT 4.300 103.860 205.700 105.020 ;
        RECT 4.000 101.660 206.000 103.860 ;
        RECT 4.000 100.500 205.700 101.660 ;
        RECT 4.000 98.300 206.000 100.500 ;
        RECT 4.000 97.140 205.700 98.300 ;
        RECT 4.000 91.580 206.000 97.140 ;
        RECT 4.300 90.420 206.000 91.580 ;
        RECT 4.000 88.220 206.000 90.420 ;
        RECT 4.300 87.060 205.700 88.220 ;
        RECT 4.000 81.500 206.000 87.060 ;
        RECT 4.000 80.340 205.700 81.500 ;
        RECT 4.000 15.540 206.000 80.340 ;
      LAYER Metal4 ;
        RECT 91.420 107.050 91.700 110.230 ;
  END
END ita27
END LIBRARY

