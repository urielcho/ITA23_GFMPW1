magic
tech gf180mcuD
magscale 1 5
timestamp 1699642741
<< metal1 >>
rect 672 19221 20328 19238
rect 672 19195 2239 19221
rect 2265 19195 2291 19221
rect 2317 19195 2343 19221
rect 2369 19195 17599 19221
rect 17625 19195 17651 19221
rect 17677 19195 17703 19221
rect 17729 19195 20328 19221
rect 672 19178 20328 19195
rect 12783 19137 12809 19143
rect 12783 19105 12809 19111
rect 12441 18999 12447 19025
rect 12473 18999 12479 19025
rect 8527 18969 8553 18975
rect 8527 18937 8553 18943
rect 672 18829 20328 18846
rect 672 18803 9919 18829
rect 9945 18803 9971 18829
rect 9997 18803 10023 18829
rect 10049 18803 20328 18829
rect 672 18786 20328 18803
rect 13119 18745 13145 18751
rect 13119 18713 13145 18719
rect 12609 18607 12615 18633
rect 12641 18607 12647 18633
rect 672 18437 20328 18454
rect 672 18411 2239 18437
rect 2265 18411 2291 18437
rect 2317 18411 2343 18437
rect 2369 18411 17599 18437
rect 17625 18411 17651 18437
rect 17677 18411 17703 18437
rect 17729 18411 20328 18437
rect 672 18394 20328 18411
rect 13063 18353 13089 18359
rect 13063 18321 13089 18327
rect 12665 18215 12671 18241
rect 12697 18215 12703 18241
rect 672 18045 20328 18062
rect 672 18019 9919 18045
rect 9945 18019 9971 18045
rect 9997 18019 10023 18045
rect 10049 18019 20328 18045
rect 672 18002 20328 18019
rect 672 17653 20328 17670
rect 672 17627 2239 17653
rect 2265 17627 2291 17653
rect 2317 17627 2343 17653
rect 2369 17627 17599 17653
rect 17625 17627 17651 17653
rect 17677 17627 17703 17653
rect 17729 17627 20328 17653
rect 672 17610 20328 17627
rect 672 17261 20328 17278
rect 672 17235 9919 17261
rect 9945 17235 9971 17261
rect 9997 17235 10023 17261
rect 10049 17235 20328 17261
rect 672 17218 20328 17235
rect 672 16869 20328 16886
rect 672 16843 2239 16869
rect 2265 16843 2291 16869
rect 2317 16843 2343 16869
rect 2369 16843 17599 16869
rect 17625 16843 17651 16869
rect 17677 16843 17703 16869
rect 17729 16843 20328 16869
rect 672 16826 20328 16843
rect 672 16477 20328 16494
rect 672 16451 9919 16477
rect 9945 16451 9971 16477
rect 9997 16451 10023 16477
rect 10049 16451 20328 16477
rect 672 16434 20328 16451
rect 672 16085 20328 16102
rect 672 16059 2239 16085
rect 2265 16059 2291 16085
rect 2317 16059 2343 16085
rect 2369 16059 17599 16085
rect 17625 16059 17651 16085
rect 17677 16059 17703 16085
rect 17729 16059 20328 16085
rect 672 16042 20328 16059
rect 672 15693 20328 15710
rect 672 15667 9919 15693
rect 9945 15667 9971 15693
rect 9997 15667 10023 15693
rect 10049 15667 20328 15693
rect 672 15650 20328 15667
rect 672 15301 20328 15318
rect 672 15275 2239 15301
rect 2265 15275 2291 15301
rect 2317 15275 2343 15301
rect 2369 15275 17599 15301
rect 17625 15275 17651 15301
rect 17677 15275 17703 15301
rect 17729 15275 20328 15301
rect 672 15258 20328 15275
rect 672 14909 20328 14926
rect 672 14883 9919 14909
rect 9945 14883 9971 14909
rect 9997 14883 10023 14909
rect 10049 14883 20328 14909
rect 672 14866 20328 14883
rect 672 14517 20328 14534
rect 672 14491 2239 14517
rect 2265 14491 2291 14517
rect 2317 14491 2343 14517
rect 2369 14491 17599 14517
rect 17625 14491 17651 14517
rect 17677 14491 17703 14517
rect 17729 14491 20328 14517
rect 672 14474 20328 14491
rect 672 14125 20328 14142
rect 672 14099 9919 14125
rect 9945 14099 9971 14125
rect 9997 14099 10023 14125
rect 10049 14099 20328 14125
rect 672 14082 20328 14099
rect 672 13733 20328 13750
rect 672 13707 2239 13733
rect 2265 13707 2291 13733
rect 2317 13707 2343 13733
rect 2369 13707 17599 13733
rect 17625 13707 17651 13733
rect 17677 13707 17703 13733
rect 17729 13707 20328 13733
rect 672 13690 20328 13707
rect 672 13341 20328 13358
rect 672 13315 9919 13341
rect 9945 13315 9971 13341
rect 9997 13315 10023 13341
rect 10049 13315 20328 13341
rect 672 13298 20328 13315
rect 7575 13257 7601 13263
rect 12217 13231 12223 13257
rect 12249 13231 12255 13257
rect 7575 13225 7601 13231
rect 7519 13145 7545 13151
rect 12105 13119 12111 13145
rect 12137 13119 12143 13145
rect 7519 13113 7545 13119
rect 7575 13033 7601 13039
rect 7575 13001 7601 13007
rect 672 12949 20328 12966
rect 672 12923 2239 12949
rect 2265 12923 2291 12949
rect 2317 12923 2343 12949
rect 2369 12923 17599 12949
rect 17625 12923 17651 12949
rect 17677 12923 17703 12949
rect 17729 12923 20328 12949
rect 672 12906 20328 12923
rect 967 12809 993 12815
rect 12391 12809 12417 12815
rect 6729 12783 6735 12809
rect 6761 12783 6767 12809
rect 10089 12783 10095 12809
rect 10121 12783 10127 12809
rect 967 12777 993 12783
rect 12391 12777 12417 12783
rect 2137 12727 2143 12753
rect 2169 12727 2175 12753
rect 8185 12727 8191 12753
rect 8217 12727 8223 12753
rect 8689 12727 8695 12753
rect 8721 12727 8727 12753
rect 10985 12727 10991 12753
rect 11017 12727 11023 12753
rect 12777 12727 12783 12753
rect 12809 12727 12815 12753
rect 7793 12671 7799 12697
rect 7825 12671 7831 12697
rect 9025 12671 9031 12697
rect 9057 12671 9063 12697
rect 11321 12671 11327 12697
rect 11353 12671 11359 12697
rect 12665 12671 12671 12697
rect 12697 12671 12703 12697
rect 672 12557 20328 12574
rect 672 12531 9919 12557
rect 9945 12531 9971 12557
rect 9997 12531 10023 12557
rect 10049 12531 20328 12557
rect 672 12514 20328 12531
rect 8079 12473 8105 12479
rect 8079 12441 8105 12447
rect 8359 12473 8385 12479
rect 8359 12441 8385 12447
rect 11159 12473 11185 12479
rect 11159 12441 11185 12447
rect 7967 12417 7993 12423
rect 7967 12385 7993 12391
rect 11551 12417 11577 12423
rect 11551 12385 11577 12391
rect 7855 12361 7881 12367
rect 2137 12335 2143 12361
rect 2169 12335 2175 12361
rect 7681 12335 7687 12361
rect 7713 12335 7719 12361
rect 7855 12329 7881 12335
rect 8303 12361 8329 12367
rect 8303 12329 8329 12335
rect 8471 12361 8497 12367
rect 10431 12361 10457 12367
rect 11383 12361 11409 12367
rect 8689 12335 8695 12361
rect 8721 12335 8727 12361
rect 11041 12335 11047 12361
rect 11073 12335 11079 12361
rect 8471 12329 8497 12335
rect 10431 12329 10457 12335
rect 11383 12329 11409 12335
rect 11607 12361 11633 12367
rect 11607 12329 11633 12335
rect 11831 12361 11857 12367
rect 11831 12329 11857 12335
rect 11943 12361 11969 12367
rect 11943 12329 11969 12335
rect 12167 12361 12193 12367
rect 18825 12335 18831 12361
rect 18857 12335 18863 12361
rect 12167 12329 12193 12335
rect 7911 12305 7937 12311
rect 10319 12305 10345 12311
rect 6225 12279 6231 12305
rect 6257 12279 6263 12305
rect 7289 12279 7295 12305
rect 7321 12279 7327 12305
rect 9081 12279 9087 12305
rect 9113 12279 9119 12305
rect 10145 12279 10151 12305
rect 10177 12279 10183 12305
rect 7911 12273 7937 12279
rect 10319 12273 10345 12279
rect 11439 12305 11465 12311
rect 11439 12273 11465 12279
rect 11887 12305 11913 12311
rect 11887 12273 11913 12279
rect 967 12249 993 12255
rect 11215 12249 11241 12255
rect 10593 12223 10599 12249
rect 10625 12223 10631 12249
rect 967 12217 993 12223
rect 11215 12217 11241 12223
rect 20007 12249 20033 12255
rect 20007 12217 20033 12223
rect 672 12165 20328 12182
rect 672 12139 2239 12165
rect 2265 12139 2291 12165
rect 2317 12139 2343 12165
rect 2369 12139 17599 12165
rect 17625 12139 17651 12165
rect 17677 12139 17703 12165
rect 17729 12139 20328 12165
rect 672 12122 20328 12139
rect 13007 12081 13033 12087
rect 13007 12049 13033 12055
rect 7295 12025 7321 12031
rect 7295 11993 7321 11999
rect 9255 12025 9281 12031
rect 11713 11999 11719 12025
rect 11745 11999 11751 12025
rect 12777 11999 12783 12025
rect 12809 11999 12815 12025
rect 9255 11993 9281 11999
rect 7519 11969 7545 11975
rect 7519 11937 7545 11943
rect 7631 11969 7657 11975
rect 7631 11937 7657 11943
rect 7855 11969 7881 11975
rect 7855 11937 7881 11943
rect 7911 11969 7937 11975
rect 9311 11969 9337 11975
rect 9025 11943 9031 11969
rect 9057 11943 9063 11969
rect 7911 11937 7937 11943
rect 9311 11937 9337 11943
rect 10095 11969 10121 11975
rect 10095 11937 10121 11943
rect 10375 11969 10401 11975
rect 11377 11943 11383 11969
rect 11409 11943 11415 11969
rect 10375 11937 10401 11943
rect 7239 11913 7265 11919
rect 7239 11881 7265 11887
rect 7407 11913 7433 11919
rect 9199 11913 9225 11919
rect 13007 11913 13033 11919
rect 8689 11887 8695 11913
rect 8721 11887 8727 11913
rect 9753 11887 9759 11913
rect 9785 11887 9791 11913
rect 7407 11881 7433 11887
rect 9199 11881 9225 11887
rect 13007 11881 13033 11887
rect 13063 11913 13089 11919
rect 13063 11881 13089 11887
rect 7799 11857 7825 11863
rect 7799 11825 7825 11831
rect 8863 11857 8889 11863
rect 8863 11825 8889 11831
rect 9927 11857 9953 11863
rect 9927 11825 9953 11831
rect 672 11773 20328 11790
rect 672 11747 9919 11773
rect 9945 11747 9971 11773
rect 9997 11747 10023 11773
rect 10049 11747 20328 11773
rect 672 11730 20328 11747
rect 7183 11689 7209 11695
rect 7183 11657 7209 11663
rect 9367 11689 9393 11695
rect 9367 11657 9393 11663
rect 9703 11689 9729 11695
rect 9703 11657 9729 11663
rect 9927 11689 9953 11695
rect 10537 11663 10543 11689
rect 10569 11663 10575 11689
rect 9927 11657 9953 11663
rect 13455 11633 13481 11639
rect 7793 11607 7799 11633
rect 7825 11607 7831 11633
rect 9529 11607 9535 11633
rect 9561 11607 9567 11633
rect 10313 11607 10319 11633
rect 10345 11607 10351 11633
rect 10425 11607 10431 11633
rect 10457 11607 10463 11633
rect 13455 11601 13481 11607
rect 13791 11633 13817 11639
rect 13791 11601 13817 11607
rect 7295 11577 7321 11583
rect 9311 11577 9337 11583
rect 2137 11551 2143 11577
rect 2169 11551 2175 11577
rect 7457 11551 7463 11577
rect 7489 11551 7495 11577
rect 7681 11551 7687 11577
rect 7713 11551 7719 11577
rect 7295 11545 7321 11551
rect 9311 11545 9337 11551
rect 9983 11577 10009 11583
rect 9983 11545 10009 11551
rect 10711 11577 10737 11583
rect 10711 11545 10737 11551
rect 13343 11577 13369 11583
rect 13343 11545 13369 11551
rect 13511 11577 13537 11583
rect 13511 11545 13537 11551
rect 13679 11577 13705 11583
rect 13679 11545 13705 11551
rect 13847 11577 13873 11583
rect 18825 11551 18831 11577
rect 18857 11551 18863 11577
rect 13847 11545 13873 11551
rect 7239 11521 7265 11527
rect 7239 11489 7265 11495
rect 967 11465 993 11471
rect 967 11433 993 11439
rect 9927 11465 9953 11471
rect 9927 11433 9953 11439
rect 20007 11465 20033 11471
rect 20007 11433 20033 11439
rect 672 11381 20328 11398
rect 672 11355 2239 11381
rect 2265 11355 2291 11381
rect 2317 11355 2343 11381
rect 2369 11355 17599 11381
rect 17625 11355 17651 11381
rect 17677 11355 17703 11381
rect 17729 11355 20328 11381
rect 672 11338 20328 11355
rect 10985 11271 10991 11297
rect 11017 11271 11023 11297
rect 11657 11271 11663 11297
rect 11689 11271 11695 11297
rect 967 11241 993 11247
rect 20007 11241 20033 11247
rect 9417 11215 9423 11241
rect 9449 11215 9455 11241
rect 10817 11215 10823 11241
rect 10849 11215 10855 11241
rect 13225 11215 13231 11241
rect 13257 11215 13263 11241
rect 14289 11215 14295 11241
rect 14321 11215 14327 11241
rect 967 11209 993 11215
rect 20007 11209 20033 11215
rect 7015 11185 7041 11191
rect 2137 11159 2143 11185
rect 2169 11159 2175 11185
rect 7015 11153 7041 11159
rect 7127 11185 7153 11191
rect 7127 11153 7153 11159
rect 7351 11185 7377 11191
rect 7351 11153 7377 11159
rect 7407 11185 7433 11191
rect 7407 11153 7433 11159
rect 7631 11185 7657 11191
rect 7631 11153 7657 11159
rect 9647 11185 9673 11191
rect 10761 11159 10767 11185
rect 10793 11159 10799 11185
rect 11657 11159 11663 11185
rect 11689 11159 11695 11185
rect 12833 11159 12839 11185
rect 12865 11159 12871 11185
rect 18825 11159 18831 11185
rect 18857 11159 18863 11185
rect 9647 11153 9673 11159
rect 6847 11129 6873 11135
rect 11943 11129 11969 11135
rect 11825 11103 11831 11129
rect 11857 11103 11863 11129
rect 6847 11097 6873 11103
rect 11943 11097 11969 11103
rect 6903 11073 6929 11079
rect 6903 11041 6929 11047
rect 7519 11073 7545 11079
rect 9983 11073 10009 11079
rect 9809 11047 9815 11073
rect 9841 11047 9847 11073
rect 7519 11041 7545 11047
rect 9983 11041 10009 11047
rect 11551 11073 11577 11079
rect 11551 11041 11577 11047
rect 672 10989 20328 11006
rect 672 10963 9919 10989
rect 9945 10963 9971 10989
rect 9997 10963 10023 10989
rect 10049 10963 20328 10989
rect 672 10946 20328 10963
rect 7519 10905 7545 10911
rect 7519 10873 7545 10879
rect 10767 10905 10793 10911
rect 10767 10873 10793 10879
rect 7463 10849 7489 10855
rect 6729 10823 6735 10849
rect 6761 10823 6767 10849
rect 7463 10817 7489 10823
rect 8191 10849 8217 10855
rect 14905 10823 14911 10849
rect 14937 10823 14943 10849
rect 8191 10817 8217 10823
rect 7575 10793 7601 10799
rect 8135 10793 8161 10799
rect 9759 10793 9785 10799
rect 10599 10793 10625 10799
rect 7065 10767 7071 10793
rect 7097 10767 7103 10793
rect 7737 10767 7743 10793
rect 7769 10767 7775 10793
rect 8969 10767 8975 10793
rect 9001 10767 9007 10793
rect 10145 10767 10151 10793
rect 10177 10767 10183 10793
rect 10369 10767 10375 10793
rect 10401 10767 10407 10793
rect 10929 10767 10935 10793
rect 10961 10767 10967 10793
rect 13169 10767 13175 10793
rect 13201 10767 13207 10793
rect 14793 10767 14799 10793
rect 14825 10767 14831 10793
rect 18825 10767 18831 10793
rect 18857 10767 18863 10793
rect 7575 10761 7601 10767
rect 8135 10761 8161 10767
rect 9759 10761 9785 10767
rect 10599 10761 10625 10767
rect 9199 10737 9225 10743
rect 5665 10711 5671 10737
rect 5697 10711 5703 10737
rect 8745 10711 8751 10737
rect 8777 10711 8783 10737
rect 9199 10705 9225 10711
rect 9647 10737 9673 10743
rect 20007 10737 20033 10743
rect 11265 10711 11271 10737
rect 11297 10711 11303 10737
rect 12329 10711 12335 10737
rect 12361 10711 12367 10737
rect 13505 10711 13511 10737
rect 13537 10711 13543 10737
rect 14569 10711 14575 10737
rect 14601 10711 14607 10737
rect 9647 10705 9673 10711
rect 20007 10705 20033 10711
rect 9927 10681 9953 10687
rect 9927 10649 9953 10655
rect 672 10597 20328 10614
rect 672 10571 2239 10597
rect 2265 10571 2291 10597
rect 2317 10571 2343 10597
rect 2369 10571 17599 10597
rect 17625 10571 17651 10597
rect 17677 10571 17703 10597
rect 17729 10571 20328 10597
rect 672 10554 20328 10571
rect 20007 10457 20033 10463
rect 20007 10425 20033 10431
rect 10033 10375 10039 10401
rect 10065 10375 10071 10401
rect 11321 10375 11327 10401
rect 11353 10375 11359 10401
rect 11657 10375 11663 10401
rect 11689 10375 11695 10401
rect 18825 10375 18831 10401
rect 18857 10375 18863 10401
rect 10655 10345 10681 10351
rect 8129 10319 8135 10345
rect 8161 10319 8167 10345
rect 11041 10319 11047 10345
rect 11073 10319 11079 10345
rect 13169 10319 13175 10345
rect 13201 10319 13207 10345
rect 10655 10313 10681 10319
rect 10711 10289 10737 10295
rect 11321 10263 11327 10289
rect 11353 10263 11359 10289
rect 10711 10257 10737 10263
rect 672 10205 20328 10222
rect 672 10179 9919 10205
rect 9945 10179 9971 10205
rect 9997 10179 10023 10205
rect 10049 10179 20328 10205
rect 672 10162 20328 10179
rect 8919 10065 8945 10071
rect 7793 10039 7799 10065
rect 7825 10039 7831 10065
rect 8919 10033 8945 10039
rect 8975 10065 9001 10071
rect 8975 10033 9001 10039
rect 9031 10065 9057 10071
rect 13287 10065 13313 10071
rect 9529 10039 9535 10065
rect 9561 10039 9567 10065
rect 11657 10039 11663 10065
rect 11689 10039 11695 10065
rect 12777 10039 12783 10065
rect 12809 10039 12815 10065
rect 9031 10033 9057 10039
rect 13287 10033 13313 10039
rect 13791 10065 13817 10071
rect 13791 10033 13817 10039
rect 13847 10065 13873 10071
rect 13847 10033 13873 10039
rect 13231 10009 13257 10015
rect 8129 9983 8135 10009
rect 8161 9983 8167 10009
rect 9417 9983 9423 10009
rect 9449 9983 9455 10009
rect 9697 9983 9703 10009
rect 9729 9983 9735 10009
rect 12665 9983 12671 10009
rect 12697 9983 12703 10009
rect 13231 9977 13257 9983
rect 13343 10009 13369 10015
rect 13343 9977 13369 9983
rect 13567 10009 13593 10015
rect 18937 9983 18943 10009
rect 18969 9983 18975 10009
rect 13567 9977 13593 9983
rect 20007 9953 20033 9959
rect 6729 9927 6735 9953
rect 6761 9927 6767 9953
rect 20007 9921 20033 9927
rect 9479 9897 9505 9903
rect 9479 9865 9505 9871
rect 13847 9897 13873 9903
rect 13847 9865 13873 9871
rect 672 9813 20328 9830
rect 672 9787 2239 9813
rect 2265 9787 2291 9813
rect 2317 9787 2343 9813
rect 2369 9787 17599 9813
rect 17625 9787 17651 9813
rect 17677 9787 17703 9813
rect 17729 9787 20328 9813
rect 672 9770 20328 9787
rect 10263 9729 10289 9735
rect 20007 9729 20033 9735
rect 12049 9703 12055 9729
rect 12081 9703 12087 9729
rect 10263 9697 10289 9703
rect 20007 9697 20033 9703
rect 9311 9673 9337 9679
rect 12279 9673 12305 9679
rect 8409 9647 8415 9673
rect 8441 9647 8447 9673
rect 9641 9647 9647 9673
rect 9673 9647 9679 9673
rect 9311 9641 9337 9647
rect 12279 9641 12305 9647
rect 12503 9673 12529 9679
rect 12503 9641 12529 9647
rect 9423 9617 9449 9623
rect 7009 9591 7015 9617
rect 7041 9591 7047 9617
rect 9423 9585 9449 9591
rect 9983 9617 10009 9623
rect 10991 9617 11017 9623
rect 10089 9591 10095 9617
rect 10121 9591 10127 9617
rect 9983 9585 10009 9591
rect 10991 9585 11017 9591
rect 11103 9617 11129 9623
rect 11103 9585 11129 9591
rect 11327 9617 11353 9623
rect 11327 9585 11353 9591
rect 11439 9617 11465 9623
rect 13679 9617 13705 9623
rect 11937 9591 11943 9617
rect 11969 9591 11975 9617
rect 11439 9585 11465 9591
rect 13679 9585 13705 9591
rect 13847 9617 13873 9623
rect 13847 9585 13873 9591
rect 14575 9617 14601 9623
rect 18825 9591 18831 9617
rect 18857 9591 18863 9617
rect 14575 9585 14601 9591
rect 12335 9561 12361 9567
rect 7345 9535 7351 9561
rect 7377 9535 7383 9561
rect 10817 9535 10823 9561
rect 10849 9535 10855 9561
rect 12217 9535 12223 9561
rect 12249 9535 12255 9561
rect 12335 9529 12361 9535
rect 12895 9561 12921 9567
rect 12895 9529 12921 9535
rect 13511 9561 13537 9567
rect 13511 9529 13537 9535
rect 9927 9505 9953 9511
rect 9927 9473 9953 9479
rect 10039 9505 10065 9511
rect 10039 9473 10065 9479
rect 11271 9505 11297 9511
rect 11271 9473 11297 9479
rect 12559 9505 12585 9511
rect 12559 9473 12585 9479
rect 12615 9505 12641 9511
rect 13735 9505 13761 9511
rect 13057 9479 13063 9505
rect 13089 9479 13095 9505
rect 14737 9479 14743 9505
rect 14769 9479 14775 9505
rect 12615 9473 12641 9479
rect 13735 9473 13761 9479
rect 672 9421 20328 9438
rect 672 9395 9919 9421
rect 9945 9395 9971 9421
rect 9997 9395 10023 9421
rect 10049 9395 20328 9421
rect 672 9378 20328 9395
rect 7575 9337 7601 9343
rect 7575 9305 7601 9311
rect 9199 9337 9225 9343
rect 12895 9337 12921 9343
rect 9697 9311 9703 9337
rect 9729 9311 9735 9337
rect 11657 9311 11663 9337
rect 11689 9311 11695 9337
rect 9199 9305 9225 9311
rect 12895 9305 12921 9311
rect 14855 9337 14881 9343
rect 14855 9305 14881 9311
rect 7687 9281 7713 9287
rect 7687 9249 7713 9255
rect 7911 9281 7937 9287
rect 7911 9249 7937 9255
rect 7967 9281 7993 9287
rect 11215 9281 11241 9287
rect 9025 9255 9031 9281
rect 9057 9255 9063 9281
rect 9921 9255 9927 9281
rect 9953 9255 9959 9281
rect 13057 9255 13063 9281
rect 13089 9255 13095 9281
rect 15353 9255 15359 9281
rect 15385 9255 15391 9281
rect 7967 9249 7993 9255
rect 11215 9249 11241 9255
rect 7351 9225 7377 9231
rect 2137 9199 2143 9225
rect 2169 9199 2175 9225
rect 7177 9199 7183 9225
rect 7209 9199 7215 9225
rect 7351 9193 7377 9199
rect 7799 9225 7825 9231
rect 7799 9193 7825 9199
rect 9535 9225 9561 9231
rect 10935 9225 10961 9231
rect 15023 9225 15049 9231
rect 9865 9199 9871 9225
rect 9897 9199 9903 9225
rect 13225 9199 13231 9225
rect 13257 9199 13263 9225
rect 9535 9193 9561 9199
rect 10935 9193 10961 9199
rect 15023 9193 15049 9199
rect 15191 9225 15217 9231
rect 18825 9199 18831 9225
rect 18857 9199 18863 9225
rect 15191 9193 15217 9199
rect 7631 9169 7657 9175
rect 20007 9169 20033 9175
rect 5777 9143 5783 9169
rect 5809 9143 5815 9169
rect 6841 9143 6847 9169
rect 6873 9143 6879 9169
rect 13617 9143 13623 9169
rect 13649 9143 13655 9169
rect 14681 9143 14687 9169
rect 14713 9143 14719 9169
rect 7631 9137 7657 9143
rect 20007 9137 20033 9143
rect 967 9113 993 9119
rect 967 9081 993 9087
rect 672 9029 20328 9046
rect 672 9003 2239 9029
rect 2265 9003 2291 9029
rect 2317 9003 2343 9029
rect 2369 9003 17599 9029
rect 17625 9003 17651 9029
rect 17677 9003 17703 9029
rect 17729 9003 20328 9029
rect 672 8986 20328 9003
rect 8863 8945 8889 8951
rect 8863 8913 8889 8919
rect 14071 8945 14097 8951
rect 14071 8913 14097 8919
rect 967 8889 993 8895
rect 13287 8889 13313 8895
rect 9865 8863 9871 8889
rect 9897 8863 9903 8889
rect 12217 8863 12223 8889
rect 12249 8863 12255 8889
rect 967 8857 993 8863
rect 13287 8857 13313 8863
rect 14127 8889 14153 8895
rect 19945 8863 19951 8889
rect 19977 8863 19983 8889
rect 14127 8857 14153 8863
rect 6847 8833 6873 8839
rect 2137 8807 2143 8833
rect 2169 8807 2175 8833
rect 6847 8801 6873 8807
rect 6959 8833 6985 8839
rect 6959 8801 6985 8807
rect 7351 8833 7377 8839
rect 9647 8833 9673 8839
rect 9249 8807 9255 8833
rect 9281 8807 9287 8833
rect 7351 8801 7377 8807
rect 9647 8801 9673 8807
rect 10095 8833 10121 8839
rect 10095 8801 10121 8807
rect 10431 8833 10457 8839
rect 14575 8833 14601 8839
rect 10705 8807 10711 8833
rect 10737 8807 10743 8833
rect 11825 8807 11831 8833
rect 11857 8807 11863 8833
rect 18825 8807 18831 8833
rect 18857 8807 18863 8833
rect 10431 8801 10457 8807
rect 14575 8801 14601 8807
rect 7463 8777 7489 8783
rect 7463 8745 7489 8751
rect 7519 8777 7545 8783
rect 7519 8745 7545 8751
rect 8919 8777 8945 8783
rect 8919 8745 8945 8751
rect 9367 8777 9393 8783
rect 9367 8745 9393 8751
rect 10207 8777 10233 8783
rect 10207 8745 10233 8751
rect 6903 8721 6929 8727
rect 6903 8689 6929 8695
rect 7071 8721 7097 8727
rect 7071 8689 7097 8695
rect 8863 8721 8889 8727
rect 8863 8689 8889 8695
rect 9479 8721 9505 8727
rect 9479 8689 9505 8695
rect 9535 8721 9561 8727
rect 9535 8689 9561 8695
rect 10151 8721 10177 8727
rect 10817 8695 10823 8721
rect 10849 8695 10855 8721
rect 14737 8695 14743 8721
rect 14769 8695 14775 8721
rect 10151 8689 10177 8695
rect 672 8637 20328 8654
rect 672 8611 9919 8637
rect 9945 8611 9971 8637
rect 9997 8611 10023 8637
rect 10049 8611 20328 8637
rect 672 8594 20328 8611
rect 7575 8553 7601 8559
rect 7575 8521 7601 8527
rect 7687 8553 7713 8559
rect 7687 8521 7713 8527
rect 9535 8553 9561 8559
rect 9535 8521 9561 8527
rect 11047 8553 11073 8559
rect 11047 8521 11073 8527
rect 7743 8497 7769 8503
rect 7065 8471 7071 8497
rect 7097 8471 7103 8497
rect 7743 8465 7769 8471
rect 8303 8497 8329 8503
rect 8303 8465 8329 8471
rect 8359 8497 8385 8503
rect 8359 8465 8385 8471
rect 9031 8497 9057 8503
rect 9031 8465 9057 8471
rect 10935 8497 10961 8503
rect 10935 8465 10961 8471
rect 11383 8497 11409 8503
rect 19665 8471 19671 8497
rect 19697 8471 19703 8497
rect 11383 8465 11409 8471
rect 8471 8441 8497 8447
rect 7457 8415 7463 8441
rect 7489 8415 7495 8441
rect 8471 8409 8497 8415
rect 8919 8441 8945 8447
rect 8919 8409 8945 8415
rect 9199 8441 9225 8447
rect 9199 8409 9225 8415
rect 9591 8441 9617 8447
rect 9591 8409 9617 8415
rect 9703 8441 9729 8447
rect 9703 8409 9729 8415
rect 9927 8441 9953 8447
rect 9927 8409 9953 8415
rect 9983 8441 10009 8447
rect 9983 8409 10009 8415
rect 11103 8441 11129 8447
rect 11103 8409 11129 8415
rect 11159 8441 11185 8447
rect 11545 8415 11551 8441
rect 11577 8415 11583 8441
rect 18825 8415 18831 8441
rect 18857 8415 18863 8441
rect 11159 8409 11185 8415
rect 9311 8385 9337 8391
rect 6001 8359 6007 8385
rect 6033 8359 6039 8385
rect 9311 8353 9337 8359
rect 9815 8385 9841 8391
rect 9815 8353 9841 8359
rect 11439 8385 11465 8391
rect 11439 8353 11465 8359
rect 8975 8329 9001 8335
rect 8975 8297 9001 8303
rect 672 8245 20328 8262
rect 672 8219 2239 8245
rect 2265 8219 2291 8245
rect 2317 8219 2343 8245
rect 2369 8219 17599 8245
rect 17625 8219 17651 8245
rect 17677 8219 17703 8245
rect 17729 8219 20328 8245
rect 672 8202 20328 8219
rect 9927 8105 9953 8111
rect 7233 8079 7239 8105
rect 7265 8079 7271 8105
rect 8297 8079 8303 8105
rect 8329 8079 8335 8105
rect 8857 8079 8863 8105
rect 8889 8079 8895 8105
rect 11153 8079 11159 8105
rect 11185 8079 11191 8105
rect 12217 8079 12223 8105
rect 12249 8079 12255 8105
rect 19889 8079 19895 8105
rect 19921 8079 19927 8105
rect 9927 8073 9953 8079
rect 6897 8023 6903 8049
rect 6929 8023 6935 8049
rect 8521 8023 8527 8049
rect 8553 8023 8559 8049
rect 10817 8023 10823 8049
rect 10849 8023 10855 8049
rect 18825 8023 18831 8049
rect 18857 8023 18863 8049
rect 672 7853 20328 7870
rect 672 7827 9919 7853
rect 9945 7827 9971 7853
rect 9997 7827 10023 7853
rect 10049 7827 20328 7853
rect 672 7810 20328 7827
rect 9809 7687 9815 7713
rect 9841 7687 9847 7713
rect 11881 7687 11887 7713
rect 11913 7687 11919 7713
rect 9417 7631 9423 7657
rect 9449 7631 9455 7657
rect 11769 7631 11775 7657
rect 11801 7631 11807 7657
rect 18825 7631 18831 7657
rect 18857 7631 18863 7657
rect 20007 7601 20033 7607
rect 10873 7575 10879 7601
rect 10905 7575 10911 7601
rect 20007 7569 20033 7575
rect 672 7461 20328 7478
rect 672 7435 2239 7461
rect 2265 7435 2291 7461
rect 2317 7435 2343 7461
rect 2369 7435 17599 7461
rect 17625 7435 17651 7461
rect 17677 7435 17703 7461
rect 17729 7435 20328 7461
rect 672 7418 20328 7435
rect 672 7069 20328 7086
rect 672 7043 9919 7069
rect 9945 7043 9971 7069
rect 9997 7043 10023 7069
rect 10049 7043 20328 7069
rect 672 7026 20328 7043
rect 672 6677 20328 6694
rect 672 6651 2239 6677
rect 2265 6651 2291 6677
rect 2317 6651 2343 6677
rect 2369 6651 17599 6677
rect 17625 6651 17651 6677
rect 17677 6651 17703 6677
rect 17729 6651 20328 6677
rect 672 6634 20328 6651
rect 672 6285 20328 6302
rect 672 6259 9919 6285
rect 9945 6259 9971 6285
rect 9997 6259 10023 6285
rect 10049 6259 20328 6285
rect 672 6242 20328 6259
rect 672 5893 20328 5910
rect 672 5867 2239 5893
rect 2265 5867 2291 5893
rect 2317 5867 2343 5893
rect 2369 5867 17599 5893
rect 17625 5867 17651 5893
rect 17677 5867 17703 5893
rect 17729 5867 20328 5893
rect 672 5850 20328 5867
rect 672 5501 20328 5518
rect 672 5475 9919 5501
rect 9945 5475 9971 5501
rect 9997 5475 10023 5501
rect 10049 5475 20328 5501
rect 672 5458 20328 5475
rect 672 5109 20328 5126
rect 672 5083 2239 5109
rect 2265 5083 2291 5109
rect 2317 5083 2343 5109
rect 2369 5083 17599 5109
rect 17625 5083 17651 5109
rect 17677 5083 17703 5109
rect 17729 5083 20328 5109
rect 672 5066 20328 5083
rect 672 4717 20328 4734
rect 672 4691 9919 4717
rect 9945 4691 9971 4717
rect 9997 4691 10023 4717
rect 10049 4691 20328 4717
rect 672 4674 20328 4691
rect 672 4325 20328 4342
rect 672 4299 2239 4325
rect 2265 4299 2291 4325
rect 2317 4299 2343 4325
rect 2369 4299 17599 4325
rect 17625 4299 17651 4325
rect 17677 4299 17703 4325
rect 17729 4299 20328 4325
rect 672 4282 20328 4299
rect 672 3933 20328 3950
rect 672 3907 9919 3933
rect 9945 3907 9971 3933
rect 9997 3907 10023 3933
rect 10049 3907 20328 3933
rect 672 3890 20328 3907
rect 672 3541 20328 3558
rect 672 3515 2239 3541
rect 2265 3515 2291 3541
rect 2317 3515 2343 3541
rect 2369 3515 17599 3541
rect 17625 3515 17651 3541
rect 17677 3515 17703 3541
rect 17729 3515 20328 3541
rect 672 3498 20328 3515
rect 672 3149 20328 3166
rect 672 3123 9919 3149
rect 9945 3123 9971 3149
rect 9997 3123 10023 3149
rect 10049 3123 20328 3149
rect 672 3106 20328 3123
rect 672 2757 20328 2774
rect 672 2731 2239 2757
rect 2265 2731 2291 2757
rect 2317 2731 2343 2757
rect 2369 2731 17599 2757
rect 17625 2731 17651 2757
rect 17677 2731 17703 2757
rect 17729 2731 20328 2757
rect 672 2714 20328 2731
rect 12391 2617 12417 2623
rect 12391 2585 12417 2591
rect 11881 2535 11887 2561
rect 11913 2535 11919 2561
rect 672 2365 20328 2382
rect 672 2339 9919 2365
rect 9945 2339 9971 2365
rect 9997 2339 10023 2365
rect 10049 2339 20328 2365
rect 672 2322 20328 2339
rect 672 1973 20328 1990
rect 672 1947 2239 1973
rect 2265 1947 2291 1973
rect 2317 1947 2343 1973
rect 2369 1947 17599 1973
rect 17625 1947 17651 1973
rect 17677 1947 17703 1973
rect 17729 1947 20328 1973
rect 672 1930 20328 1947
rect 9311 1833 9337 1839
rect 9311 1801 9337 1807
rect 11047 1833 11073 1839
rect 11047 1801 11073 1807
rect 12783 1833 12809 1839
rect 12783 1801 12809 1807
rect 8801 1751 8807 1777
rect 8833 1751 8839 1777
rect 10537 1751 10543 1777
rect 10569 1751 10575 1777
rect 12273 1751 12279 1777
rect 12305 1751 12311 1777
rect 672 1581 20328 1598
rect 672 1555 9919 1581
rect 9945 1555 9971 1581
rect 9997 1555 10023 1581
rect 10049 1555 20328 1581
rect 672 1538 20328 1555
<< via1 >>
rect 2239 19195 2265 19221
rect 2291 19195 2317 19221
rect 2343 19195 2369 19221
rect 17599 19195 17625 19221
rect 17651 19195 17677 19221
rect 17703 19195 17729 19221
rect 12783 19111 12809 19137
rect 12447 18999 12473 19025
rect 8527 18943 8553 18969
rect 9919 18803 9945 18829
rect 9971 18803 9997 18829
rect 10023 18803 10049 18829
rect 13119 18719 13145 18745
rect 12615 18607 12641 18633
rect 2239 18411 2265 18437
rect 2291 18411 2317 18437
rect 2343 18411 2369 18437
rect 17599 18411 17625 18437
rect 17651 18411 17677 18437
rect 17703 18411 17729 18437
rect 13063 18327 13089 18353
rect 12671 18215 12697 18241
rect 9919 18019 9945 18045
rect 9971 18019 9997 18045
rect 10023 18019 10049 18045
rect 2239 17627 2265 17653
rect 2291 17627 2317 17653
rect 2343 17627 2369 17653
rect 17599 17627 17625 17653
rect 17651 17627 17677 17653
rect 17703 17627 17729 17653
rect 9919 17235 9945 17261
rect 9971 17235 9997 17261
rect 10023 17235 10049 17261
rect 2239 16843 2265 16869
rect 2291 16843 2317 16869
rect 2343 16843 2369 16869
rect 17599 16843 17625 16869
rect 17651 16843 17677 16869
rect 17703 16843 17729 16869
rect 9919 16451 9945 16477
rect 9971 16451 9997 16477
rect 10023 16451 10049 16477
rect 2239 16059 2265 16085
rect 2291 16059 2317 16085
rect 2343 16059 2369 16085
rect 17599 16059 17625 16085
rect 17651 16059 17677 16085
rect 17703 16059 17729 16085
rect 9919 15667 9945 15693
rect 9971 15667 9997 15693
rect 10023 15667 10049 15693
rect 2239 15275 2265 15301
rect 2291 15275 2317 15301
rect 2343 15275 2369 15301
rect 17599 15275 17625 15301
rect 17651 15275 17677 15301
rect 17703 15275 17729 15301
rect 9919 14883 9945 14909
rect 9971 14883 9997 14909
rect 10023 14883 10049 14909
rect 2239 14491 2265 14517
rect 2291 14491 2317 14517
rect 2343 14491 2369 14517
rect 17599 14491 17625 14517
rect 17651 14491 17677 14517
rect 17703 14491 17729 14517
rect 9919 14099 9945 14125
rect 9971 14099 9997 14125
rect 10023 14099 10049 14125
rect 2239 13707 2265 13733
rect 2291 13707 2317 13733
rect 2343 13707 2369 13733
rect 17599 13707 17625 13733
rect 17651 13707 17677 13733
rect 17703 13707 17729 13733
rect 9919 13315 9945 13341
rect 9971 13315 9997 13341
rect 10023 13315 10049 13341
rect 7575 13231 7601 13257
rect 12223 13231 12249 13257
rect 7519 13119 7545 13145
rect 12111 13119 12137 13145
rect 7575 13007 7601 13033
rect 2239 12923 2265 12949
rect 2291 12923 2317 12949
rect 2343 12923 2369 12949
rect 17599 12923 17625 12949
rect 17651 12923 17677 12949
rect 17703 12923 17729 12949
rect 967 12783 993 12809
rect 6735 12783 6761 12809
rect 10095 12783 10121 12809
rect 12391 12783 12417 12809
rect 2143 12727 2169 12753
rect 8191 12727 8217 12753
rect 8695 12727 8721 12753
rect 10991 12727 11017 12753
rect 12783 12727 12809 12753
rect 7799 12671 7825 12697
rect 9031 12671 9057 12697
rect 11327 12671 11353 12697
rect 12671 12671 12697 12697
rect 9919 12531 9945 12557
rect 9971 12531 9997 12557
rect 10023 12531 10049 12557
rect 8079 12447 8105 12473
rect 8359 12447 8385 12473
rect 11159 12447 11185 12473
rect 7967 12391 7993 12417
rect 11551 12391 11577 12417
rect 2143 12335 2169 12361
rect 7687 12335 7713 12361
rect 7855 12335 7881 12361
rect 8303 12335 8329 12361
rect 8471 12335 8497 12361
rect 8695 12335 8721 12361
rect 10431 12335 10457 12361
rect 11047 12335 11073 12361
rect 11383 12335 11409 12361
rect 11607 12335 11633 12361
rect 11831 12335 11857 12361
rect 11943 12335 11969 12361
rect 12167 12335 12193 12361
rect 18831 12335 18857 12361
rect 6231 12279 6257 12305
rect 7295 12279 7321 12305
rect 7911 12279 7937 12305
rect 9087 12279 9113 12305
rect 10151 12279 10177 12305
rect 10319 12279 10345 12305
rect 11439 12279 11465 12305
rect 11887 12279 11913 12305
rect 967 12223 993 12249
rect 10599 12223 10625 12249
rect 11215 12223 11241 12249
rect 20007 12223 20033 12249
rect 2239 12139 2265 12165
rect 2291 12139 2317 12165
rect 2343 12139 2369 12165
rect 17599 12139 17625 12165
rect 17651 12139 17677 12165
rect 17703 12139 17729 12165
rect 13007 12055 13033 12081
rect 7295 11999 7321 12025
rect 9255 11999 9281 12025
rect 11719 11999 11745 12025
rect 12783 11999 12809 12025
rect 7519 11943 7545 11969
rect 7631 11943 7657 11969
rect 7855 11943 7881 11969
rect 7911 11943 7937 11969
rect 9031 11943 9057 11969
rect 9311 11943 9337 11969
rect 10095 11943 10121 11969
rect 10375 11943 10401 11969
rect 11383 11943 11409 11969
rect 7239 11887 7265 11913
rect 7407 11887 7433 11913
rect 8695 11887 8721 11913
rect 9199 11887 9225 11913
rect 9759 11887 9785 11913
rect 13007 11887 13033 11913
rect 13063 11887 13089 11913
rect 7799 11831 7825 11857
rect 8863 11831 8889 11857
rect 9927 11831 9953 11857
rect 9919 11747 9945 11773
rect 9971 11747 9997 11773
rect 10023 11747 10049 11773
rect 7183 11663 7209 11689
rect 9367 11663 9393 11689
rect 9703 11663 9729 11689
rect 9927 11663 9953 11689
rect 10543 11663 10569 11689
rect 7799 11607 7825 11633
rect 9535 11607 9561 11633
rect 10319 11607 10345 11633
rect 10431 11607 10457 11633
rect 13455 11607 13481 11633
rect 13791 11607 13817 11633
rect 2143 11551 2169 11577
rect 7295 11551 7321 11577
rect 7463 11551 7489 11577
rect 7687 11551 7713 11577
rect 9311 11551 9337 11577
rect 9983 11551 10009 11577
rect 10711 11551 10737 11577
rect 13343 11551 13369 11577
rect 13511 11551 13537 11577
rect 13679 11551 13705 11577
rect 13847 11551 13873 11577
rect 18831 11551 18857 11577
rect 7239 11495 7265 11521
rect 967 11439 993 11465
rect 9927 11439 9953 11465
rect 20007 11439 20033 11465
rect 2239 11355 2265 11381
rect 2291 11355 2317 11381
rect 2343 11355 2369 11381
rect 17599 11355 17625 11381
rect 17651 11355 17677 11381
rect 17703 11355 17729 11381
rect 10991 11271 11017 11297
rect 11663 11271 11689 11297
rect 967 11215 993 11241
rect 9423 11215 9449 11241
rect 10823 11215 10849 11241
rect 13231 11215 13257 11241
rect 14295 11215 14321 11241
rect 20007 11215 20033 11241
rect 2143 11159 2169 11185
rect 7015 11159 7041 11185
rect 7127 11159 7153 11185
rect 7351 11159 7377 11185
rect 7407 11159 7433 11185
rect 7631 11159 7657 11185
rect 9647 11159 9673 11185
rect 10767 11159 10793 11185
rect 11663 11159 11689 11185
rect 12839 11159 12865 11185
rect 18831 11159 18857 11185
rect 6847 11103 6873 11129
rect 11831 11103 11857 11129
rect 11943 11103 11969 11129
rect 6903 11047 6929 11073
rect 7519 11047 7545 11073
rect 9815 11047 9841 11073
rect 9983 11047 10009 11073
rect 11551 11047 11577 11073
rect 9919 10963 9945 10989
rect 9971 10963 9997 10989
rect 10023 10963 10049 10989
rect 7519 10879 7545 10905
rect 10767 10879 10793 10905
rect 6735 10823 6761 10849
rect 7463 10823 7489 10849
rect 8191 10823 8217 10849
rect 14911 10823 14937 10849
rect 7071 10767 7097 10793
rect 7575 10767 7601 10793
rect 7743 10767 7769 10793
rect 8135 10767 8161 10793
rect 8975 10767 9001 10793
rect 9759 10767 9785 10793
rect 10151 10767 10177 10793
rect 10375 10767 10401 10793
rect 10599 10767 10625 10793
rect 10935 10767 10961 10793
rect 13175 10767 13201 10793
rect 14799 10767 14825 10793
rect 18831 10767 18857 10793
rect 5671 10711 5697 10737
rect 8751 10711 8777 10737
rect 9199 10711 9225 10737
rect 9647 10711 9673 10737
rect 11271 10711 11297 10737
rect 12335 10711 12361 10737
rect 13511 10711 13537 10737
rect 14575 10711 14601 10737
rect 20007 10711 20033 10737
rect 9927 10655 9953 10681
rect 2239 10571 2265 10597
rect 2291 10571 2317 10597
rect 2343 10571 2369 10597
rect 17599 10571 17625 10597
rect 17651 10571 17677 10597
rect 17703 10571 17729 10597
rect 20007 10431 20033 10457
rect 10039 10375 10065 10401
rect 11327 10375 11353 10401
rect 11663 10375 11689 10401
rect 18831 10375 18857 10401
rect 8135 10319 8161 10345
rect 10655 10319 10681 10345
rect 11047 10319 11073 10345
rect 13175 10319 13201 10345
rect 10711 10263 10737 10289
rect 11327 10263 11353 10289
rect 9919 10179 9945 10205
rect 9971 10179 9997 10205
rect 10023 10179 10049 10205
rect 7799 10039 7825 10065
rect 8919 10039 8945 10065
rect 8975 10039 9001 10065
rect 9031 10039 9057 10065
rect 9535 10039 9561 10065
rect 11663 10039 11689 10065
rect 12783 10039 12809 10065
rect 13287 10039 13313 10065
rect 13791 10039 13817 10065
rect 13847 10039 13873 10065
rect 8135 9983 8161 10009
rect 9423 9983 9449 10009
rect 9703 9983 9729 10009
rect 12671 9983 12697 10009
rect 13231 9983 13257 10009
rect 13343 9983 13369 10009
rect 13567 9983 13593 10009
rect 18943 9983 18969 10009
rect 6735 9927 6761 9953
rect 20007 9927 20033 9953
rect 9479 9871 9505 9897
rect 13847 9871 13873 9897
rect 2239 9787 2265 9813
rect 2291 9787 2317 9813
rect 2343 9787 2369 9813
rect 17599 9787 17625 9813
rect 17651 9787 17677 9813
rect 17703 9787 17729 9813
rect 10263 9703 10289 9729
rect 12055 9703 12081 9729
rect 20007 9703 20033 9729
rect 8415 9647 8441 9673
rect 9311 9647 9337 9673
rect 9647 9647 9673 9673
rect 12279 9647 12305 9673
rect 12503 9647 12529 9673
rect 7015 9591 7041 9617
rect 9423 9591 9449 9617
rect 9983 9591 10009 9617
rect 10095 9591 10121 9617
rect 10991 9591 11017 9617
rect 11103 9591 11129 9617
rect 11327 9591 11353 9617
rect 11439 9591 11465 9617
rect 11943 9591 11969 9617
rect 13679 9591 13705 9617
rect 13847 9591 13873 9617
rect 14575 9591 14601 9617
rect 18831 9591 18857 9617
rect 7351 9535 7377 9561
rect 10823 9535 10849 9561
rect 12223 9535 12249 9561
rect 12335 9535 12361 9561
rect 12895 9535 12921 9561
rect 13511 9535 13537 9561
rect 9927 9479 9953 9505
rect 10039 9479 10065 9505
rect 11271 9479 11297 9505
rect 12559 9479 12585 9505
rect 12615 9479 12641 9505
rect 13063 9479 13089 9505
rect 13735 9479 13761 9505
rect 14743 9479 14769 9505
rect 9919 9395 9945 9421
rect 9971 9395 9997 9421
rect 10023 9395 10049 9421
rect 7575 9311 7601 9337
rect 9199 9311 9225 9337
rect 9703 9311 9729 9337
rect 11663 9311 11689 9337
rect 12895 9311 12921 9337
rect 14855 9311 14881 9337
rect 7687 9255 7713 9281
rect 7911 9255 7937 9281
rect 7967 9255 7993 9281
rect 9031 9255 9057 9281
rect 9927 9255 9953 9281
rect 11215 9255 11241 9281
rect 13063 9255 13089 9281
rect 15359 9255 15385 9281
rect 2143 9199 2169 9225
rect 7183 9199 7209 9225
rect 7351 9199 7377 9225
rect 7799 9199 7825 9225
rect 9535 9199 9561 9225
rect 9871 9199 9897 9225
rect 10935 9199 10961 9225
rect 13231 9199 13257 9225
rect 15023 9199 15049 9225
rect 15191 9199 15217 9225
rect 18831 9199 18857 9225
rect 5783 9143 5809 9169
rect 6847 9143 6873 9169
rect 7631 9143 7657 9169
rect 13623 9143 13649 9169
rect 14687 9143 14713 9169
rect 20007 9143 20033 9169
rect 967 9087 993 9113
rect 2239 9003 2265 9029
rect 2291 9003 2317 9029
rect 2343 9003 2369 9029
rect 17599 9003 17625 9029
rect 17651 9003 17677 9029
rect 17703 9003 17729 9029
rect 8863 8919 8889 8945
rect 14071 8919 14097 8945
rect 967 8863 993 8889
rect 9871 8863 9897 8889
rect 12223 8863 12249 8889
rect 13287 8863 13313 8889
rect 14127 8863 14153 8889
rect 19951 8863 19977 8889
rect 2143 8807 2169 8833
rect 6847 8807 6873 8833
rect 6959 8807 6985 8833
rect 7351 8807 7377 8833
rect 9255 8807 9281 8833
rect 9647 8807 9673 8833
rect 10095 8807 10121 8833
rect 10431 8807 10457 8833
rect 10711 8807 10737 8833
rect 11831 8807 11857 8833
rect 14575 8807 14601 8833
rect 18831 8807 18857 8833
rect 7463 8751 7489 8777
rect 7519 8751 7545 8777
rect 8919 8751 8945 8777
rect 9367 8751 9393 8777
rect 10207 8751 10233 8777
rect 6903 8695 6929 8721
rect 7071 8695 7097 8721
rect 8863 8695 8889 8721
rect 9479 8695 9505 8721
rect 9535 8695 9561 8721
rect 10151 8695 10177 8721
rect 10823 8695 10849 8721
rect 14743 8695 14769 8721
rect 9919 8611 9945 8637
rect 9971 8611 9997 8637
rect 10023 8611 10049 8637
rect 7575 8527 7601 8553
rect 7687 8527 7713 8553
rect 9535 8527 9561 8553
rect 11047 8527 11073 8553
rect 7071 8471 7097 8497
rect 7743 8471 7769 8497
rect 8303 8471 8329 8497
rect 8359 8471 8385 8497
rect 9031 8471 9057 8497
rect 10935 8471 10961 8497
rect 11383 8471 11409 8497
rect 19671 8471 19697 8497
rect 7463 8415 7489 8441
rect 8471 8415 8497 8441
rect 8919 8415 8945 8441
rect 9199 8415 9225 8441
rect 9591 8415 9617 8441
rect 9703 8415 9729 8441
rect 9927 8415 9953 8441
rect 9983 8415 10009 8441
rect 11103 8415 11129 8441
rect 11159 8415 11185 8441
rect 11551 8415 11577 8441
rect 18831 8415 18857 8441
rect 6007 8359 6033 8385
rect 9311 8359 9337 8385
rect 9815 8359 9841 8385
rect 11439 8359 11465 8385
rect 8975 8303 9001 8329
rect 2239 8219 2265 8245
rect 2291 8219 2317 8245
rect 2343 8219 2369 8245
rect 17599 8219 17625 8245
rect 17651 8219 17677 8245
rect 17703 8219 17729 8245
rect 7239 8079 7265 8105
rect 8303 8079 8329 8105
rect 8863 8079 8889 8105
rect 9927 8079 9953 8105
rect 11159 8079 11185 8105
rect 12223 8079 12249 8105
rect 19895 8079 19921 8105
rect 6903 8023 6929 8049
rect 8527 8023 8553 8049
rect 10823 8023 10849 8049
rect 18831 8023 18857 8049
rect 9919 7827 9945 7853
rect 9971 7827 9997 7853
rect 10023 7827 10049 7853
rect 9815 7687 9841 7713
rect 11887 7687 11913 7713
rect 9423 7631 9449 7657
rect 11775 7631 11801 7657
rect 18831 7631 18857 7657
rect 10879 7575 10905 7601
rect 20007 7575 20033 7601
rect 2239 7435 2265 7461
rect 2291 7435 2317 7461
rect 2343 7435 2369 7461
rect 17599 7435 17625 7461
rect 17651 7435 17677 7461
rect 17703 7435 17729 7461
rect 9919 7043 9945 7069
rect 9971 7043 9997 7069
rect 10023 7043 10049 7069
rect 2239 6651 2265 6677
rect 2291 6651 2317 6677
rect 2343 6651 2369 6677
rect 17599 6651 17625 6677
rect 17651 6651 17677 6677
rect 17703 6651 17729 6677
rect 9919 6259 9945 6285
rect 9971 6259 9997 6285
rect 10023 6259 10049 6285
rect 2239 5867 2265 5893
rect 2291 5867 2317 5893
rect 2343 5867 2369 5893
rect 17599 5867 17625 5893
rect 17651 5867 17677 5893
rect 17703 5867 17729 5893
rect 9919 5475 9945 5501
rect 9971 5475 9997 5501
rect 10023 5475 10049 5501
rect 2239 5083 2265 5109
rect 2291 5083 2317 5109
rect 2343 5083 2369 5109
rect 17599 5083 17625 5109
rect 17651 5083 17677 5109
rect 17703 5083 17729 5109
rect 9919 4691 9945 4717
rect 9971 4691 9997 4717
rect 10023 4691 10049 4717
rect 2239 4299 2265 4325
rect 2291 4299 2317 4325
rect 2343 4299 2369 4325
rect 17599 4299 17625 4325
rect 17651 4299 17677 4325
rect 17703 4299 17729 4325
rect 9919 3907 9945 3933
rect 9971 3907 9997 3933
rect 10023 3907 10049 3933
rect 2239 3515 2265 3541
rect 2291 3515 2317 3541
rect 2343 3515 2369 3541
rect 17599 3515 17625 3541
rect 17651 3515 17677 3541
rect 17703 3515 17729 3541
rect 9919 3123 9945 3149
rect 9971 3123 9997 3149
rect 10023 3123 10049 3149
rect 2239 2731 2265 2757
rect 2291 2731 2317 2757
rect 2343 2731 2369 2757
rect 17599 2731 17625 2757
rect 17651 2731 17677 2757
rect 17703 2731 17729 2757
rect 12391 2591 12417 2617
rect 11887 2535 11913 2561
rect 9919 2339 9945 2365
rect 9971 2339 9997 2365
rect 10023 2339 10049 2365
rect 2239 1947 2265 1973
rect 2291 1947 2317 1973
rect 2343 1947 2369 1973
rect 17599 1947 17625 1973
rect 17651 1947 17677 1973
rect 17703 1947 17729 1973
rect 9311 1807 9337 1833
rect 11047 1807 11073 1833
rect 12783 1807 12809 1833
rect 8807 1751 8833 1777
rect 10543 1751 10569 1777
rect 12279 1751 12305 1777
rect 9919 1555 9945 1581
rect 9971 1555 9997 1581
rect 10023 1555 10049 1581
<< metal2 >>
rect 8400 20600 8456 21000
rect 11760 20600 11816 21000
rect 12096 20600 12152 21000
rect 12432 20600 12488 21000
rect 2238 19222 2370 19227
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2238 19189 2370 19194
rect 8414 18970 8442 20600
rect 11774 19138 11802 20600
rect 11774 19105 11802 19110
rect 8526 18970 8554 18975
rect 8414 18969 8554 18970
rect 8414 18943 8527 18969
rect 8553 18943 8554 18969
rect 8414 18942 8554 18943
rect 8526 18937 8554 18942
rect 9918 18830 10050 18835
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 9918 18797 10050 18802
rect 12110 18746 12138 20600
rect 12446 19922 12474 20600
rect 12446 19894 12530 19922
rect 12110 18713 12138 18718
rect 12446 19025 12474 19031
rect 12446 18999 12447 19025
rect 12473 18999 12474 19025
rect 2238 18438 2370 18443
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2238 18405 2370 18410
rect 9918 18046 10050 18051
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 9918 18013 10050 18018
rect 2238 17654 2370 17659
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2238 17621 2370 17626
rect 9918 17262 10050 17267
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 9918 17229 10050 17234
rect 2238 16870 2370 16875
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2238 16837 2370 16842
rect 9918 16478 10050 16483
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 9918 16445 10050 16450
rect 2238 16086 2370 16091
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2238 16053 2370 16058
rect 9918 15694 10050 15699
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 9918 15661 10050 15666
rect 2238 15302 2370 15307
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2238 15269 2370 15274
rect 9918 14910 10050 14915
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 9918 14877 10050 14882
rect 2238 14518 2370 14523
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2238 14485 2370 14490
rect 9918 14126 10050 14131
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 9918 14093 10050 14098
rect 2238 13734 2370 13739
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2238 13701 2370 13706
rect 12446 13454 12474 18999
rect 12502 18354 12530 19894
rect 17598 19222 17730 19227
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17598 19189 17730 19194
rect 12782 19138 12810 19143
rect 12782 19091 12810 19110
rect 13118 18746 13146 18751
rect 13118 18699 13146 18718
rect 12614 18633 12642 18639
rect 12614 18607 12615 18633
rect 12641 18607 12642 18633
rect 12558 18354 12586 18359
rect 12502 18326 12558 18354
rect 12558 18321 12586 18326
rect 12390 13426 12474 13454
rect 9918 13342 10050 13347
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 9918 13309 10050 13314
rect 7574 13258 7602 13263
rect 7462 13257 7602 13258
rect 7462 13231 7575 13257
rect 7601 13231 7602 13257
rect 7462 13230 7602 13231
rect 2238 12950 2370 12955
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2238 12917 2370 12922
rect 966 12809 994 12815
rect 966 12783 967 12809
rect 993 12783 994 12809
rect 966 12474 994 12783
rect 966 12441 994 12446
rect 2086 12810 2114 12815
rect 966 12250 994 12255
rect 966 12203 994 12222
rect 966 11466 994 11471
rect 966 11419 994 11438
rect 966 11241 994 11247
rect 966 11215 967 11241
rect 993 11215 994 11241
rect 966 10794 994 11215
rect 966 10761 994 10766
rect 2086 9506 2114 12782
rect 6734 12809 6762 12815
rect 6734 12783 6735 12809
rect 6761 12783 6762 12809
rect 2142 12754 2170 12759
rect 2142 12707 2170 12726
rect 6734 12754 6762 12783
rect 6734 12721 6762 12726
rect 7462 12754 7490 13230
rect 7574 13225 7602 13230
rect 12222 13258 12250 13263
rect 12222 13211 12250 13230
rect 7462 12721 7490 12726
rect 7518 13145 7546 13151
rect 7518 13119 7519 13145
rect 7545 13119 7546 13145
rect 7518 12474 7546 13119
rect 12110 13145 12138 13151
rect 12110 13119 12111 13145
rect 12137 13119 12138 13145
rect 7574 13034 7602 13039
rect 7574 13033 7658 13034
rect 7574 13007 7575 13033
rect 7601 13007 7658 13033
rect 7574 13006 7658 13007
rect 7574 13001 7602 13006
rect 7462 12446 7518 12474
rect 2142 12362 2170 12367
rect 2142 12315 2170 12334
rect 6230 12362 6258 12367
rect 6230 12305 6258 12334
rect 6230 12279 6231 12305
rect 6257 12279 6258 12305
rect 6230 12273 6258 12279
rect 7294 12305 7322 12311
rect 7294 12279 7295 12305
rect 7321 12279 7322 12305
rect 2238 12166 2370 12171
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2238 12133 2370 12138
rect 7294 12025 7322 12279
rect 7294 11999 7295 12025
rect 7321 11999 7322 12025
rect 7294 11993 7322 11999
rect 7238 11913 7266 11919
rect 7238 11887 7239 11913
rect 7265 11887 7266 11913
rect 7238 11802 7266 11887
rect 7238 11769 7266 11774
rect 7406 11913 7434 11919
rect 7406 11887 7407 11913
rect 7433 11887 7434 11913
rect 7182 11690 7210 11695
rect 7182 11643 7210 11662
rect 7350 11690 7378 11695
rect 2142 11578 2170 11583
rect 2142 11531 2170 11550
rect 5670 11578 5698 11583
rect 2238 11382 2370 11387
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2238 11349 2370 11354
rect 2142 11186 2170 11191
rect 2142 11139 2170 11158
rect 5670 10737 5698 11550
rect 7294 11578 7322 11583
rect 7294 11531 7322 11550
rect 7238 11521 7266 11527
rect 7238 11495 7239 11521
rect 7265 11495 7266 11521
rect 6734 11186 6762 11191
rect 7014 11186 7042 11191
rect 6734 10962 6762 11158
rect 6846 11158 6986 11186
rect 6846 11129 6874 11158
rect 6846 11103 6847 11129
rect 6873 11103 6874 11129
rect 6846 11097 6874 11103
rect 5670 10711 5671 10737
rect 5697 10711 5698 10737
rect 5670 10705 5698 10711
rect 6678 10934 6762 10962
rect 6902 11073 6930 11079
rect 6902 11047 6903 11073
rect 6929 11047 6930 11073
rect 6678 10738 6706 10934
rect 6902 10906 6930 11047
rect 6734 10878 6930 10906
rect 6734 10849 6762 10878
rect 6734 10823 6735 10849
rect 6761 10823 6762 10849
rect 6734 10817 6762 10823
rect 6790 10738 6818 10743
rect 6678 10710 6790 10738
rect 2238 10598 2370 10603
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2238 10565 2370 10570
rect 6790 10094 6818 10710
rect 6958 10094 6986 11158
rect 7014 11139 7042 11158
rect 7126 11186 7154 11191
rect 7238 11186 7266 11495
rect 7350 11298 7378 11662
rect 7126 11185 7266 11186
rect 7126 11159 7127 11185
rect 7153 11159 7266 11185
rect 7126 11158 7266 11159
rect 7294 11270 7378 11298
rect 7406 11634 7434 11887
rect 7126 11153 7154 11158
rect 7294 10850 7322 11270
rect 7350 11185 7378 11191
rect 7350 11159 7351 11185
rect 7377 11159 7378 11185
rect 7350 10962 7378 11159
rect 7406 11186 7434 11606
rect 7462 11577 7490 12446
rect 7518 12441 7546 12446
rect 7518 12306 7546 12311
rect 7518 11969 7546 12278
rect 7518 11943 7519 11969
rect 7545 11943 7546 11969
rect 7518 11937 7546 11943
rect 7630 11969 7658 13006
rect 10094 12810 10122 12815
rect 10094 12809 10458 12810
rect 10094 12783 10095 12809
rect 10121 12783 10458 12809
rect 10094 12782 10458 12783
rect 10094 12777 10122 12782
rect 8190 12753 8218 12759
rect 8190 12727 8191 12753
rect 8217 12727 8218 12753
rect 7798 12698 7826 12703
rect 7742 12697 7826 12698
rect 7742 12671 7799 12697
rect 7825 12671 7826 12697
rect 7742 12670 7826 12671
rect 7686 12361 7714 12367
rect 7686 12335 7687 12361
rect 7713 12335 7714 12361
rect 7686 12026 7714 12335
rect 7742 12026 7770 12670
rect 7798 12665 7826 12670
rect 8078 12474 8106 12479
rect 8078 12427 8106 12446
rect 7966 12418 7994 12423
rect 7966 12371 7994 12390
rect 7854 12361 7882 12367
rect 7854 12335 7855 12361
rect 7881 12335 7882 12361
rect 7854 12138 7882 12335
rect 7910 12306 7938 12311
rect 7910 12259 7938 12278
rect 7854 12110 7994 12138
rect 7742 11998 7826 12026
rect 7686 11993 7714 11998
rect 7630 11943 7631 11969
rect 7657 11943 7658 11969
rect 7630 11937 7658 11943
rect 7798 11857 7826 11998
rect 7854 11970 7882 11975
rect 7854 11923 7882 11942
rect 7910 11969 7938 11975
rect 7910 11943 7911 11969
rect 7937 11943 7938 11969
rect 7798 11831 7799 11857
rect 7825 11831 7826 11857
rect 7798 11825 7826 11831
rect 7462 11551 7463 11577
rect 7489 11551 7490 11577
rect 7462 11545 7490 11551
rect 7686 11690 7714 11695
rect 7686 11577 7714 11662
rect 7798 11634 7826 11639
rect 7910 11634 7938 11943
rect 7966 11690 7994 12110
rect 8190 12026 8218 12727
rect 8694 12753 8722 12759
rect 8694 12727 8695 12753
rect 8721 12727 8722 12753
rect 8358 12474 8386 12479
rect 8358 12427 8386 12446
rect 8638 12474 8666 12479
rect 8190 11993 8218 11998
rect 8302 12361 8330 12367
rect 8302 12335 8303 12361
rect 8329 12335 8330 12361
rect 8302 11802 8330 12335
rect 8470 12362 8498 12367
rect 8470 12315 8498 12334
rect 8302 11769 8330 11774
rect 8414 12026 8442 12031
rect 7966 11657 7994 11662
rect 7826 11606 7938 11634
rect 7798 11587 7826 11606
rect 7686 11551 7687 11577
rect 7713 11551 7714 11577
rect 7686 11545 7714 11551
rect 7406 11139 7434 11158
rect 7630 11185 7658 11191
rect 7630 11159 7631 11185
rect 7657 11159 7658 11185
rect 7518 11073 7546 11079
rect 7518 11047 7519 11073
rect 7545 11047 7546 11073
rect 7518 11018 7546 11047
rect 7518 10990 7602 11018
rect 7350 10934 7546 10962
rect 7518 10905 7546 10934
rect 7518 10879 7519 10905
rect 7545 10879 7546 10905
rect 7518 10873 7546 10879
rect 7574 10906 7602 10990
rect 7630 10962 7658 11159
rect 7630 10934 7882 10962
rect 7574 10878 7826 10906
rect 7462 10850 7490 10855
rect 7294 10849 7490 10850
rect 7294 10823 7463 10849
rect 7489 10823 7490 10849
rect 7294 10822 7490 10823
rect 7070 10793 7098 10799
rect 7070 10767 7071 10793
rect 7097 10767 7098 10793
rect 7070 10094 7098 10767
rect 7462 10794 7490 10822
rect 7462 10761 7490 10766
rect 7574 10793 7602 10799
rect 7574 10767 7575 10793
rect 7601 10767 7602 10793
rect 7574 10738 7602 10767
rect 7574 10705 7602 10710
rect 7742 10793 7770 10799
rect 7742 10767 7743 10793
rect 7769 10767 7770 10793
rect 7742 10738 7770 10767
rect 7742 10705 7770 10710
rect 6734 10066 6818 10094
rect 6902 10066 6986 10094
rect 7014 10066 7098 10094
rect 6734 9953 6762 10066
rect 6734 9927 6735 9953
rect 6761 9927 6762 9953
rect 6734 9921 6762 9927
rect 2238 9814 2370 9819
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2238 9781 2370 9786
rect 2086 9473 2114 9478
rect 2142 9225 2170 9231
rect 2142 9199 2143 9225
rect 2169 9199 2170 9225
rect 2142 9170 2170 9199
rect 2142 9137 2170 9142
rect 5782 9170 5810 9175
rect 966 9114 994 9119
rect 966 9067 994 9086
rect 2238 9030 2370 9035
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2238 8997 2370 9002
rect 966 8889 994 8895
rect 966 8863 967 8889
rect 993 8863 994 8889
rect 966 8442 994 8863
rect 2142 8834 2170 8839
rect 2142 8787 2170 8806
rect 5782 8778 5810 9142
rect 6846 9170 6874 9175
rect 6846 9123 6874 9142
rect 6902 9114 6930 10066
rect 7014 10010 7042 10066
rect 7798 10065 7826 10878
rect 7798 10039 7799 10065
rect 7825 10039 7826 10065
rect 7798 10033 7826 10039
rect 7014 9617 7042 9982
rect 7854 9954 7882 10934
rect 8190 10849 8218 10855
rect 8190 10823 8191 10849
rect 8217 10823 8218 10849
rect 8134 10794 8162 10799
rect 8190 10794 8218 10823
rect 8246 10794 8274 10799
rect 8190 10766 8246 10794
rect 8134 10747 8162 10766
rect 8246 10761 8274 10766
rect 8134 10346 8162 10351
rect 8134 10010 8162 10318
rect 8414 10346 8442 11998
rect 8638 11914 8666 12446
rect 8694 12361 8722 12727
rect 9030 12698 9058 12703
rect 8694 12335 8695 12361
rect 8721 12335 8722 12361
rect 8694 12026 8722 12335
rect 8694 11993 8722 11998
rect 8918 12697 9058 12698
rect 8918 12671 9031 12697
rect 9057 12671 9058 12697
rect 8918 12670 9058 12671
rect 8694 11914 8722 11919
rect 8638 11913 8722 11914
rect 8638 11887 8695 11913
rect 8721 11887 8722 11913
rect 8638 11886 8722 11887
rect 8694 11881 8722 11886
rect 8862 11857 8890 11863
rect 8862 11831 8863 11857
rect 8889 11831 8890 11857
rect 8414 10313 8442 10318
rect 8750 11802 8778 11807
rect 8750 10737 8778 11774
rect 8862 11578 8890 11831
rect 8862 11545 8890 11550
rect 8750 10711 8751 10737
rect 8777 10711 8778 10737
rect 8134 9963 8162 9982
rect 7966 9954 7994 9959
rect 7854 9926 7966 9954
rect 7014 9591 7015 9617
rect 7041 9591 7042 9617
rect 5782 8745 5810 8750
rect 6006 8834 6034 8839
rect 966 8409 994 8414
rect 6006 8554 6034 8806
rect 6846 8834 6874 8839
rect 6902 8834 6930 9086
rect 6846 8833 6930 8834
rect 6846 8807 6847 8833
rect 6873 8807 6930 8833
rect 6846 8806 6930 8807
rect 6958 9338 6986 9343
rect 6958 8833 6986 9310
rect 7014 9226 7042 9591
rect 7350 9562 7378 9567
rect 7350 9561 7434 9562
rect 7350 9535 7351 9561
rect 7377 9535 7434 9561
rect 7350 9534 7434 9535
rect 7350 9529 7378 9534
rect 7182 9226 7210 9231
rect 7014 9225 7210 9226
rect 7014 9199 7183 9225
rect 7209 9199 7210 9225
rect 7014 9198 7210 9199
rect 6958 8807 6959 8833
rect 6985 8807 6986 8833
rect 6846 8801 6874 8806
rect 6958 8801 6986 8807
rect 6902 8721 6930 8727
rect 6902 8695 6903 8721
rect 6929 8695 6930 8721
rect 6902 8554 6930 8695
rect 7070 8722 7098 8727
rect 7070 8675 7098 8694
rect 6902 8526 7098 8554
rect 6006 8385 6034 8526
rect 7070 8497 7098 8526
rect 7070 8471 7071 8497
rect 7097 8471 7098 8497
rect 7070 8465 7098 8471
rect 6006 8359 6007 8385
rect 6033 8359 6034 8385
rect 6006 8353 6034 8359
rect 2238 8246 2370 8251
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2238 8213 2370 8218
rect 6902 8050 6930 8055
rect 6902 8003 6930 8022
rect 7182 8050 7210 9198
rect 7350 9225 7378 9231
rect 7350 9199 7351 9225
rect 7377 9199 7378 9225
rect 7350 8833 7378 9199
rect 7406 9226 7434 9534
rect 7574 9338 7602 9343
rect 7574 9291 7602 9310
rect 7686 9282 7714 9287
rect 7686 9235 7714 9254
rect 7910 9281 7938 9287
rect 7910 9255 7911 9281
rect 7937 9255 7938 9281
rect 7406 9193 7434 9198
rect 7798 9226 7826 9231
rect 7798 9179 7826 9198
rect 7630 9170 7658 9175
rect 7630 9123 7658 9142
rect 7910 9114 7938 9255
rect 7966 9282 7994 9926
rect 8750 9898 8778 10711
rect 8918 10514 8946 12670
rect 9030 12665 9058 12670
rect 9918 12558 10050 12563
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 9918 12525 10050 12530
rect 8974 12362 9002 12367
rect 9758 12362 9786 12367
rect 10430 12362 10458 12782
rect 10990 12753 11018 12759
rect 10990 12727 10991 12753
rect 11017 12727 11018 12753
rect 10990 12474 11018 12727
rect 11326 12698 11354 12703
rect 11158 12697 11354 12698
rect 11158 12671 11327 12697
rect 11353 12671 11354 12697
rect 11158 12670 11354 12671
rect 10990 12446 11130 12474
rect 11046 12362 11074 12367
rect 9002 12334 9058 12362
rect 8974 12329 9002 12334
rect 9030 11969 9058 12334
rect 9086 12306 9114 12311
rect 9086 12305 9226 12306
rect 9086 12279 9087 12305
rect 9113 12279 9226 12305
rect 9086 12278 9226 12279
rect 9086 12273 9114 12278
rect 9198 12026 9226 12278
rect 9702 12082 9730 12087
rect 9254 12026 9282 12031
rect 9198 12025 9282 12026
rect 9198 11999 9255 12025
rect 9281 11999 9282 12025
rect 9198 11998 9282 11999
rect 9254 11993 9282 11998
rect 9030 11943 9031 11969
rect 9057 11943 9058 11969
rect 9030 11937 9058 11943
rect 9310 11970 9338 11975
rect 9310 11923 9338 11942
rect 9198 11914 9226 11919
rect 9198 11867 9226 11886
rect 9366 11690 9394 11695
rect 9366 11643 9394 11662
rect 9702 11689 9730 12054
rect 9702 11663 9703 11689
rect 9729 11663 9730 11689
rect 9702 11657 9730 11663
rect 9758 11914 9786 12334
rect 10374 12361 10458 12362
rect 10374 12335 10431 12361
rect 10457 12335 10458 12361
rect 10374 12334 10458 12335
rect 10150 12306 10178 12311
rect 10318 12306 10346 12311
rect 10150 12305 10346 12306
rect 10150 12279 10151 12305
rect 10177 12279 10319 12305
rect 10345 12279 10346 12305
rect 10150 12278 10346 12279
rect 10150 12082 10178 12278
rect 10318 12273 10346 12278
rect 10150 12049 10178 12054
rect 9534 11633 9562 11639
rect 9534 11607 9535 11633
rect 9561 11607 9562 11633
rect 9310 11578 9338 11583
rect 9534 11578 9562 11607
rect 9338 11550 9562 11578
rect 9758 11578 9786 11886
rect 10094 11969 10122 11975
rect 10094 11943 10095 11969
rect 10121 11943 10122 11969
rect 9926 11858 9954 11863
rect 10094 11858 10122 11943
rect 10374 11969 10402 12334
rect 10430 12329 10458 12334
rect 10934 12361 11074 12362
rect 10934 12335 11047 12361
rect 11073 12335 11074 12361
rect 10934 12334 11074 12335
rect 10598 12250 10626 12255
rect 10598 12249 10682 12250
rect 10598 12223 10599 12249
rect 10625 12223 10682 12249
rect 10598 12222 10682 12223
rect 10598 12217 10626 12222
rect 10374 11943 10375 11969
rect 10401 11943 10402 11969
rect 10374 11937 10402 11943
rect 10542 12194 10570 12199
rect 10542 11970 10570 12166
rect 9926 11857 10122 11858
rect 9926 11831 9927 11857
rect 9953 11831 10122 11857
rect 9926 11830 10122 11831
rect 9926 11825 9954 11830
rect 9918 11774 10050 11779
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 9918 11741 10050 11746
rect 9926 11690 9954 11695
rect 9926 11643 9954 11662
rect 9982 11578 10010 11583
rect 9758 11577 10010 11578
rect 9758 11551 9983 11577
rect 10009 11551 10010 11577
rect 9758 11550 10010 11551
rect 9310 11531 9338 11550
rect 9422 11241 9450 11247
rect 9422 11215 9423 11241
rect 9449 11215 9450 11241
rect 8974 10794 9002 10799
rect 8974 10747 9002 10766
rect 9198 10738 9226 10743
rect 9030 10737 9226 10738
rect 9030 10711 9199 10737
rect 9225 10711 9226 10737
rect 9030 10710 9226 10711
rect 8918 10486 9002 10514
rect 8750 9865 8778 9870
rect 8918 10065 8946 10071
rect 8918 10039 8919 10065
rect 8945 10039 8946 10065
rect 8414 9674 8442 9679
rect 8414 9627 8442 9646
rect 7966 9235 7994 9254
rect 8918 9562 8946 10039
rect 8974 10065 9002 10486
rect 8974 10039 8975 10065
rect 9001 10039 9002 10065
rect 8974 10033 9002 10039
rect 9030 10065 9058 10710
rect 9198 10705 9226 10710
rect 9422 10738 9450 11215
rect 9534 11186 9562 11550
rect 9982 11545 10010 11550
rect 9926 11466 9954 11471
rect 9702 11465 9954 11466
rect 9702 11439 9927 11465
rect 9953 11439 9954 11465
rect 9702 11438 9954 11439
rect 9646 11186 9674 11191
rect 9534 11158 9646 11186
rect 9646 11139 9674 11158
rect 9646 10738 9674 10743
rect 9450 10737 9674 10738
rect 9450 10711 9647 10737
rect 9673 10711 9674 10737
rect 9450 10710 9674 10711
rect 9422 10691 9450 10710
rect 9646 10122 9674 10710
rect 9702 10402 9730 11438
rect 9926 11433 9954 11438
rect 9814 11074 9842 11079
rect 9758 11073 9842 11074
rect 9758 11047 9815 11073
rect 9841 11047 9842 11073
rect 9758 11046 9842 11047
rect 9758 10794 9786 11046
rect 9814 11041 9842 11046
rect 9982 11074 10010 11079
rect 10094 11074 10122 11830
rect 10318 11718 10514 11746
rect 10318 11633 10346 11718
rect 10430 11634 10458 11639
rect 10318 11607 10319 11633
rect 10345 11607 10346 11633
rect 10318 11601 10346 11607
rect 10374 11633 10458 11634
rect 10374 11607 10431 11633
rect 10457 11607 10458 11633
rect 10374 11606 10458 11607
rect 9982 11073 10122 11074
rect 9982 11047 9983 11073
rect 10009 11047 10122 11073
rect 9982 11046 10122 11047
rect 9982 11041 10010 11046
rect 9918 10990 10050 10995
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 9918 10957 10050 10962
rect 10094 10850 10122 11046
rect 10094 10817 10122 10822
rect 9758 10747 9786 10766
rect 10150 10794 10178 10799
rect 10150 10747 10178 10766
rect 10374 10793 10402 11606
rect 10430 11601 10458 11606
rect 10374 10767 10375 10793
rect 10401 10767 10402 10793
rect 9926 10681 9954 10687
rect 9926 10655 9927 10681
rect 9953 10655 9954 10681
rect 9702 10374 9842 10402
rect 9646 10089 9674 10094
rect 9758 10290 9786 10295
rect 9030 10039 9031 10065
rect 9057 10039 9058 10065
rect 9030 10033 9058 10039
rect 9534 10066 9562 10071
rect 9534 10065 9618 10066
rect 9534 10039 9535 10065
rect 9561 10039 9618 10065
rect 9534 10038 9618 10039
rect 9534 10033 9562 10038
rect 8918 9282 8946 9534
rect 9310 10010 9338 10015
rect 9310 9673 9338 9982
rect 9310 9647 9311 9673
rect 9337 9647 9338 9673
rect 9310 9506 9338 9647
rect 9422 10009 9450 10015
rect 9422 9983 9423 10009
rect 9449 9983 9450 10009
rect 9422 9674 9450 9983
rect 9422 9618 9450 9646
rect 9310 9473 9338 9478
rect 9366 9617 9450 9618
rect 9366 9591 9423 9617
rect 9449 9591 9450 9617
rect 9366 9590 9450 9591
rect 9366 9394 9394 9590
rect 9422 9585 9450 9590
rect 9478 9898 9506 9903
rect 9478 9506 9506 9870
rect 9478 9473 9506 9478
rect 9534 9730 9562 9735
rect 9198 9366 9394 9394
rect 9198 9337 9226 9366
rect 9422 9338 9450 9343
rect 9534 9338 9562 9702
rect 9198 9311 9199 9337
rect 9225 9311 9226 9337
rect 9198 9305 9226 9311
rect 9310 9310 9422 9338
rect 9450 9310 9562 9338
rect 8918 9249 8946 9254
rect 9030 9281 9058 9287
rect 9030 9255 9031 9281
rect 9057 9255 9058 9281
rect 7910 8946 7938 9086
rect 7910 8913 7938 8918
rect 8862 8946 8890 8951
rect 8862 8899 8890 8918
rect 7350 8807 7351 8833
rect 7377 8807 7378 8833
rect 7350 8801 7378 8807
rect 7462 8778 7490 8783
rect 7462 8731 7490 8750
rect 7518 8777 7546 8783
rect 7518 8751 7519 8777
rect 7545 8751 7546 8777
rect 7518 8666 7546 8751
rect 8918 8778 8946 8783
rect 9030 8778 9058 9255
rect 9254 9282 9282 9287
rect 8946 8750 9058 8778
rect 9086 8834 9114 8839
rect 8918 8731 8946 8750
rect 7518 8633 7546 8638
rect 7574 8722 7602 8727
rect 7574 8553 7602 8694
rect 8862 8722 8890 8727
rect 7574 8527 7575 8553
rect 7601 8527 7602 8553
rect 7574 8521 7602 8527
rect 7686 8554 7714 8559
rect 7686 8507 7714 8526
rect 7742 8498 7770 8503
rect 7742 8451 7770 8470
rect 8302 8498 8330 8503
rect 8302 8451 8330 8470
rect 8358 8497 8386 8503
rect 8358 8471 8359 8497
rect 8385 8471 8386 8497
rect 7462 8442 7490 8447
rect 7462 8441 7546 8442
rect 7462 8415 7463 8441
rect 7489 8415 7546 8441
rect 7462 8414 7546 8415
rect 7462 8409 7490 8414
rect 7238 8330 7266 8335
rect 7238 8105 7266 8302
rect 7238 8079 7239 8105
rect 7265 8079 7266 8105
rect 7238 8073 7266 8079
rect 7182 8017 7210 8022
rect 7518 8050 7546 8414
rect 8302 8106 8330 8111
rect 8358 8106 8386 8471
rect 8470 8442 8498 8447
rect 8470 8395 8498 8414
rect 8330 8078 8386 8106
rect 8806 8106 8834 8111
rect 8302 8059 8330 8078
rect 7518 8017 7546 8022
rect 8526 8050 8554 8055
rect 8526 7658 8554 8022
rect 8526 7625 8554 7630
rect 2238 7462 2370 7467
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2238 7429 2370 7434
rect 2238 6678 2370 6683
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2238 6645 2370 6650
rect 2238 5894 2370 5899
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2238 5861 2370 5866
rect 2238 5110 2370 5115
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2238 5077 2370 5082
rect 2238 4326 2370 4331
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2238 4293 2370 4298
rect 2238 3542 2370 3547
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2238 3509 2370 3514
rect 2238 2758 2370 2763
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2238 2725 2370 2730
rect 2238 1974 2370 1979
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2238 1941 2370 1946
rect 8806 1777 8834 8078
rect 8862 8105 8890 8694
rect 9030 8498 9058 8503
rect 9086 8498 9114 8806
rect 9254 8833 9282 9254
rect 9254 8807 9255 8833
rect 9281 8807 9282 8833
rect 9254 8801 9282 8807
rect 9030 8497 9114 8498
rect 9030 8471 9031 8497
rect 9057 8471 9114 8497
rect 9030 8470 9114 8471
rect 9198 8778 9226 8783
rect 9030 8465 9058 8470
rect 8918 8442 8946 8447
rect 8918 8395 8946 8414
rect 9198 8441 9226 8750
rect 9198 8415 9199 8441
rect 9225 8415 9226 8441
rect 9198 8409 9226 8415
rect 9310 8385 9338 9310
rect 9422 9291 9450 9310
rect 9590 9282 9618 10038
rect 9702 10010 9730 10015
rect 9702 9963 9730 9982
rect 9646 9673 9674 9679
rect 9646 9647 9647 9673
rect 9673 9647 9674 9673
rect 9646 9338 9674 9647
rect 9646 9305 9674 9310
rect 9702 9618 9730 9623
rect 9702 9337 9730 9590
rect 9702 9311 9703 9337
rect 9729 9311 9730 9337
rect 9702 9305 9730 9311
rect 9534 9226 9562 9231
rect 9534 9179 9562 9198
rect 9590 8834 9618 9254
rect 9646 8834 9674 8839
rect 9758 8834 9786 10262
rect 9814 9730 9842 10374
rect 9926 10290 9954 10655
rect 10038 10402 10066 10407
rect 10038 10355 10066 10374
rect 10374 10290 10402 10767
rect 10486 10794 10514 11718
rect 10542 11689 10570 11942
rect 10542 11663 10543 11689
rect 10569 11663 10570 11689
rect 10542 11657 10570 11663
rect 10598 10794 10626 10799
rect 10486 10793 10626 10794
rect 10486 10767 10599 10793
rect 10625 10767 10626 10793
rect 10486 10766 10626 10767
rect 10598 10346 10626 10766
rect 10654 10458 10682 12222
rect 10934 11746 10962 12334
rect 11046 12329 11074 12334
rect 11102 11970 11130 12446
rect 11158 12473 11186 12670
rect 11326 12665 11354 12670
rect 11158 12447 11159 12473
rect 11185 12447 11186 12473
rect 11158 12441 11186 12447
rect 11550 12642 11578 12647
rect 11550 12417 11578 12614
rect 12110 12642 12138 13119
rect 12110 12609 12138 12614
rect 12390 12809 12418 13426
rect 12614 13258 12642 18607
rect 17598 18438 17730 18443
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17598 18405 17730 18410
rect 13062 18354 13090 18359
rect 13062 18307 13090 18326
rect 12614 13225 12642 13230
rect 12670 18241 12698 18247
rect 12670 18215 12671 18241
rect 12697 18215 12698 18241
rect 12390 12783 12391 12809
rect 12417 12783 12418 12809
rect 12390 12642 12418 12783
rect 12670 12697 12698 18215
rect 17598 17654 17730 17659
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17598 17621 17730 17626
rect 17598 16870 17730 16875
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17598 16837 17730 16842
rect 17598 16086 17730 16091
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17598 16053 17730 16058
rect 17598 15302 17730 15307
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17598 15269 17730 15274
rect 17598 14518 17730 14523
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17598 14485 17730 14490
rect 17598 13734 17730 13739
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17598 13701 17730 13706
rect 17598 12950 17730 12955
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17598 12917 17730 12922
rect 12670 12671 12671 12697
rect 12697 12671 12698 12697
rect 12670 12665 12698 12671
rect 12782 12753 12810 12759
rect 12782 12727 12783 12753
rect 12809 12727 12810 12753
rect 12390 12609 12418 12614
rect 12782 12642 12810 12727
rect 12782 12609 12810 12614
rect 11550 12391 11551 12417
rect 11577 12391 11578 12417
rect 11550 12385 11578 12391
rect 11382 12362 11410 12367
rect 11382 12315 11410 12334
rect 11606 12361 11634 12367
rect 11606 12335 11607 12361
rect 11633 12335 11634 12361
rect 11438 12305 11466 12311
rect 11438 12279 11439 12305
rect 11465 12279 11466 12305
rect 11214 12250 11242 12255
rect 11438 12250 11466 12279
rect 11214 12249 11466 12250
rect 11214 12223 11215 12249
rect 11241 12223 11466 12249
rect 11214 12222 11466 12223
rect 11214 12217 11242 12222
rect 11382 11970 11410 11975
rect 11102 11969 11410 11970
rect 11102 11943 11383 11969
rect 11409 11943 11410 11969
rect 11102 11942 11410 11943
rect 10710 11718 10962 11746
rect 10710 11690 10738 11718
rect 10710 11577 10738 11662
rect 10710 11551 10711 11577
rect 10737 11551 10738 11577
rect 10710 11545 10738 11551
rect 10990 11298 11018 11303
rect 10822 11241 10850 11247
rect 10822 11215 10823 11241
rect 10849 11215 10850 11241
rect 10766 11186 10794 11191
rect 10766 11139 10794 11158
rect 10766 10906 10794 10911
rect 10766 10859 10794 10878
rect 10822 10850 10850 11215
rect 10822 10817 10850 10822
rect 10934 10794 10962 10799
rect 10934 10747 10962 10766
rect 10654 10430 10794 10458
rect 10654 10346 10682 10351
rect 10598 10345 10682 10346
rect 10598 10319 10655 10345
rect 10681 10319 10682 10345
rect 10598 10318 10682 10319
rect 9926 10262 10122 10290
rect 9918 10206 10050 10211
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 9918 10173 10050 10178
rect 9814 9697 9842 9702
rect 10038 10122 10066 10127
rect 9982 9618 10010 9623
rect 9422 8833 9730 8834
rect 9422 8807 9647 8833
rect 9673 8807 9730 8833
rect 9422 8806 9730 8807
rect 9366 8778 9394 8783
rect 9366 8731 9394 8750
rect 9422 8442 9450 8806
rect 9646 8801 9674 8806
rect 9478 8722 9506 8727
rect 9478 8554 9506 8694
rect 9534 8722 9562 8727
rect 9534 8721 9674 8722
rect 9534 8695 9535 8721
rect 9561 8695 9674 8721
rect 9534 8694 9674 8695
rect 9534 8689 9562 8694
rect 9646 8610 9674 8694
rect 9702 8666 9730 8806
rect 9758 8801 9786 8806
rect 9814 9617 10010 9618
rect 9814 9591 9983 9617
rect 10009 9591 10010 9617
rect 9814 9590 10010 9591
rect 9702 8638 9786 8666
rect 9646 8582 9730 8610
rect 9534 8554 9562 8559
rect 9478 8553 9562 8554
rect 9478 8527 9535 8553
rect 9561 8527 9562 8553
rect 9478 8526 9562 8527
rect 9534 8521 9562 8526
rect 9590 8442 9618 8447
rect 9422 8441 9618 8442
rect 9422 8415 9591 8441
rect 9617 8415 9618 8441
rect 9422 8414 9618 8415
rect 9590 8409 9618 8414
rect 9702 8441 9730 8582
rect 9758 8498 9786 8638
rect 9814 8554 9842 9590
rect 9982 9585 10010 9590
rect 9926 9506 9954 9525
rect 9926 9473 9954 9478
rect 10038 9506 10066 10094
rect 10094 10010 10122 10262
rect 10374 10257 10402 10262
rect 10094 9730 10122 9982
rect 10262 9730 10290 9735
rect 10094 9702 10178 9730
rect 10094 9618 10122 9623
rect 10094 9571 10122 9590
rect 10038 9505 10122 9506
rect 10038 9479 10039 9505
rect 10065 9479 10122 9505
rect 10038 9478 10122 9479
rect 10038 9473 10066 9478
rect 9918 9422 10050 9427
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 9918 9389 10050 9394
rect 9870 9338 9898 9343
rect 10094 9338 10122 9478
rect 9870 9225 9898 9310
rect 10038 9310 10122 9338
rect 9926 9282 9954 9287
rect 9926 9235 9954 9254
rect 9870 9199 9871 9225
rect 9897 9199 9898 9225
rect 9870 9193 9898 9199
rect 10038 9170 10066 9310
rect 10038 9137 10066 9142
rect 9870 8889 9898 8895
rect 9870 8863 9871 8889
rect 9897 8863 9898 8889
rect 9870 8834 9898 8863
rect 9870 8801 9898 8806
rect 10094 8834 10122 8839
rect 10150 8834 10178 9702
rect 10262 9683 10290 9702
rect 10654 9338 10682 10318
rect 10710 10290 10738 10295
rect 10710 10243 10738 10262
rect 10654 9305 10682 9310
rect 10766 9226 10794 10430
rect 10990 9730 11018 11270
rect 11214 10850 11242 10855
rect 11046 10346 11074 10351
rect 11046 10299 11074 10318
rect 10990 9617 11018 9702
rect 10990 9591 10991 9617
rect 11017 9591 11018 9617
rect 10990 9585 11018 9591
rect 11102 9617 11130 9623
rect 11102 9591 11103 9617
rect 11129 9591 11130 9617
rect 10822 9562 10850 9567
rect 10822 9515 10850 9534
rect 11102 9562 11130 9591
rect 11130 9534 11186 9562
rect 11102 9529 11130 9534
rect 10094 8833 10178 8834
rect 10094 8807 10095 8833
rect 10121 8807 10178 8833
rect 10094 8806 10178 8807
rect 10430 8833 10458 8839
rect 10430 8807 10431 8833
rect 10457 8807 10458 8833
rect 10094 8801 10122 8806
rect 10206 8778 10234 8783
rect 10206 8731 10234 8750
rect 10150 8721 10178 8727
rect 10150 8695 10151 8721
rect 10177 8695 10178 8721
rect 9918 8638 10050 8643
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 9918 8605 10050 8610
rect 9814 8526 10010 8554
rect 9758 8470 9898 8498
rect 9702 8415 9703 8441
rect 9729 8415 9730 8441
rect 9702 8409 9730 8415
rect 9310 8359 9311 8385
rect 9337 8359 9338 8385
rect 9310 8353 9338 8359
rect 9814 8385 9842 8391
rect 9814 8359 9815 8385
rect 9841 8359 9842 8385
rect 8974 8330 9002 8335
rect 8974 8283 9002 8302
rect 8862 8079 8863 8105
rect 8889 8079 8890 8105
rect 8862 8073 8890 8079
rect 9814 7713 9842 8359
rect 9870 8106 9898 8470
rect 9926 8442 9954 8447
rect 9926 8395 9954 8414
rect 9982 8441 10010 8526
rect 9982 8415 9983 8441
rect 10009 8415 10010 8441
rect 9982 8409 10010 8415
rect 10150 8442 10178 8695
rect 10150 8409 10178 8414
rect 9926 8106 9954 8111
rect 9870 8105 9954 8106
rect 9870 8079 9927 8105
rect 9953 8079 9954 8105
rect 9870 8078 9954 8079
rect 9926 8073 9954 8078
rect 9918 7854 10050 7859
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 9918 7821 10050 7826
rect 9814 7687 9815 7713
rect 9841 7687 9842 7713
rect 9814 7681 9842 7687
rect 9422 7658 9450 7663
rect 9422 7611 9450 7630
rect 10430 7574 10458 8807
rect 10710 8834 10738 8839
rect 10766 8834 10794 9198
rect 10934 9225 10962 9231
rect 10934 9199 10935 9225
rect 10961 9199 10962 9225
rect 10934 9170 10962 9199
rect 10934 9137 10962 9142
rect 10710 8833 10794 8834
rect 10710 8807 10711 8833
rect 10737 8807 10794 8833
rect 10710 8806 10794 8807
rect 10710 8801 10738 8806
rect 10822 8722 10850 8727
rect 10822 8721 10962 8722
rect 10822 8695 10823 8721
rect 10849 8695 10962 8721
rect 10822 8694 10962 8695
rect 10822 8689 10850 8694
rect 10822 8610 10850 8615
rect 10822 8049 10850 8582
rect 10934 8498 10962 8694
rect 10934 8451 10962 8470
rect 11046 8553 11074 8559
rect 11046 8527 11047 8553
rect 11073 8527 11074 8553
rect 11046 8330 11074 8527
rect 11102 8442 11130 8447
rect 11102 8395 11130 8414
rect 11158 8441 11186 9534
rect 11214 9281 11242 10822
rect 11382 10794 11410 11942
rect 11606 11186 11634 12335
rect 11830 12361 11858 12367
rect 11830 12335 11831 12361
rect 11857 12335 11858 12361
rect 11830 12194 11858 12335
rect 11942 12362 11970 12367
rect 11942 12315 11970 12334
rect 12166 12362 12194 12367
rect 12166 12315 12194 12334
rect 13006 12362 13034 12367
rect 11830 12161 11858 12166
rect 11886 12305 11914 12311
rect 11886 12279 11887 12305
rect 11913 12279 11914 12305
rect 11886 12082 11914 12279
rect 11718 12054 11914 12082
rect 13006 12081 13034 12334
rect 18830 12361 18858 12367
rect 18830 12335 18831 12361
rect 18857 12335 18858 12361
rect 17598 12166 17730 12171
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17598 12133 17730 12138
rect 13006 12055 13007 12081
rect 13033 12055 13034 12081
rect 11718 12025 11746 12054
rect 13006 12049 13034 12055
rect 11718 11999 11719 12025
rect 11745 11999 11746 12025
rect 11718 11993 11746 11999
rect 12782 12026 12810 12031
rect 12782 11979 12810 11998
rect 18830 12026 18858 12335
rect 20006 12249 20034 12255
rect 20006 12223 20007 12249
rect 20033 12223 20034 12249
rect 20006 12138 20034 12223
rect 20006 12105 20034 12110
rect 18830 11993 18858 11998
rect 13006 11970 13034 11975
rect 13006 11913 13034 11942
rect 13006 11887 13007 11913
rect 13033 11887 13034 11913
rect 13006 11881 13034 11887
rect 13062 11913 13090 11919
rect 13062 11887 13063 11913
rect 13089 11887 13090 11913
rect 13062 11634 13090 11887
rect 13062 11601 13090 11606
rect 13454 11633 13482 11639
rect 13454 11607 13455 11633
rect 13481 11607 13482 11633
rect 13342 11578 13370 11583
rect 13230 11577 13370 11578
rect 13230 11551 13343 11577
rect 13369 11551 13370 11577
rect 13230 11550 13370 11551
rect 11662 11298 11690 11303
rect 11662 11251 11690 11270
rect 13230 11241 13258 11550
rect 13342 11545 13370 11550
rect 13230 11215 13231 11241
rect 13257 11215 13258 11241
rect 13230 11209 13258 11215
rect 11662 11186 11690 11191
rect 11606 11185 11690 11186
rect 11606 11159 11663 11185
rect 11689 11159 11690 11185
rect 11606 11158 11690 11159
rect 11550 11074 11578 11079
rect 11382 10761 11410 10766
rect 11438 11073 11578 11074
rect 11438 11047 11551 11073
rect 11577 11047 11578 11073
rect 11438 11046 11578 11047
rect 11270 10737 11298 10743
rect 11270 10711 11271 10737
rect 11297 10711 11298 10737
rect 11270 9505 11298 10711
rect 11326 10402 11354 10407
rect 11326 10401 11410 10402
rect 11326 10375 11327 10401
rect 11353 10375 11410 10401
rect 11326 10374 11410 10375
rect 11326 10369 11354 10374
rect 11326 10289 11354 10295
rect 11326 10263 11327 10289
rect 11353 10263 11354 10289
rect 11326 9954 11354 10263
rect 11326 9921 11354 9926
rect 11382 10290 11410 10374
rect 11326 9618 11354 9623
rect 11382 9618 11410 10262
rect 11326 9617 11410 9618
rect 11326 9591 11327 9617
rect 11353 9591 11410 9617
rect 11326 9590 11410 9591
rect 11438 9617 11466 11046
rect 11550 11041 11578 11046
rect 11662 10906 11690 11158
rect 12838 11185 12866 11191
rect 12838 11159 12839 11185
rect 12865 11159 12866 11185
rect 11830 11129 11858 11135
rect 11830 11103 11831 11129
rect 11857 11103 11858 11129
rect 11690 10878 11802 10906
rect 11662 10859 11690 10878
rect 11662 10402 11690 10407
rect 11662 10065 11690 10374
rect 11662 10039 11663 10065
rect 11689 10039 11690 10065
rect 11662 10033 11690 10039
rect 11438 9591 11439 9617
rect 11465 9591 11466 9617
rect 11326 9585 11354 9590
rect 11438 9585 11466 9591
rect 11774 9618 11802 10878
rect 11830 10738 11858 11103
rect 11942 11130 11970 11135
rect 11942 11129 12026 11130
rect 11942 11103 11943 11129
rect 11969 11103 12026 11129
rect 11942 11102 12026 11103
rect 11942 11097 11970 11102
rect 11830 10705 11858 10710
rect 11942 9618 11970 9623
rect 11774 9617 11970 9618
rect 11774 9591 11943 9617
rect 11969 9591 11970 9617
rect 11774 9590 11970 9591
rect 11942 9585 11970 9590
rect 11998 9618 12026 11102
rect 12838 10794 12866 11159
rect 13454 10850 13482 11607
rect 13790 11633 13818 11639
rect 13790 11607 13791 11633
rect 13817 11607 13818 11633
rect 13510 11578 13538 11583
rect 13678 11578 13706 11583
rect 13510 11577 13706 11578
rect 13510 11551 13511 11577
rect 13537 11551 13679 11577
rect 13705 11551 13706 11577
rect 13510 11550 13706 11551
rect 13510 11545 13538 11550
rect 13678 11545 13706 11550
rect 13790 11578 13818 11607
rect 13790 11545 13818 11550
rect 13846 11634 13874 11639
rect 13846 11577 13874 11606
rect 13846 11551 13847 11577
rect 13873 11551 13874 11577
rect 13846 11186 13874 11551
rect 14294 11578 14322 11583
rect 14294 11241 14322 11550
rect 18830 11578 18858 11583
rect 18830 11531 18858 11550
rect 20006 11466 20034 11471
rect 20006 11419 20034 11438
rect 17598 11382 17730 11387
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17598 11349 17730 11354
rect 14294 11215 14295 11241
rect 14321 11215 14322 11241
rect 14294 11209 14322 11215
rect 20006 11241 20034 11247
rect 20006 11215 20007 11241
rect 20033 11215 20034 11241
rect 13790 11158 13874 11186
rect 18830 11185 18858 11191
rect 18830 11159 18831 11185
rect 18857 11159 18858 11185
rect 13454 10822 13594 10850
rect 12838 10761 12866 10766
rect 13174 10794 13202 10799
rect 12334 10738 12362 10743
rect 12334 10402 12362 10710
rect 12334 10369 12362 10374
rect 13174 10345 13202 10766
rect 13510 10738 13538 10743
rect 13174 10319 13175 10345
rect 13201 10319 13202 10345
rect 12782 10066 12810 10071
rect 12782 10019 12810 10038
rect 12670 10009 12698 10015
rect 12670 9983 12671 10009
rect 12697 9983 12698 10009
rect 12054 9730 12082 9735
rect 12054 9683 12082 9702
rect 12278 9674 12306 9679
rect 12502 9674 12530 9679
rect 12278 9673 12530 9674
rect 12278 9647 12279 9673
rect 12305 9647 12503 9673
rect 12529 9647 12530 9673
rect 12278 9646 12530 9647
rect 12278 9641 12306 9646
rect 12502 9641 12530 9646
rect 11998 9585 12026 9590
rect 12222 9562 12250 9567
rect 12222 9515 12250 9534
rect 12334 9561 12362 9567
rect 12334 9535 12335 9561
rect 12361 9535 12362 9561
rect 11270 9479 11271 9505
rect 11297 9479 11298 9505
rect 11270 9473 11298 9479
rect 12334 9506 12362 9535
rect 12334 9473 12362 9478
rect 12558 9505 12586 9511
rect 12558 9479 12559 9505
rect 12585 9479 12586 9505
rect 11662 9338 11690 9343
rect 11214 9255 11215 9281
rect 11241 9255 11242 9281
rect 11214 9249 11242 9255
rect 11550 9310 11662 9338
rect 11382 8497 11410 8503
rect 11382 8471 11383 8497
rect 11409 8471 11410 8497
rect 11382 8442 11410 8471
rect 11158 8415 11159 8441
rect 11185 8415 11186 8441
rect 11158 8409 11186 8415
rect 11214 8414 11410 8442
rect 11550 8441 11578 9310
rect 11662 9291 11690 9310
rect 12558 9170 12586 9479
rect 12614 9505 12642 9511
rect 12614 9479 12615 9505
rect 12641 9479 12642 9505
rect 12614 9338 12642 9479
rect 12670 9506 12698 9983
rect 12670 9473 12698 9478
rect 12894 9562 12922 9567
rect 12614 9305 12642 9310
rect 12894 9394 12922 9534
rect 13062 9506 13090 9511
rect 13062 9459 13090 9478
rect 12894 9337 12922 9366
rect 12894 9311 12895 9337
rect 12921 9311 12922 9337
rect 12894 9305 12922 9311
rect 12222 9142 12586 9170
rect 13062 9281 13090 9287
rect 13062 9255 13063 9281
rect 13089 9255 13090 9281
rect 12222 8889 12250 9142
rect 13062 9114 13090 9255
rect 13174 9226 13202 10319
rect 13286 10737 13538 10738
rect 13286 10711 13511 10737
rect 13537 10711 13538 10737
rect 13286 10710 13538 10711
rect 13286 10065 13314 10710
rect 13510 10705 13538 10710
rect 13566 10094 13594 10822
rect 13286 10039 13287 10065
rect 13313 10039 13314 10065
rect 13286 10033 13314 10039
rect 13510 10066 13594 10094
rect 13790 10066 13818 11158
rect 18830 10906 18858 11159
rect 20006 11130 20034 11215
rect 20006 11097 20034 11102
rect 18830 10873 18858 10878
rect 14910 10850 14938 10855
rect 14910 10803 14938 10822
rect 14798 10794 14826 10799
rect 14574 10766 14798 10794
rect 13230 10010 13258 10015
rect 13230 9963 13258 9982
rect 13342 10009 13370 10015
rect 13342 9983 13343 10009
rect 13369 9983 13370 10009
rect 13342 9954 13370 9983
rect 13342 9921 13370 9926
rect 13510 9954 13538 10066
rect 13790 10019 13818 10038
rect 13846 10738 13874 10743
rect 13846 10065 13874 10710
rect 14574 10738 14602 10766
rect 14798 10747 14826 10766
rect 18830 10794 18858 10799
rect 18830 10747 18858 10766
rect 20006 10794 20034 10799
rect 14574 10691 14602 10710
rect 20006 10737 20034 10766
rect 20006 10711 20007 10737
rect 20033 10711 20034 10737
rect 20006 10705 20034 10711
rect 17598 10598 17730 10603
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17598 10565 17730 10570
rect 20006 10458 20034 10463
rect 20006 10411 20034 10430
rect 18830 10402 18858 10407
rect 18830 10355 18858 10374
rect 13846 10039 13847 10065
rect 13873 10039 13874 10065
rect 13846 10033 13874 10039
rect 13902 10066 13930 10071
rect 13510 9921 13538 9926
rect 13566 10009 13594 10015
rect 13566 9983 13567 10009
rect 13593 9983 13594 10009
rect 13566 9898 13594 9983
rect 13846 9898 13874 9903
rect 13566 9897 13874 9898
rect 13566 9871 13847 9897
rect 13873 9871 13874 9897
rect 13566 9870 13874 9871
rect 13846 9865 13874 9870
rect 13678 9618 13706 9623
rect 13678 9571 13706 9590
rect 13846 9618 13874 9623
rect 13902 9618 13930 10038
rect 20006 10066 20034 10071
rect 18942 10009 18970 10015
rect 18942 9983 18943 10009
rect 18969 9983 18970 10009
rect 17598 9814 17730 9819
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17598 9781 17730 9786
rect 13846 9617 13930 9618
rect 13846 9591 13847 9617
rect 13873 9591 13930 9617
rect 13846 9590 13930 9591
rect 14574 9618 14602 9623
rect 13846 9585 13874 9590
rect 13510 9561 13538 9567
rect 13510 9535 13511 9561
rect 13537 9535 13538 9561
rect 13286 9394 13314 9399
rect 13230 9226 13258 9231
rect 13174 9225 13258 9226
rect 13174 9199 13231 9225
rect 13257 9199 13258 9225
rect 13174 9198 13258 9199
rect 13062 9081 13090 9086
rect 12222 8863 12223 8889
rect 12249 8863 12250 8889
rect 12222 8857 12250 8863
rect 11830 8833 11858 8839
rect 11830 8807 11831 8833
rect 11857 8807 11858 8833
rect 11830 8610 11858 8807
rect 11830 8577 11858 8582
rect 13230 8610 13258 9198
rect 13286 8889 13314 9366
rect 13510 9338 13538 9535
rect 13510 9305 13538 9310
rect 13734 9505 13762 9511
rect 13734 9479 13735 9505
rect 13761 9479 13762 9505
rect 13734 9282 13762 9479
rect 13734 9254 14154 9282
rect 13622 9170 13650 9175
rect 13622 9169 14098 9170
rect 13622 9143 13623 9169
rect 13649 9143 14098 9169
rect 13622 9142 14098 9143
rect 13622 9137 13650 9142
rect 14070 8945 14098 9142
rect 14070 8919 14071 8945
rect 14097 8919 14098 8945
rect 14070 8913 14098 8919
rect 13286 8863 13287 8889
rect 13313 8863 13314 8889
rect 13286 8857 13314 8863
rect 14126 8889 14154 9254
rect 14126 8863 14127 8889
rect 14153 8863 14154 8889
rect 14126 8857 14154 8863
rect 14574 8833 14602 9590
rect 14854 9618 14882 9623
rect 14742 9506 14770 9511
rect 14742 9459 14770 9478
rect 14854 9337 14882 9590
rect 18830 9617 18858 9623
rect 18830 9591 18831 9617
rect 18857 9591 18858 9617
rect 14854 9311 14855 9337
rect 14881 9311 14882 9337
rect 14854 9226 14882 9311
rect 18774 9506 18802 9511
rect 15358 9281 15386 9287
rect 15358 9255 15359 9281
rect 15385 9255 15386 9281
rect 14854 9193 14882 9198
rect 15022 9225 15050 9231
rect 15022 9199 15023 9225
rect 15049 9199 15050 9225
rect 14686 9170 14714 9175
rect 14686 9123 14714 9142
rect 15022 9170 15050 9199
rect 15190 9226 15218 9231
rect 15190 9179 15218 9198
rect 15022 9137 15050 9142
rect 14574 8807 14575 8833
rect 14601 8807 14602 8833
rect 14574 8801 14602 8807
rect 14742 8722 14770 8727
rect 14742 8675 14770 8694
rect 13230 8577 13258 8582
rect 11550 8415 11551 8441
rect 11577 8415 11578 8441
rect 11214 8330 11242 8414
rect 11550 8409 11578 8415
rect 11718 8442 11746 8447
rect 12222 8442 12250 8447
rect 11746 8414 11802 8442
rect 11718 8409 11746 8414
rect 11438 8386 11466 8391
rect 11046 8302 11242 8330
rect 11270 8385 11466 8386
rect 11270 8359 11439 8385
rect 11465 8359 11466 8385
rect 11270 8358 11466 8359
rect 11270 8162 11298 8358
rect 11438 8353 11466 8358
rect 11158 8134 11298 8162
rect 11158 8105 11186 8134
rect 11158 8079 11159 8105
rect 11185 8079 11186 8105
rect 11158 8073 11186 8079
rect 10822 8023 10823 8049
rect 10849 8023 10850 8049
rect 10822 8017 10850 8023
rect 11774 7657 11802 8414
rect 12222 8105 12250 8414
rect 12222 8079 12223 8105
rect 12249 8079 12250 8105
rect 11774 7631 11775 7657
rect 11801 7631 11802 7657
rect 11774 7625 11802 7631
rect 11886 7713 11914 7719
rect 11886 7687 11887 7713
rect 11913 7687 11914 7713
rect 10878 7601 10906 7607
rect 10878 7575 10879 7601
rect 10905 7575 10906 7601
rect 10878 7574 10906 7575
rect 10430 7546 10906 7574
rect 9918 7070 10050 7075
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 9918 7037 10050 7042
rect 9918 6286 10050 6291
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 9918 6253 10050 6258
rect 9918 5502 10050 5507
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 9918 5469 10050 5474
rect 9918 4718 10050 4723
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 9918 4685 10050 4690
rect 10878 4214 10906 7546
rect 10542 4186 10906 4214
rect 9918 3934 10050 3939
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 9918 3901 10050 3906
rect 9918 3150 10050 3155
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 9918 3117 10050 3122
rect 9918 2366 10050 2371
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 9918 2333 10050 2338
rect 9310 1834 9338 1839
rect 8806 1751 8807 1777
rect 8833 1751 8834 1777
rect 8806 1745 8834 1751
rect 9086 1833 9338 1834
rect 9086 1807 9311 1833
rect 9337 1807 9338 1833
rect 9086 1806 9338 1807
rect 9086 400 9114 1806
rect 9310 1801 9338 1806
rect 10430 1834 10458 1839
rect 9918 1582 10050 1587
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 9918 1549 10050 1554
rect 10430 400 10458 1806
rect 10542 1777 10570 4186
rect 11774 2618 11802 2623
rect 11046 1834 11074 1839
rect 11046 1787 11074 1806
rect 11438 1834 11466 1839
rect 10542 1751 10543 1777
rect 10569 1751 10570 1777
rect 10542 1745 10570 1751
rect 11438 400 11466 1806
rect 11774 400 11802 2590
rect 11886 2561 11914 7687
rect 12222 7574 12250 8079
rect 15358 8050 15386 9255
rect 18718 9170 18746 9175
rect 17598 9030 17730 9035
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17598 8997 17730 9002
rect 17598 8246 17730 8251
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17598 8213 17730 8218
rect 15358 8017 15386 8022
rect 18718 7658 18746 9142
rect 18774 8834 18802 9478
rect 18830 9450 18858 9591
rect 18830 9417 18858 9422
rect 18942 9394 18970 9983
rect 20006 9953 20034 10038
rect 20006 9927 20007 9953
rect 20033 9927 20034 9953
rect 20006 9921 20034 9927
rect 20006 9786 20034 9791
rect 20006 9729 20034 9758
rect 20006 9703 20007 9729
rect 20033 9703 20034 9729
rect 20006 9697 20034 9703
rect 18942 9361 18970 9366
rect 20006 9450 20034 9455
rect 18830 9226 18858 9231
rect 18830 9179 18858 9198
rect 20006 9169 20034 9422
rect 20006 9143 20007 9169
rect 20033 9143 20034 9169
rect 20006 9137 20034 9143
rect 19950 9114 19978 9119
rect 19950 8889 19978 9086
rect 19950 8863 19951 8889
rect 19977 8863 19978 8889
rect 19950 8857 19978 8863
rect 18830 8834 18858 8839
rect 18774 8833 18858 8834
rect 18774 8807 18831 8833
rect 18857 8807 18858 8833
rect 18774 8806 18858 8807
rect 18830 8801 18858 8806
rect 19670 8778 19698 8783
rect 18830 8722 18858 8727
rect 18830 8441 18858 8694
rect 19670 8497 19698 8750
rect 19670 8471 19671 8497
rect 19697 8471 19698 8497
rect 19670 8465 19698 8471
rect 18830 8415 18831 8441
rect 18857 8415 18858 8441
rect 18830 8409 18858 8415
rect 19894 8386 19922 8391
rect 19894 8105 19922 8358
rect 19894 8079 19895 8105
rect 19921 8079 19922 8105
rect 19894 8073 19922 8079
rect 20006 8106 20034 8111
rect 18830 8050 18858 8055
rect 18830 8003 18858 8022
rect 18830 7658 18858 7663
rect 18718 7657 18858 7658
rect 18718 7631 18831 7657
rect 18857 7631 18858 7657
rect 18718 7630 18858 7631
rect 18830 7625 18858 7630
rect 20006 7601 20034 8078
rect 20006 7575 20007 7601
rect 20033 7575 20034 7601
rect 12222 7546 12306 7574
rect 20006 7569 20034 7575
rect 11886 2535 11887 2561
rect 11913 2535 11914 2561
rect 11886 2529 11914 2535
rect 12278 1777 12306 7546
rect 17598 7462 17730 7467
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17598 7429 17730 7434
rect 17598 6678 17730 6683
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17598 6645 17730 6650
rect 17598 5894 17730 5899
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17598 5861 17730 5866
rect 17598 5110 17730 5115
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17598 5077 17730 5082
rect 17598 4326 17730 4331
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17598 4293 17730 4298
rect 17598 3542 17730 3547
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17598 3509 17730 3514
rect 17598 2758 17730 2763
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17598 2725 17730 2730
rect 12390 2618 12418 2623
rect 12390 2571 12418 2590
rect 17598 1974 17730 1979
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17598 1941 17730 1946
rect 12782 1834 12810 1839
rect 12782 1787 12810 1806
rect 12278 1751 12279 1777
rect 12305 1751 12306 1777
rect 12278 1745 12306 1751
rect 9072 0 9128 400
rect 10416 0 10472 400
rect 11424 0 11480 400
rect 11760 0 11816 400
<< via2 >>
rect 2238 19221 2266 19222
rect 2238 19195 2239 19221
rect 2239 19195 2265 19221
rect 2265 19195 2266 19221
rect 2238 19194 2266 19195
rect 2290 19221 2318 19222
rect 2290 19195 2291 19221
rect 2291 19195 2317 19221
rect 2317 19195 2318 19221
rect 2290 19194 2318 19195
rect 2342 19221 2370 19222
rect 2342 19195 2343 19221
rect 2343 19195 2369 19221
rect 2369 19195 2370 19221
rect 2342 19194 2370 19195
rect 11774 19110 11802 19138
rect 9918 18829 9946 18830
rect 9918 18803 9919 18829
rect 9919 18803 9945 18829
rect 9945 18803 9946 18829
rect 9918 18802 9946 18803
rect 9970 18829 9998 18830
rect 9970 18803 9971 18829
rect 9971 18803 9997 18829
rect 9997 18803 9998 18829
rect 9970 18802 9998 18803
rect 10022 18829 10050 18830
rect 10022 18803 10023 18829
rect 10023 18803 10049 18829
rect 10049 18803 10050 18829
rect 10022 18802 10050 18803
rect 12110 18718 12138 18746
rect 2238 18437 2266 18438
rect 2238 18411 2239 18437
rect 2239 18411 2265 18437
rect 2265 18411 2266 18437
rect 2238 18410 2266 18411
rect 2290 18437 2318 18438
rect 2290 18411 2291 18437
rect 2291 18411 2317 18437
rect 2317 18411 2318 18437
rect 2290 18410 2318 18411
rect 2342 18437 2370 18438
rect 2342 18411 2343 18437
rect 2343 18411 2369 18437
rect 2369 18411 2370 18437
rect 2342 18410 2370 18411
rect 9918 18045 9946 18046
rect 9918 18019 9919 18045
rect 9919 18019 9945 18045
rect 9945 18019 9946 18045
rect 9918 18018 9946 18019
rect 9970 18045 9998 18046
rect 9970 18019 9971 18045
rect 9971 18019 9997 18045
rect 9997 18019 9998 18045
rect 9970 18018 9998 18019
rect 10022 18045 10050 18046
rect 10022 18019 10023 18045
rect 10023 18019 10049 18045
rect 10049 18019 10050 18045
rect 10022 18018 10050 18019
rect 2238 17653 2266 17654
rect 2238 17627 2239 17653
rect 2239 17627 2265 17653
rect 2265 17627 2266 17653
rect 2238 17626 2266 17627
rect 2290 17653 2318 17654
rect 2290 17627 2291 17653
rect 2291 17627 2317 17653
rect 2317 17627 2318 17653
rect 2290 17626 2318 17627
rect 2342 17653 2370 17654
rect 2342 17627 2343 17653
rect 2343 17627 2369 17653
rect 2369 17627 2370 17653
rect 2342 17626 2370 17627
rect 9918 17261 9946 17262
rect 9918 17235 9919 17261
rect 9919 17235 9945 17261
rect 9945 17235 9946 17261
rect 9918 17234 9946 17235
rect 9970 17261 9998 17262
rect 9970 17235 9971 17261
rect 9971 17235 9997 17261
rect 9997 17235 9998 17261
rect 9970 17234 9998 17235
rect 10022 17261 10050 17262
rect 10022 17235 10023 17261
rect 10023 17235 10049 17261
rect 10049 17235 10050 17261
rect 10022 17234 10050 17235
rect 2238 16869 2266 16870
rect 2238 16843 2239 16869
rect 2239 16843 2265 16869
rect 2265 16843 2266 16869
rect 2238 16842 2266 16843
rect 2290 16869 2318 16870
rect 2290 16843 2291 16869
rect 2291 16843 2317 16869
rect 2317 16843 2318 16869
rect 2290 16842 2318 16843
rect 2342 16869 2370 16870
rect 2342 16843 2343 16869
rect 2343 16843 2369 16869
rect 2369 16843 2370 16869
rect 2342 16842 2370 16843
rect 9918 16477 9946 16478
rect 9918 16451 9919 16477
rect 9919 16451 9945 16477
rect 9945 16451 9946 16477
rect 9918 16450 9946 16451
rect 9970 16477 9998 16478
rect 9970 16451 9971 16477
rect 9971 16451 9997 16477
rect 9997 16451 9998 16477
rect 9970 16450 9998 16451
rect 10022 16477 10050 16478
rect 10022 16451 10023 16477
rect 10023 16451 10049 16477
rect 10049 16451 10050 16477
rect 10022 16450 10050 16451
rect 2238 16085 2266 16086
rect 2238 16059 2239 16085
rect 2239 16059 2265 16085
rect 2265 16059 2266 16085
rect 2238 16058 2266 16059
rect 2290 16085 2318 16086
rect 2290 16059 2291 16085
rect 2291 16059 2317 16085
rect 2317 16059 2318 16085
rect 2290 16058 2318 16059
rect 2342 16085 2370 16086
rect 2342 16059 2343 16085
rect 2343 16059 2369 16085
rect 2369 16059 2370 16085
rect 2342 16058 2370 16059
rect 9918 15693 9946 15694
rect 9918 15667 9919 15693
rect 9919 15667 9945 15693
rect 9945 15667 9946 15693
rect 9918 15666 9946 15667
rect 9970 15693 9998 15694
rect 9970 15667 9971 15693
rect 9971 15667 9997 15693
rect 9997 15667 9998 15693
rect 9970 15666 9998 15667
rect 10022 15693 10050 15694
rect 10022 15667 10023 15693
rect 10023 15667 10049 15693
rect 10049 15667 10050 15693
rect 10022 15666 10050 15667
rect 2238 15301 2266 15302
rect 2238 15275 2239 15301
rect 2239 15275 2265 15301
rect 2265 15275 2266 15301
rect 2238 15274 2266 15275
rect 2290 15301 2318 15302
rect 2290 15275 2291 15301
rect 2291 15275 2317 15301
rect 2317 15275 2318 15301
rect 2290 15274 2318 15275
rect 2342 15301 2370 15302
rect 2342 15275 2343 15301
rect 2343 15275 2369 15301
rect 2369 15275 2370 15301
rect 2342 15274 2370 15275
rect 9918 14909 9946 14910
rect 9918 14883 9919 14909
rect 9919 14883 9945 14909
rect 9945 14883 9946 14909
rect 9918 14882 9946 14883
rect 9970 14909 9998 14910
rect 9970 14883 9971 14909
rect 9971 14883 9997 14909
rect 9997 14883 9998 14909
rect 9970 14882 9998 14883
rect 10022 14909 10050 14910
rect 10022 14883 10023 14909
rect 10023 14883 10049 14909
rect 10049 14883 10050 14909
rect 10022 14882 10050 14883
rect 2238 14517 2266 14518
rect 2238 14491 2239 14517
rect 2239 14491 2265 14517
rect 2265 14491 2266 14517
rect 2238 14490 2266 14491
rect 2290 14517 2318 14518
rect 2290 14491 2291 14517
rect 2291 14491 2317 14517
rect 2317 14491 2318 14517
rect 2290 14490 2318 14491
rect 2342 14517 2370 14518
rect 2342 14491 2343 14517
rect 2343 14491 2369 14517
rect 2369 14491 2370 14517
rect 2342 14490 2370 14491
rect 9918 14125 9946 14126
rect 9918 14099 9919 14125
rect 9919 14099 9945 14125
rect 9945 14099 9946 14125
rect 9918 14098 9946 14099
rect 9970 14125 9998 14126
rect 9970 14099 9971 14125
rect 9971 14099 9997 14125
rect 9997 14099 9998 14125
rect 9970 14098 9998 14099
rect 10022 14125 10050 14126
rect 10022 14099 10023 14125
rect 10023 14099 10049 14125
rect 10049 14099 10050 14125
rect 10022 14098 10050 14099
rect 2238 13733 2266 13734
rect 2238 13707 2239 13733
rect 2239 13707 2265 13733
rect 2265 13707 2266 13733
rect 2238 13706 2266 13707
rect 2290 13733 2318 13734
rect 2290 13707 2291 13733
rect 2291 13707 2317 13733
rect 2317 13707 2318 13733
rect 2290 13706 2318 13707
rect 2342 13733 2370 13734
rect 2342 13707 2343 13733
rect 2343 13707 2369 13733
rect 2369 13707 2370 13733
rect 2342 13706 2370 13707
rect 17598 19221 17626 19222
rect 17598 19195 17599 19221
rect 17599 19195 17625 19221
rect 17625 19195 17626 19221
rect 17598 19194 17626 19195
rect 17650 19221 17678 19222
rect 17650 19195 17651 19221
rect 17651 19195 17677 19221
rect 17677 19195 17678 19221
rect 17650 19194 17678 19195
rect 17702 19221 17730 19222
rect 17702 19195 17703 19221
rect 17703 19195 17729 19221
rect 17729 19195 17730 19221
rect 17702 19194 17730 19195
rect 12782 19137 12810 19138
rect 12782 19111 12783 19137
rect 12783 19111 12809 19137
rect 12809 19111 12810 19137
rect 12782 19110 12810 19111
rect 13118 18745 13146 18746
rect 13118 18719 13119 18745
rect 13119 18719 13145 18745
rect 13145 18719 13146 18745
rect 13118 18718 13146 18719
rect 12558 18326 12586 18354
rect 9918 13341 9946 13342
rect 9918 13315 9919 13341
rect 9919 13315 9945 13341
rect 9945 13315 9946 13341
rect 9918 13314 9946 13315
rect 9970 13341 9998 13342
rect 9970 13315 9971 13341
rect 9971 13315 9997 13341
rect 9997 13315 9998 13341
rect 9970 13314 9998 13315
rect 10022 13341 10050 13342
rect 10022 13315 10023 13341
rect 10023 13315 10049 13341
rect 10049 13315 10050 13341
rect 10022 13314 10050 13315
rect 2238 12949 2266 12950
rect 2238 12923 2239 12949
rect 2239 12923 2265 12949
rect 2265 12923 2266 12949
rect 2238 12922 2266 12923
rect 2290 12949 2318 12950
rect 2290 12923 2291 12949
rect 2291 12923 2317 12949
rect 2317 12923 2318 12949
rect 2290 12922 2318 12923
rect 2342 12949 2370 12950
rect 2342 12923 2343 12949
rect 2343 12923 2369 12949
rect 2369 12923 2370 12949
rect 2342 12922 2370 12923
rect 966 12446 994 12474
rect 2086 12782 2114 12810
rect 966 12249 994 12250
rect 966 12223 967 12249
rect 967 12223 993 12249
rect 993 12223 994 12249
rect 966 12222 994 12223
rect 966 11465 994 11466
rect 966 11439 967 11465
rect 967 11439 993 11465
rect 993 11439 994 11465
rect 966 11438 994 11439
rect 966 10766 994 10794
rect 2142 12753 2170 12754
rect 2142 12727 2143 12753
rect 2143 12727 2169 12753
rect 2169 12727 2170 12753
rect 2142 12726 2170 12727
rect 6734 12726 6762 12754
rect 12222 13257 12250 13258
rect 12222 13231 12223 13257
rect 12223 13231 12249 13257
rect 12249 13231 12250 13257
rect 12222 13230 12250 13231
rect 7462 12726 7490 12754
rect 7518 12446 7546 12474
rect 2142 12361 2170 12362
rect 2142 12335 2143 12361
rect 2143 12335 2169 12361
rect 2169 12335 2170 12361
rect 2142 12334 2170 12335
rect 6230 12334 6258 12362
rect 2238 12165 2266 12166
rect 2238 12139 2239 12165
rect 2239 12139 2265 12165
rect 2265 12139 2266 12165
rect 2238 12138 2266 12139
rect 2290 12165 2318 12166
rect 2290 12139 2291 12165
rect 2291 12139 2317 12165
rect 2317 12139 2318 12165
rect 2290 12138 2318 12139
rect 2342 12165 2370 12166
rect 2342 12139 2343 12165
rect 2343 12139 2369 12165
rect 2369 12139 2370 12165
rect 2342 12138 2370 12139
rect 7238 11774 7266 11802
rect 7182 11689 7210 11690
rect 7182 11663 7183 11689
rect 7183 11663 7209 11689
rect 7209 11663 7210 11689
rect 7182 11662 7210 11663
rect 7350 11662 7378 11690
rect 2142 11577 2170 11578
rect 2142 11551 2143 11577
rect 2143 11551 2169 11577
rect 2169 11551 2170 11577
rect 2142 11550 2170 11551
rect 5670 11550 5698 11578
rect 2238 11381 2266 11382
rect 2238 11355 2239 11381
rect 2239 11355 2265 11381
rect 2265 11355 2266 11381
rect 2238 11354 2266 11355
rect 2290 11381 2318 11382
rect 2290 11355 2291 11381
rect 2291 11355 2317 11381
rect 2317 11355 2318 11381
rect 2290 11354 2318 11355
rect 2342 11381 2370 11382
rect 2342 11355 2343 11381
rect 2343 11355 2369 11381
rect 2369 11355 2370 11381
rect 2342 11354 2370 11355
rect 2142 11185 2170 11186
rect 2142 11159 2143 11185
rect 2143 11159 2169 11185
rect 2169 11159 2170 11185
rect 2142 11158 2170 11159
rect 7294 11577 7322 11578
rect 7294 11551 7295 11577
rect 7295 11551 7321 11577
rect 7321 11551 7322 11577
rect 7294 11550 7322 11551
rect 6734 11158 6762 11186
rect 6790 10710 6818 10738
rect 2238 10597 2266 10598
rect 2238 10571 2239 10597
rect 2239 10571 2265 10597
rect 2265 10571 2266 10597
rect 2238 10570 2266 10571
rect 2290 10597 2318 10598
rect 2290 10571 2291 10597
rect 2291 10571 2317 10597
rect 2317 10571 2318 10597
rect 2290 10570 2318 10571
rect 2342 10597 2370 10598
rect 2342 10571 2343 10597
rect 2343 10571 2369 10597
rect 2369 10571 2370 10597
rect 2342 10570 2370 10571
rect 7014 11185 7042 11186
rect 7014 11159 7015 11185
rect 7015 11159 7041 11185
rect 7041 11159 7042 11185
rect 7014 11158 7042 11159
rect 7406 11606 7434 11634
rect 7518 12278 7546 12306
rect 7686 11998 7714 12026
rect 8078 12473 8106 12474
rect 8078 12447 8079 12473
rect 8079 12447 8105 12473
rect 8105 12447 8106 12473
rect 8078 12446 8106 12447
rect 7966 12417 7994 12418
rect 7966 12391 7967 12417
rect 7967 12391 7993 12417
rect 7993 12391 7994 12417
rect 7966 12390 7994 12391
rect 7910 12305 7938 12306
rect 7910 12279 7911 12305
rect 7911 12279 7937 12305
rect 7937 12279 7938 12305
rect 7910 12278 7938 12279
rect 7854 11969 7882 11970
rect 7854 11943 7855 11969
rect 7855 11943 7881 11969
rect 7881 11943 7882 11969
rect 7854 11942 7882 11943
rect 7686 11662 7714 11690
rect 8358 12473 8386 12474
rect 8358 12447 8359 12473
rect 8359 12447 8385 12473
rect 8385 12447 8386 12473
rect 8358 12446 8386 12447
rect 8638 12446 8666 12474
rect 8190 11998 8218 12026
rect 8470 12361 8498 12362
rect 8470 12335 8471 12361
rect 8471 12335 8497 12361
rect 8497 12335 8498 12361
rect 8470 12334 8498 12335
rect 8302 11774 8330 11802
rect 8414 11998 8442 12026
rect 7966 11662 7994 11690
rect 7798 11633 7826 11634
rect 7798 11607 7799 11633
rect 7799 11607 7825 11633
rect 7825 11607 7826 11633
rect 7798 11606 7826 11607
rect 7406 11185 7434 11186
rect 7406 11159 7407 11185
rect 7407 11159 7433 11185
rect 7433 11159 7434 11185
rect 7406 11158 7434 11159
rect 7462 10766 7490 10794
rect 7574 10710 7602 10738
rect 7742 10710 7770 10738
rect 2238 9813 2266 9814
rect 2238 9787 2239 9813
rect 2239 9787 2265 9813
rect 2265 9787 2266 9813
rect 2238 9786 2266 9787
rect 2290 9813 2318 9814
rect 2290 9787 2291 9813
rect 2291 9787 2317 9813
rect 2317 9787 2318 9813
rect 2290 9786 2318 9787
rect 2342 9813 2370 9814
rect 2342 9787 2343 9813
rect 2343 9787 2369 9813
rect 2369 9787 2370 9813
rect 2342 9786 2370 9787
rect 2086 9478 2114 9506
rect 2142 9142 2170 9170
rect 5782 9169 5810 9170
rect 5782 9143 5783 9169
rect 5783 9143 5809 9169
rect 5809 9143 5810 9169
rect 5782 9142 5810 9143
rect 966 9113 994 9114
rect 966 9087 967 9113
rect 967 9087 993 9113
rect 993 9087 994 9113
rect 966 9086 994 9087
rect 2238 9029 2266 9030
rect 2238 9003 2239 9029
rect 2239 9003 2265 9029
rect 2265 9003 2266 9029
rect 2238 9002 2266 9003
rect 2290 9029 2318 9030
rect 2290 9003 2291 9029
rect 2291 9003 2317 9029
rect 2317 9003 2318 9029
rect 2290 9002 2318 9003
rect 2342 9029 2370 9030
rect 2342 9003 2343 9029
rect 2343 9003 2369 9029
rect 2369 9003 2370 9029
rect 2342 9002 2370 9003
rect 2142 8833 2170 8834
rect 2142 8807 2143 8833
rect 2143 8807 2169 8833
rect 2169 8807 2170 8833
rect 2142 8806 2170 8807
rect 6846 9169 6874 9170
rect 6846 9143 6847 9169
rect 6847 9143 6873 9169
rect 6873 9143 6874 9169
rect 6846 9142 6874 9143
rect 7014 9982 7042 10010
rect 8134 10793 8162 10794
rect 8134 10767 8135 10793
rect 8135 10767 8161 10793
rect 8161 10767 8162 10793
rect 8134 10766 8162 10767
rect 8246 10766 8274 10794
rect 8134 10345 8162 10346
rect 8134 10319 8135 10345
rect 8135 10319 8161 10345
rect 8161 10319 8162 10345
rect 8134 10318 8162 10319
rect 8694 11998 8722 12026
rect 8414 10318 8442 10346
rect 8750 11774 8778 11802
rect 8862 11550 8890 11578
rect 8134 10009 8162 10010
rect 8134 9983 8135 10009
rect 8135 9983 8161 10009
rect 8161 9983 8162 10009
rect 8134 9982 8162 9983
rect 7966 9926 7994 9954
rect 6902 9086 6930 9114
rect 5782 8750 5810 8778
rect 6006 8806 6034 8834
rect 966 8414 994 8442
rect 6958 9310 6986 9338
rect 6006 8526 6034 8554
rect 7070 8721 7098 8722
rect 7070 8695 7071 8721
rect 7071 8695 7097 8721
rect 7097 8695 7098 8721
rect 7070 8694 7098 8695
rect 2238 8245 2266 8246
rect 2238 8219 2239 8245
rect 2239 8219 2265 8245
rect 2265 8219 2266 8245
rect 2238 8218 2266 8219
rect 2290 8245 2318 8246
rect 2290 8219 2291 8245
rect 2291 8219 2317 8245
rect 2317 8219 2318 8245
rect 2290 8218 2318 8219
rect 2342 8245 2370 8246
rect 2342 8219 2343 8245
rect 2343 8219 2369 8245
rect 2369 8219 2370 8245
rect 2342 8218 2370 8219
rect 6902 8049 6930 8050
rect 6902 8023 6903 8049
rect 6903 8023 6929 8049
rect 6929 8023 6930 8049
rect 6902 8022 6930 8023
rect 7574 9337 7602 9338
rect 7574 9311 7575 9337
rect 7575 9311 7601 9337
rect 7601 9311 7602 9337
rect 7574 9310 7602 9311
rect 7686 9281 7714 9282
rect 7686 9255 7687 9281
rect 7687 9255 7713 9281
rect 7713 9255 7714 9281
rect 7686 9254 7714 9255
rect 7406 9198 7434 9226
rect 7798 9225 7826 9226
rect 7798 9199 7799 9225
rect 7799 9199 7825 9225
rect 7825 9199 7826 9225
rect 7798 9198 7826 9199
rect 7630 9169 7658 9170
rect 7630 9143 7631 9169
rect 7631 9143 7657 9169
rect 7657 9143 7658 9169
rect 7630 9142 7658 9143
rect 9918 12557 9946 12558
rect 9918 12531 9919 12557
rect 9919 12531 9945 12557
rect 9945 12531 9946 12557
rect 9918 12530 9946 12531
rect 9970 12557 9998 12558
rect 9970 12531 9971 12557
rect 9971 12531 9997 12557
rect 9997 12531 9998 12557
rect 9970 12530 9998 12531
rect 10022 12557 10050 12558
rect 10022 12531 10023 12557
rect 10023 12531 10049 12557
rect 10049 12531 10050 12557
rect 10022 12530 10050 12531
rect 8974 12334 9002 12362
rect 9758 12334 9786 12362
rect 9702 12054 9730 12082
rect 9310 11969 9338 11970
rect 9310 11943 9311 11969
rect 9311 11943 9337 11969
rect 9337 11943 9338 11969
rect 9310 11942 9338 11943
rect 9198 11913 9226 11914
rect 9198 11887 9199 11913
rect 9199 11887 9225 11913
rect 9225 11887 9226 11913
rect 9198 11886 9226 11887
rect 9366 11689 9394 11690
rect 9366 11663 9367 11689
rect 9367 11663 9393 11689
rect 9393 11663 9394 11689
rect 9366 11662 9394 11663
rect 10150 12054 10178 12082
rect 9758 11913 9786 11914
rect 9758 11887 9759 11913
rect 9759 11887 9785 11913
rect 9785 11887 9786 11913
rect 9758 11886 9786 11887
rect 9310 11577 9338 11578
rect 9310 11551 9311 11577
rect 9311 11551 9337 11577
rect 9337 11551 9338 11577
rect 9310 11550 9338 11551
rect 10542 12166 10570 12194
rect 10542 11942 10570 11970
rect 9918 11773 9946 11774
rect 9918 11747 9919 11773
rect 9919 11747 9945 11773
rect 9945 11747 9946 11773
rect 9918 11746 9946 11747
rect 9970 11773 9998 11774
rect 9970 11747 9971 11773
rect 9971 11747 9997 11773
rect 9997 11747 9998 11773
rect 9970 11746 9998 11747
rect 10022 11773 10050 11774
rect 10022 11747 10023 11773
rect 10023 11747 10049 11773
rect 10049 11747 10050 11773
rect 10022 11746 10050 11747
rect 9926 11689 9954 11690
rect 9926 11663 9927 11689
rect 9927 11663 9953 11689
rect 9953 11663 9954 11689
rect 9926 11662 9954 11663
rect 8974 10793 9002 10794
rect 8974 10767 8975 10793
rect 8975 10767 9001 10793
rect 9001 10767 9002 10793
rect 8974 10766 9002 10767
rect 8750 9870 8778 9898
rect 8414 9673 8442 9674
rect 8414 9647 8415 9673
rect 8415 9647 8441 9673
rect 8441 9647 8442 9673
rect 8414 9646 8442 9647
rect 7966 9281 7994 9282
rect 7966 9255 7967 9281
rect 7967 9255 7993 9281
rect 7993 9255 7994 9281
rect 7966 9254 7994 9255
rect 9646 11185 9674 11186
rect 9646 11159 9647 11185
rect 9647 11159 9673 11185
rect 9673 11159 9674 11185
rect 9646 11158 9674 11159
rect 9422 10710 9450 10738
rect 9918 10989 9946 10990
rect 9918 10963 9919 10989
rect 9919 10963 9945 10989
rect 9945 10963 9946 10989
rect 9918 10962 9946 10963
rect 9970 10989 9998 10990
rect 9970 10963 9971 10989
rect 9971 10963 9997 10989
rect 9997 10963 9998 10989
rect 9970 10962 9998 10963
rect 10022 10989 10050 10990
rect 10022 10963 10023 10989
rect 10023 10963 10049 10989
rect 10049 10963 10050 10989
rect 10022 10962 10050 10963
rect 10094 10822 10122 10850
rect 9758 10793 9786 10794
rect 9758 10767 9759 10793
rect 9759 10767 9785 10793
rect 9785 10767 9786 10793
rect 9758 10766 9786 10767
rect 10150 10793 10178 10794
rect 10150 10767 10151 10793
rect 10151 10767 10177 10793
rect 10177 10767 10178 10793
rect 10150 10766 10178 10767
rect 9646 10094 9674 10122
rect 9758 10262 9786 10290
rect 8918 9534 8946 9562
rect 9310 9982 9338 10010
rect 9422 9646 9450 9674
rect 9310 9478 9338 9506
rect 9478 9897 9506 9898
rect 9478 9871 9479 9897
rect 9479 9871 9505 9897
rect 9505 9871 9506 9897
rect 9478 9870 9506 9871
rect 9478 9478 9506 9506
rect 9534 9702 9562 9730
rect 9422 9310 9450 9338
rect 8918 9254 8946 9282
rect 7910 9086 7938 9114
rect 7910 8918 7938 8946
rect 8862 8945 8890 8946
rect 8862 8919 8863 8945
rect 8863 8919 8889 8945
rect 8889 8919 8890 8945
rect 8862 8918 8890 8919
rect 7462 8777 7490 8778
rect 7462 8751 7463 8777
rect 7463 8751 7489 8777
rect 7489 8751 7490 8777
rect 7462 8750 7490 8751
rect 9254 9254 9282 9282
rect 8918 8777 8946 8778
rect 8918 8751 8919 8777
rect 8919 8751 8945 8777
rect 8945 8751 8946 8777
rect 8918 8750 8946 8751
rect 9086 8806 9114 8834
rect 7518 8638 7546 8666
rect 7574 8694 7602 8722
rect 8862 8721 8890 8722
rect 8862 8695 8863 8721
rect 8863 8695 8889 8721
rect 8889 8695 8890 8721
rect 8862 8694 8890 8695
rect 7686 8553 7714 8554
rect 7686 8527 7687 8553
rect 7687 8527 7713 8553
rect 7713 8527 7714 8553
rect 7686 8526 7714 8527
rect 7742 8497 7770 8498
rect 7742 8471 7743 8497
rect 7743 8471 7769 8497
rect 7769 8471 7770 8497
rect 7742 8470 7770 8471
rect 8302 8497 8330 8498
rect 8302 8471 8303 8497
rect 8303 8471 8329 8497
rect 8329 8471 8330 8497
rect 8302 8470 8330 8471
rect 7238 8302 7266 8330
rect 7182 8022 7210 8050
rect 8470 8441 8498 8442
rect 8470 8415 8471 8441
rect 8471 8415 8497 8441
rect 8497 8415 8498 8441
rect 8470 8414 8498 8415
rect 8302 8105 8330 8106
rect 8302 8079 8303 8105
rect 8303 8079 8329 8105
rect 8329 8079 8330 8105
rect 8302 8078 8330 8079
rect 8806 8078 8834 8106
rect 7518 8022 7546 8050
rect 8526 8049 8554 8050
rect 8526 8023 8527 8049
rect 8527 8023 8553 8049
rect 8553 8023 8554 8049
rect 8526 8022 8554 8023
rect 8526 7630 8554 7658
rect 2238 7461 2266 7462
rect 2238 7435 2239 7461
rect 2239 7435 2265 7461
rect 2265 7435 2266 7461
rect 2238 7434 2266 7435
rect 2290 7461 2318 7462
rect 2290 7435 2291 7461
rect 2291 7435 2317 7461
rect 2317 7435 2318 7461
rect 2290 7434 2318 7435
rect 2342 7461 2370 7462
rect 2342 7435 2343 7461
rect 2343 7435 2369 7461
rect 2369 7435 2370 7461
rect 2342 7434 2370 7435
rect 2238 6677 2266 6678
rect 2238 6651 2239 6677
rect 2239 6651 2265 6677
rect 2265 6651 2266 6677
rect 2238 6650 2266 6651
rect 2290 6677 2318 6678
rect 2290 6651 2291 6677
rect 2291 6651 2317 6677
rect 2317 6651 2318 6677
rect 2290 6650 2318 6651
rect 2342 6677 2370 6678
rect 2342 6651 2343 6677
rect 2343 6651 2369 6677
rect 2369 6651 2370 6677
rect 2342 6650 2370 6651
rect 2238 5893 2266 5894
rect 2238 5867 2239 5893
rect 2239 5867 2265 5893
rect 2265 5867 2266 5893
rect 2238 5866 2266 5867
rect 2290 5893 2318 5894
rect 2290 5867 2291 5893
rect 2291 5867 2317 5893
rect 2317 5867 2318 5893
rect 2290 5866 2318 5867
rect 2342 5893 2370 5894
rect 2342 5867 2343 5893
rect 2343 5867 2369 5893
rect 2369 5867 2370 5893
rect 2342 5866 2370 5867
rect 2238 5109 2266 5110
rect 2238 5083 2239 5109
rect 2239 5083 2265 5109
rect 2265 5083 2266 5109
rect 2238 5082 2266 5083
rect 2290 5109 2318 5110
rect 2290 5083 2291 5109
rect 2291 5083 2317 5109
rect 2317 5083 2318 5109
rect 2290 5082 2318 5083
rect 2342 5109 2370 5110
rect 2342 5083 2343 5109
rect 2343 5083 2369 5109
rect 2369 5083 2370 5109
rect 2342 5082 2370 5083
rect 2238 4325 2266 4326
rect 2238 4299 2239 4325
rect 2239 4299 2265 4325
rect 2265 4299 2266 4325
rect 2238 4298 2266 4299
rect 2290 4325 2318 4326
rect 2290 4299 2291 4325
rect 2291 4299 2317 4325
rect 2317 4299 2318 4325
rect 2290 4298 2318 4299
rect 2342 4325 2370 4326
rect 2342 4299 2343 4325
rect 2343 4299 2369 4325
rect 2369 4299 2370 4325
rect 2342 4298 2370 4299
rect 2238 3541 2266 3542
rect 2238 3515 2239 3541
rect 2239 3515 2265 3541
rect 2265 3515 2266 3541
rect 2238 3514 2266 3515
rect 2290 3541 2318 3542
rect 2290 3515 2291 3541
rect 2291 3515 2317 3541
rect 2317 3515 2318 3541
rect 2290 3514 2318 3515
rect 2342 3541 2370 3542
rect 2342 3515 2343 3541
rect 2343 3515 2369 3541
rect 2369 3515 2370 3541
rect 2342 3514 2370 3515
rect 2238 2757 2266 2758
rect 2238 2731 2239 2757
rect 2239 2731 2265 2757
rect 2265 2731 2266 2757
rect 2238 2730 2266 2731
rect 2290 2757 2318 2758
rect 2290 2731 2291 2757
rect 2291 2731 2317 2757
rect 2317 2731 2318 2757
rect 2290 2730 2318 2731
rect 2342 2757 2370 2758
rect 2342 2731 2343 2757
rect 2343 2731 2369 2757
rect 2369 2731 2370 2757
rect 2342 2730 2370 2731
rect 2238 1973 2266 1974
rect 2238 1947 2239 1973
rect 2239 1947 2265 1973
rect 2265 1947 2266 1973
rect 2238 1946 2266 1947
rect 2290 1973 2318 1974
rect 2290 1947 2291 1973
rect 2291 1947 2317 1973
rect 2317 1947 2318 1973
rect 2290 1946 2318 1947
rect 2342 1973 2370 1974
rect 2342 1947 2343 1973
rect 2343 1947 2369 1973
rect 2369 1947 2370 1973
rect 2342 1946 2370 1947
rect 9198 8750 9226 8778
rect 8918 8441 8946 8442
rect 8918 8415 8919 8441
rect 8919 8415 8945 8441
rect 8945 8415 8946 8441
rect 8918 8414 8946 8415
rect 9702 10009 9730 10010
rect 9702 9983 9703 10009
rect 9703 9983 9729 10009
rect 9729 9983 9730 10009
rect 9702 9982 9730 9983
rect 9646 9310 9674 9338
rect 9702 9590 9730 9618
rect 9590 9254 9618 9282
rect 9534 9225 9562 9226
rect 9534 9199 9535 9225
rect 9535 9199 9561 9225
rect 9561 9199 9562 9225
rect 9534 9198 9562 9199
rect 10038 10401 10066 10402
rect 10038 10375 10039 10401
rect 10039 10375 10065 10401
rect 10065 10375 10066 10401
rect 10038 10374 10066 10375
rect 11550 12614 11578 12642
rect 12110 12614 12138 12642
rect 17598 18437 17626 18438
rect 17598 18411 17599 18437
rect 17599 18411 17625 18437
rect 17625 18411 17626 18437
rect 17598 18410 17626 18411
rect 17650 18437 17678 18438
rect 17650 18411 17651 18437
rect 17651 18411 17677 18437
rect 17677 18411 17678 18437
rect 17650 18410 17678 18411
rect 17702 18437 17730 18438
rect 17702 18411 17703 18437
rect 17703 18411 17729 18437
rect 17729 18411 17730 18437
rect 17702 18410 17730 18411
rect 13062 18353 13090 18354
rect 13062 18327 13063 18353
rect 13063 18327 13089 18353
rect 13089 18327 13090 18353
rect 13062 18326 13090 18327
rect 12614 13230 12642 13258
rect 17598 17653 17626 17654
rect 17598 17627 17599 17653
rect 17599 17627 17625 17653
rect 17625 17627 17626 17653
rect 17598 17626 17626 17627
rect 17650 17653 17678 17654
rect 17650 17627 17651 17653
rect 17651 17627 17677 17653
rect 17677 17627 17678 17653
rect 17650 17626 17678 17627
rect 17702 17653 17730 17654
rect 17702 17627 17703 17653
rect 17703 17627 17729 17653
rect 17729 17627 17730 17653
rect 17702 17626 17730 17627
rect 17598 16869 17626 16870
rect 17598 16843 17599 16869
rect 17599 16843 17625 16869
rect 17625 16843 17626 16869
rect 17598 16842 17626 16843
rect 17650 16869 17678 16870
rect 17650 16843 17651 16869
rect 17651 16843 17677 16869
rect 17677 16843 17678 16869
rect 17650 16842 17678 16843
rect 17702 16869 17730 16870
rect 17702 16843 17703 16869
rect 17703 16843 17729 16869
rect 17729 16843 17730 16869
rect 17702 16842 17730 16843
rect 17598 16085 17626 16086
rect 17598 16059 17599 16085
rect 17599 16059 17625 16085
rect 17625 16059 17626 16085
rect 17598 16058 17626 16059
rect 17650 16085 17678 16086
rect 17650 16059 17651 16085
rect 17651 16059 17677 16085
rect 17677 16059 17678 16085
rect 17650 16058 17678 16059
rect 17702 16085 17730 16086
rect 17702 16059 17703 16085
rect 17703 16059 17729 16085
rect 17729 16059 17730 16085
rect 17702 16058 17730 16059
rect 17598 15301 17626 15302
rect 17598 15275 17599 15301
rect 17599 15275 17625 15301
rect 17625 15275 17626 15301
rect 17598 15274 17626 15275
rect 17650 15301 17678 15302
rect 17650 15275 17651 15301
rect 17651 15275 17677 15301
rect 17677 15275 17678 15301
rect 17650 15274 17678 15275
rect 17702 15301 17730 15302
rect 17702 15275 17703 15301
rect 17703 15275 17729 15301
rect 17729 15275 17730 15301
rect 17702 15274 17730 15275
rect 17598 14517 17626 14518
rect 17598 14491 17599 14517
rect 17599 14491 17625 14517
rect 17625 14491 17626 14517
rect 17598 14490 17626 14491
rect 17650 14517 17678 14518
rect 17650 14491 17651 14517
rect 17651 14491 17677 14517
rect 17677 14491 17678 14517
rect 17650 14490 17678 14491
rect 17702 14517 17730 14518
rect 17702 14491 17703 14517
rect 17703 14491 17729 14517
rect 17729 14491 17730 14517
rect 17702 14490 17730 14491
rect 17598 13733 17626 13734
rect 17598 13707 17599 13733
rect 17599 13707 17625 13733
rect 17625 13707 17626 13733
rect 17598 13706 17626 13707
rect 17650 13733 17678 13734
rect 17650 13707 17651 13733
rect 17651 13707 17677 13733
rect 17677 13707 17678 13733
rect 17650 13706 17678 13707
rect 17702 13733 17730 13734
rect 17702 13707 17703 13733
rect 17703 13707 17729 13733
rect 17729 13707 17730 13733
rect 17702 13706 17730 13707
rect 17598 12949 17626 12950
rect 17598 12923 17599 12949
rect 17599 12923 17625 12949
rect 17625 12923 17626 12949
rect 17598 12922 17626 12923
rect 17650 12949 17678 12950
rect 17650 12923 17651 12949
rect 17651 12923 17677 12949
rect 17677 12923 17678 12949
rect 17650 12922 17678 12923
rect 17702 12949 17730 12950
rect 17702 12923 17703 12949
rect 17703 12923 17729 12949
rect 17729 12923 17730 12949
rect 17702 12922 17730 12923
rect 12390 12614 12418 12642
rect 12782 12614 12810 12642
rect 11382 12361 11410 12362
rect 11382 12335 11383 12361
rect 11383 12335 11409 12361
rect 11409 12335 11410 12361
rect 11382 12334 11410 12335
rect 10710 11662 10738 11690
rect 10990 11297 11018 11298
rect 10990 11271 10991 11297
rect 10991 11271 11017 11297
rect 11017 11271 11018 11297
rect 10990 11270 11018 11271
rect 10766 11185 10794 11186
rect 10766 11159 10767 11185
rect 10767 11159 10793 11185
rect 10793 11159 10794 11185
rect 10766 11158 10794 11159
rect 10766 10905 10794 10906
rect 10766 10879 10767 10905
rect 10767 10879 10793 10905
rect 10793 10879 10794 10905
rect 10766 10878 10794 10879
rect 10822 10822 10850 10850
rect 10934 10793 10962 10794
rect 10934 10767 10935 10793
rect 10935 10767 10961 10793
rect 10961 10767 10962 10793
rect 10934 10766 10962 10767
rect 9918 10205 9946 10206
rect 9918 10179 9919 10205
rect 9919 10179 9945 10205
rect 9945 10179 9946 10205
rect 9918 10178 9946 10179
rect 9970 10205 9998 10206
rect 9970 10179 9971 10205
rect 9971 10179 9997 10205
rect 9997 10179 9998 10205
rect 9970 10178 9998 10179
rect 10022 10205 10050 10206
rect 10022 10179 10023 10205
rect 10023 10179 10049 10205
rect 10049 10179 10050 10205
rect 10022 10178 10050 10179
rect 9814 9702 9842 9730
rect 10038 10094 10066 10122
rect 9366 8777 9394 8778
rect 9366 8751 9367 8777
rect 9367 8751 9393 8777
rect 9393 8751 9394 8777
rect 9366 8750 9394 8751
rect 9478 8721 9506 8722
rect 9478 8695 9479 8721
rect 9479 8695 9505 8721
rect 9505 8695 9506 8721
rect 9478 8694 9506 8695
rect 9758 8806 9786 8834
rect 9926 9505 9954 9506
rect 9926 9479 9927 9505
rect 9927 9479 9953 9505
rect 9953 9479 9954 9505
rect 9926 9478 9954 9479
rect 10374 10262 10402 10290
rect 10094 9982 10122 10010
rect 10094 9617 10122 9618
rect 10094 9591 10095 9617
rect 10095 9591 10121 9617
rect 10121 9591 10122 9617
rect 10094 9590 10122 9591
rect 9918 9421 9946 9422
rect 9918 9395 9919 9421
rect 9919 9395 9945 9421
rect 9945 9395 9946 9421
rect 9918 9394 9946 9395
rect 9970 9421 9998 9422
rect 9970 9395 9971 9421
rect 9971 9395 9997 9421
rect 9997 9395 9998 9421
rect 9970 9394 9998 9395
rect 10022 9421 10050 9422
rect 10022 9395 10023 9421
rect 10023 9395 10049 9421
rect 10049 9395 10050 9421
rect 10022 9394 10050 9395
rect 9870 9310 9898 9338
rect 9926 9281 9954 9282
rect 9926 9255 9927 9281
rect 9927 9255 9953 9281
rect 9953 9255 9954 9281
rect 9926 9254 9954 9255
rect 10038 9142 10066 9170
rect 9870 8806 9898 8834
rect 10262 9729 10290 9730
rect 10262 9703 10263 9729
rect 10263 9703 10289 9729
rect 10289 9703 10290 9729
rect 10262 9702 10290 9703
rect 10710 10289 10738 10290
rect 10710 10263 10711 10289
rect 10711 10263 10737 10289
rect 10737 10263 10738 10289
rect 10710 10262 10738 10263
rect 10654 9310 10682 9338
rect 11214 10822 11242 10850
rect 11046 10345 11074 10346
rect 11046 10319 11047 10345
rect 11047 10319 11073 10345
rect 11073 10319 11074 10345
rect 11046 10318 11074 10319
rect 10990 9702 11018 9730
rect 10822 9561 10850 9562
rect 10822 9535 10823 9561
rect 10823 9535 10849 9561
rect 10849 9535 10850 9561
rect 10822 9534 10850 9535
rect 11102 9534 11130 9562
rect 10766 9198 10794 9226
rect 10206 8777 10234 8778
rect 10206 8751 10207 8777
rect 10207 8751 10233 8777
rect 10233 8751 10234 8777
rect 10206 8750 10234 8751
rect 9918 8637 9946 8638
rect 9918 8611 9919 8637
rect 9919 8611 9945 8637
rect 9945 8611 9946 8637
rect 9918 8610 9946 8611
rect 9970 8637 9998 8638
rect 9970 8611 9971 8637
rect 9971 8611 9997 8637
rect 9997 8611 9998 8637
rect 9970 8610 9998 8611
rect 10022 8637 10050 8638
rect 10022 8611 10023 8637
rect 10023 8611 10049 8637
rect 10049 8611 10050 8637
rect 10022 8610 10050 8611
rect 8974 8329 9002 8330
rect 8974 8303 8975 8329
rect 8975 8303 9001 8329
rect 9001 8303 9002 8329
rect 8974 8302 9002 8303
rect 9926 8441 9954 8442
rect 9926 8415 9927 8441
rect 9927 8415 9953 8441
rect 9953 8415 9954 8441
rect 9926 8414 9954 8415
rect 10150 8414 10178 8442
rect 9918 7853 9946 7854
rect 9918 7827 9919 7853
rect 9919 7827 9945 7853
rect 9945 7827 9946 7853
rect 9918 7826 9946 7827
rect 9970 7853 9998 7854
rect 9970 7827 9971 7853
rect 9971 7827 9997 7853
rect 9997 7827 9998 7853
rect 9970 7826 9998 7827
rect 10022 7853 10050 7854
rect 10022 7827 10023 7853
rect 10023 7827 10049 7853
rect 10049 7827 10050 7853
rect 10022 7826 10050 7827
rect 9422 7657 9450 7658
rect 9422 7631 9423 7657
rect 9423 7631 9449 7657
rect 9449 7631 9450 7657
rect 9422 7630 9450 7631
rect 10934 9142 10962 9170
rect 10822 8582 10850 8610
rect 10934 8497 10962 8498
rect 10934 8471 10935 8497
rect 10935 8471 10961 8497
rect 10961 8471 10962 8497
rect 10934 8470 10962 8471
rect 11102 8441 11130 8442
rect 11102 8415 11103 8441
rect 11103 8415 11129 8441
rect 11129 8415 11130 8441
rect 11102 8414 11130 8415
rect 11942 12361 11970 12362
rect 11942 12335 11943 12361
rect 11943 12335 11969 12361
rect 11969 12335 11970 12361
rect 11942 12334 11970 12335
rect 12166 12361 12194 12362
rect 12166 12335 12167 12361
rect 12167 12335 12193 12361
rect 12193 12335 12194 12361
rect 12166 12334 12194 12335
rect 13006 12334 13034 12362
rect 11830 12166 11858 12194
rect 17598 12165 17626 12166
rect 17598 12139 17599 12165
rect 17599 12139 17625 12165
rect 17625 12139 17626 12165
rect 17598 12138 17626 12139
rect 17650 12165 17678 12166
rect 17650 12139 17651 12165
rect 17651 12139 17677 12165
rect 17677 12139 17678 12165
rect 17650 12138 17678 12139
rect 17702 12165 17730 12166
rect 17702 12139 17703 12165
rect 17703 12139 17729 12165
rect 17729 12139 17730 12165
rect 17702 12138 17730 12139
rect 12782 12025 12810 12026
rect 12782 11999 12783 12025
rect 12783 11999 12809 12025
rect 12809 11999 12810 12025
rect 12782 11998 12810 11999
rect 20006 12110 20034 12138
rect 18830 11998 18858 12026
rect 13006 11942 13034 11970
rect 13062 11606 13090 11634
rect 11662 11297 11690 11298
rect 11662 11271 11663 11297
rect 11663 11271 11689 11297
rect 11689 11271 11690 11297
rect 11662 11270 11690 11271
rect 11382 10766 11410 10794
rect 11326 9926 11354 9954
rect 11382 10262 11410 10290
rect 11662 10878 11690 10906
rect 11662 10401 11690 10402
rect 11662 10375 11663 10401
rect 11663 10375 11689 10401
rect 11689 10375 11690 10401
rect 11662 10374 11690 10375
rect 11830 10710 11858 10738
rect 13790 11550 13818 11578
rect 13846 11606 13874 11634
rect 14294 11550 14322 11578
rect 18830 11577 18858 11578
rect 18830 11551 18831 11577
rect 18831 11551 18857 11577
rect 18857 11551 18858 11577
rect 18830 11550 18858 11551
rect 20006 11465 20034 11466
rect 20006 11439 20007 11465
rect 20007 11439 20033 11465
rect 20033 11439 20034 11465
rect 20006 11438 20034 11439
rect 17598 11381 17626 11382
rect 17598 11355 17599 11381
rect 17599 11355 17625 11381
rect 17625 11355 17626 11381
rect 17598 11354 17626 11355
rect 17650 11381 17678 11382
rect 17650 11355 17651 11381
rect 17651 11355 17677 11381
rect 17677 11355 17678 11381
rect 17650 11354 17678 11355
rect 17702 11381 17730 11382
rect 17702 11355 17703 11381
rect 17703 11355 17729 11381
rect 17729 11355 17730 11381
rect 17702 11354 17730 11355
rect 12838 10766 12866 10794
rect 13174 10793 13202 10794
rect 13174 10767 13175 10793
rect 13175 10767 13201 10793
rect 13201 10767 13202 10793
rect 13174 10766 13202 10767
rect 12334 10737 12362 10738
rect 12334 10711 12335 10737
rect 12335 10711 12361 10737
rect 12361 10711 12362 10737
rect 12334 10710 12362 10711
rect 12334 10374 12362 10402
rect 12782 10065 12810 10066
rect 12782 10039 12783 10065
rect 12783 10039 12809 10065
rect 12809 10039 12810 10065
rect 12782 10038 12810 10039
rect 12054 9729 12082 9730
rect 12054 9703 12055 9729
rect 12055 9703 12081 9729
rect 12081 9703 12082 9729
rect 12054 9702 12082 9703
rect 11998 9590 12026 9618
rect 12222 9561 12250 9562
rect 12222 9535 12223 9561
rect 12223 9535 12249 9561
rect 12249 9535 12250 9561
rect 12222 9534 12250 9535
rect 12334 9478 12362 9506
rect 11662 9337 11690 9338
rect 11662 9311 11663 9337
rect 11663 9311 11689 9337
rect 11689 9311 11690 9337
rect 11662 9310 11690 9311
rect 12670 9478 12698 9506
rect 12894 9561 12922 9562
rect 12894 9535 12895 9561
rect 12895 9535 12921 9561
rect 12921 9535 12922 9561
rect 12894 9534 12922 9535
rect 12614 9310 12642 9338
rect 13062 9505 13090 9506
rect 13062 9479 13063 9505
rect 13063 9479 13089 9505
rect 13089 9479 13090 9505
rect 13062 9478 13090 9479
rect 12894 9366 12922 9394
rect 20006 11102 20034 11130
rect 18830 10878 18858 10906
rect 14910 10849 14938 10850
rect 14910 10823 14911 10849
rect 14911 10823 14937 10849
rect 14937 10823 14938 10849
rect 14910 10822 14938 10823
rect 14798 10793 14826 10794
rect 14798 10767 14799 10793
rect 14799 10767 14825 10793
rect 14825 10767 14826 10793
rect 14798 10766 14826 10767
rect 13230 10009 13258 10010
rect 13230 9983 13231 10009
rect 13231 9983 13257 10009
rect 13257 9983 13258 10009
rect 13230 9982 13258 9983
rect 13342 9926 13370 9954
rect 13790 10065 13818 10066
rect 13790 10039 13791 10065
rect 13791 10039 13817 10065
rect 13817 10039 13818 10065
rect 13790 10038 13818 10039
rect 13846 10710 13874 10738
rect 18830 10793 18858 10794
rect 18830 10767 18831 10793
rect 18831 10767 18857 10793
rect 18857 10767 18858 10793
rect 18830 10766 18858 10767
rect 20006 10766 20034 10794
rect 14574 10737 14602 10738
rect 14574 10711 14575 10737
rect 14575 10711 14601 10737
rect 14601 10711 14602 10737
rect 14574 10710 14602 10711
rect 17598 10597 17626 10598
rect 17598 10571 17599 10597
rect 17599 10571 17625 10597
rect 17625 10571 17626 10597
rect 17598 10570 17626 10571
rect 17650 10597 17678 10598
rect 17650 10571 17651 10597
rect 17651 10571 17677 10597
rect 17677 10571 17678 10597
rect 17650 10570 17678 10571
rect 17702 10597 17730 10598
rect 17702 10571 17703 10597
rect 17703 10571 17729 10597
rect 17729 10571 17730 10597
rect 17702 10570 17730 10571
rect 20006 10457 20034 10458
rect 20006 10431 20007 10457
rect 20007 10431 20033 10457
rect 20033 10431 20034 10457
rect 20006 10430 20034 10431
rect 18830 10401 18858 10402
rect 18830 10375 18831 10401
rect 18831 10375 18857 10401
rect 18857 10375 18858 10401
rect 18830 10374 18858 10375
rect 13902 10038 13930 10066
rect 13510 9926 13538 9954
rect 13678 9617 13706 9618
rect 13678 9591 13679 9617
rect 13679 9591 13705 9617
rect 13705 9591 13706 9617
rect 13678 9590 13706 9591
rect 20006 10038 20034 10066
rect 17598 9813 17626 9814
rect 17598 9787 17599 9813
rect 17599 9787 17625 9813
rect 17625 9787 17626 9813
rect 17598 9786 17626 9787
rect 17650 9813 17678 9814
rect 17650 9787 17651 9813
rect 17651 9787 17677 9813
rect 17677 9787 17678 9813
rect 17650 9786 17678 9787
rect 17702 9813 17730 9814
rect 17702 9787 17703 9813
rect 17703 9787 17729 9813
rect 17729 9787 17730 9813
rect 17702 9786 17730 9787
rect 14574 9617 14602 9618
rect 14574 9591 14575 9617
rect 14575 9591 14601 9617
rect 14601 9591 14602 9617
rect 14574 9590 14602 9591
rect 13286 9366 13314 9394
rect 13062 9086 13090 9114
rect 11830 8582 11858 8610
rect 13510 9310 13538 9338
rect 14854 9590 14882 9618
rect 14742 9505 14770 9506
rect 14742 9479 14743 9505
rect 14743 9479 14769 9505
rect 14769 9479 14770 9505
rect 14742 9478 14770 9479
rect 18774 9478 18802 9506
rect 14854 9198 14882 9226
rect 14686 9169 14714 9170
rect 14686 9143 14687 9169
rect 14687 9143 14713 9169
rect 14713 9143 14714 9169
rect 14686 9142 14714 9143
rect 15190 9225 15218 9226
rect 15190 9199 15191 9225
rect 15191 9199 15217 9225
rect 15217 9199 15218 9225
rect 15190 9198 15218 9199
rect 15022 9142 15050 9170
rect 14742 8721 14770 8722
rect 14742 8695 14743 8721
rect 14743 8695 14769 8721
rect 14769 8695 14770 8721
rect 14742 8694 14770 8695
rect 13230 8582 13258 8610
rect 11718 8414 11746 8442
rect 12222 8414 12250 8442
rect 9918 7069 9946 7070
rect 9918 7043 9919 7069
rect 9919 7043 9945 7069
rect 9945 7043 9946 7069
rect 9918 7042 9946 7043
rect 9970 7069 9998 7070
rect 9970 7043 9971 7069
rect 9971 7043 9997 7069
rect 9997 7043 9998 7069
rect 9970 7042 9998 7043
rect 10022 7069 10050 7070
rect 10022 7043 10023 7069
rect 10023 7043 10049 7069
rect 10049 7043 10050 7069
rect 10022 7042 10050 7043
rect 9918 6285 9946 6286
rect 9918 6259 9919 6285
rect 9919 6259 9945 6285
rect 9945 6259 9946 6285
rect 9918 6258 9946 6259
rect 9970 6285 9998 6286
rect 9970 6259 9971 6285
rect 9971 6259 9997 6285
rect 9997 6259 9998 6285
rect 9970 6258 9998 6259
rect 10022 6285 10050 6286
rect 10022 6259 10023 6285
rect 10023 6259 10049 6285
rect 10049 6259 10050 6285
rect 10022 6258 10050 6259
rect 9918 5501 9946 5502
rect 9918 5475 9919 5501
rect 9919 5475 9945 5501
rect 9945 5475 9946 5501
rect 9918 5474 9946 5475
rect 9970 5501 9998 5502
rect 9970 5475 9971 5501
rect 9971 5475 9997 5501
rect 9997 5475 9998 5501
rect 9970 5474 9998 5475
rect 10022 5501 10050 5502
rect 10022 5475 10023 5501
rect 10023 5475 10049 5501
rect 10049 5475 10050 5501
rect 10022 5474 10050 5475
rect 9918 4717 9946 4718
rect 9918 4691 9919 4717
rect 9919 4691 9945 4717
rect 9945 4691 9946 4717
rect 9918 4690 9946 4691
rect 9970 4717 9998 4718
rect 9970 4691 9971 4717
rect 9971 4691 9997 4717
rect 9997 4691 9998 4717
rect 9970 4690 9998 4691
rect 10022 4717 10050 4718
rect 10022 4691 10023 4717
rect 10023 4691 10049 4717
rect 10049 4691 10050 4717
rect 10022 4690 10050 4691
rect 9918 3933 9946 3934
rect 9918 3907 9919 3933
rect 9919 3907 9945 3933
rect 9945 3907 9946 3933
rect 9918 3906 9946 3907
rect 9970 3933 9998 3934
rect 9970 3907 9971 3933
rect 9971 3907 9997 3933
rect 9997 3907 9998 3933
rect 9970 3906 9998 3907
rect 10022 3933 10050 3934
rect 10022 3907 10023 3933
rect 10023 3907 10049 3933
rect 10049 3907 10050 3933
rect 10022 3906 10050 3907
rect 9918 3149 9946 3150
rect 9918 3123 9919 3149
rect 9919 3123 9945 3149
rect 9945 3123 9946 3149
rect 9918 3122 9946 3123
rect 9970 3149 9998 3150
rect 9970 3123 9971 3149
rect 9971 3123 9997 3149
rect 9997 3123 9998 3149
rect 9970 3122 9998 3123
rect 10022 3149 10050 3150
rect 10022 3123 10023 3149
rect 10023 3123 10049 3149
rect 10049 3123 10050 3149
rect 10022 3122 10050 3123
rect 9918 2365 9946 2366
rect 9918 2339 9919 2365
rect 9919 2339 9945 2365
rect 9945 2339 9946 2365
rect 9918 2338 9946 2339
rect 9970 2365 9998 2366
rect 9970 2339 9971 2365
rect 9971 2339 9997 2365
rect 9997 2339 9998 2365
rect 9970 2338 9998 2339
rect 10022 2365 10050 2366
rect 10022 2339 10023 2365
rect 10023 2339 10049 2365
rect 10049 2339 10050 2365
rect 10022 2338 10050 2339
rect 10430 1806 10458 1834
rect 9918 1581 9946 1582
rect 9918 1555 9919 1581
rect 9919 1555 9945 1581
rect 9945 1555 9946 1581
rect 9918 1554 9946 1555
rect 9970 1581 9998 1582
rect 9970 1555 9971 1581
rect 9971 1555 9997 1581
rect 9997 1555 9998 1581
rect 9970 1554 9998 1555
rect 10022 1581 10050 1582
rect 10022 1555 10023 1581
rect 10023 1555 10049 1581
rect 10049 1555 10050 1581
rect 10022 1554 10050 1555
rect 11774 2590 11802 2618
rect 11046 1833 11074 1834
rect 11046 1807 11047 1833
rect 11047 1807 11073 1833
rect 11073 1807 11074 1833
rect 11046 1806 11074 1807
rect 11438 1806 11466 1834
rect 18718 9142 18746 9170
rect 17598 9029 17626 9030
rect 17598 9003 17599 9029
rect 17599 9003 17625 9029
rect 17625 9003 17626 9029
rect 17598 9002 17626 9003
rect 17650 9029 17678 9030
rect 17650 9003 17651 9029
rect 17651 9003 17677 9029
rect 17677 9003 17678 9029
rect 17650 9002 17678 9003
rect 17702 9029 17730 9030
rect 17702 9003 17703 9029
rect 17703 9003 17729 9029
rect 17729 9003 17730 9029
rect 17702 9002 17730 9003
rect 17598 8245 17626 8246
rect 17598 8219 17599 8245
rect 17599 8219 17625 8245
rect 17625 8219 17626 8245
rect 17598 8218 17626 8219
rect 17650 8245 17678 8246
rect 17650 8219 17651 8245
rect 17651 8219 17677 8245
rect 17677 8219 17678 8245
rect 17650 8218 17678 8219
rect 17702 8245 17730 8246
rect 17702 8219 17703 8245
rect 17703 8219 17729 8245
rect 17729 8219 17730 8245
rect 17702 8218 17730 8219
rect 15358 8022 15386 8050
rect 18830 9422 18858 9450
rect 20006 9758 20034 9786
rect 18942 9366 18970 9394
rect 20006 9422 20034 9450
rect 18830 9225 18858 9226
rect 18830 9199 18831 9225
rect 18831 9199 18857 9225
rect 18857 9199 18858 9225
rect 18830 9198 18858 9199
rect 19950 9086 19978 9114
rect 19670 8750 19698 8778
rect 18830 8694 18858 8722
rect 19894 8358 19922 8386
rect 20006 8078 20034 8106
rect 18830 8049 18858 8050
rect 18830 8023 18831 8049
rect 18831 8023 18857 8049
rect 18857 8023 18858 8049
rect 18830 8022 18858 8023
rect 17598 7461 17626 7462
rect 17598 7435 17599 7461
rect 17599 7435 17625 7461
rect 17625 7435 17626 7461
rect 17598 7434 17626 7435
rect 17650 7461 17678 7462
rect 17650 7435 17651 7461
rect 17651 7435 17677 7461
rect 17677 7435 17678 7461
rect 17650 7434 17678 7435
rect 17702 7461 17730 7462
rect 17702 7435 17703 7461
rect 17703 7435 17729 7461
rect 17729 7435 17730 7461
rect 17702 7434 17730 7435
rect 17598 6677 17626 6678
rect 17598 6651 17599 6677
rect 17599 6651 17625 6677
rect 17625 6651 17626 6677
rect 17598 6650 17626 6651
rect 17650 6677 17678 6678
rect 17650 6651 17651 6677
rect 17651 6651 17677 6677
rect 17677 6651 17678 6677
rect 17650 6650 17678 6651
rect 17702 6677 17730 6678
rect 17702 6651 17703 6677
rect 17703 6651 17729 6677
rect 17729 6651 17730 6677
rect 17702 6650 17730 6651
rect 17598 5893 17626 5894
rect 17598 5867 17599 5893
rect 17599 5867 17625 5893
rect 17625 5867 17626 5893
rect 17598 5866 17626 5867
rect 17650 5893 17678 5894
rect 17650 5867 17651 5893
rect 17651 5867 17677 5893
rect 17677 5867 17678 5893
rect 17650 5866 17678 5867
rect 17702 5893 17730 5894
rect 17702 5867 17703 5893
rect 17703 5867 17729 5893
rect 17729 5867 17730 5893
rect 17702 5866 17730 5867
rect 17598 5109 17626 5110
rect 17598 5083 17599 5109
rect 17599 5083 17625 5109
rect 17625 5083 17626 5109
rect 17598 5082 17626 5083
rect 17650 5109 17678 5110
rect 17650 5083 17651 5109
rect 17651 5083 17677 5109
rect 17677 5083 17678 5109
rect 17650 5082 17678 5083
rect 17702 5109 17730 5110
rect 17702 5083 17703 5109
rect 17703 5083 17729 5109
rect 17729 5083 17730 5109
rect 17702 5082 17730 5083
rect 17598 4325 17626 4326
rect 17598 4299 17599 4325
rect 17599 4299 17625 4325
rect 17625 4299 17626 4325
rect 17598 4298 17626 4299
rect 17650 4325 17678 4326
rect 17650 4299 17651 4325
rect 17651 4299 17677 4325
rect 17677 4299 17678 4325
rect 17650 4298 17678 4299
rect 17702 4325 17730 4326
rect 17702 4299 17703 4325
rect 17703 4299 17729 4325
rect 17729 4299 17730 4325
rect 17702 4298 17730 4299
rect 17598 3541 17626 3542
rect 17598 3515 17599 3541
rect 17599 3515 17625 3541
rect 17625 3515 17626 3541
rect 17598 3514 17626 3515
rect 17650 3541 17678 3542
rect 17650 3515 17651 3541
rect 17651 3515 17677 3541
rect 17677 3515 17678 3541
rect 17650 3514 17678 3515
rect 17702 3541 17730 3542
rect 17702 3515 17703 3541
rect 17703 3515 17729 3541
rect 17729 3515 17730 3541
rect 17702 3514 17730 3515
rect 17598 2757 17626 2758
rect 17598 2731 17599 2757
rect 17599 2731 17625 2757
rect 17625 2731 17626 2757
rect 17598 2730 17626 2731
rect 17650 2757 17678 2758
rect 17650 2731 17651 2757
rect 17651 2731 17677 2757
rect 17677 2731 17678 2757
rect 17650 2730 17678 2731
rect 17702 2757 17730 2758
rect 17702 2731 17703 2757
rect 17703 2731 17729 2757
rect 17729 2731 17730 2757
rect 17702 2730 17730 2731
rect 12390 2617 12418 2618
rect 12390 2591 12391 2617
rect 12391 2591 12417 2617
rect 12417 2591 12418 2617
rect 12390 2590 12418 2591
rect 17598 1973 17626 1974
rect 17598 1947 17599 1973
rect 17599 1947 17625 1973
rect 17625 1947 17626 1973
rect 17598 1946 17626 1947
rect 17650 1973 17678 1974
rect 17650 1947 17651 1973
rect 17651 1947 17677 1973
rect 17677 1947 17678 1973
rect 17650 1946 17678 1947
rect 17702 1973 17730 1974
rect 17702 1947 17703 1973
rect 17703 1947 17729 1973
rect 17729 1947 17730 1973
rect 17702 1946 17730 1947
rect 12782 1833 12810 1834
rect 12782 1807 12783 1833
rect 12783 1807 12809 1833
rect 12809 1807 12810 1833
rect 12782 1806 12810 1807
<< metal3 >>
rect 2233 19194 2238 19222
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2370 19194 2375 19222
rect 17593 19194 17598 19222
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17730 19194 17735 19222
rect 11769 19110 11774 19138
rect 11802 19110 12782 19138
rect 12810 19110 12815 19138
rect 9913 18802 9918 18830
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 10050 18802 10055 18830
rect 12105 18718 12110 18746
rect 12138 18718 13118 18746
rect 13146 18718 13151 18746
rect 2233 18410 2238 18438
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2370 18410 2375 18438
rect 17593 18410 17598 18438
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17730 18410 17735 18438
rect 12553 18326 12558 18354
rect 12586 18326 13062 18354
rect 13090 18326 13095 18354
rect 9913 18018 9918 18046
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 10050 18018 10055 18046
rect 2233 17626 2238 17654
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2370 17626 2375 17654
rect 17593 17626 17598 17654
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17730 17626 17735 17654
rect 9913 17234 9918 17262
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 10050 17234 10055 17262
rect 2233 16842 2238 16870
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2370 16842 2375 16870
rect 17593 16842 17598 16870
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17730 16842 17735 16870
rect 9913 16450 9918 16478
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 10050 16450 10055 16478
rect 2233 16058 2238 16086
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2370 16058 2375 16086
rect 17593 16058 17598 16086
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17730 16058 17735 16086
rect 9913 15666 9918 15694
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 10050 15666 10055 15694
rect 2233 15274 2238 15302
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2370 15274 2375 15302
rect 17593 15274 17598 15302
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17730 15274 17735 15302
rect 9913 14882 9918 14910
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 10050 14882 10055 14910
rect 2233 14490 2238 14518
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2370 14490 2375 14518
rect 17593 14490 17598 14518
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17730 14490 17735 14518
rect 9913 14098 9918 14126
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 10050 14098 10055 14126
rect 2233 13706 2238 13734
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2370 13706 2375 13734
rect 17593 13706 17598 13734
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17730 13706 17735 13734
rect 9913 13314 9918 13342
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 10050 13314 10055 13342
rect 12217 13230 12222 13258
rect 12250 13230 12614 13258
rect 12642 13230 12647 13258
rect 2233 12922 2238 12950
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2370 12922 2375 12950
rect 17593 12922 17598 12950
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17730 12922 17735 12950
rect 0 12810 400 12824
rect 0 12782 2086 12810
rect 2114 12782 2119 12810
rect 0 12768 400 12782
rect 2137 12726 2142 12754
rect 2170 12726 6734 12754
rect 6762 12726 7462 12754
rect 7490 12726 7495 12754
rect 11545 12614 11550 12642
rect 11578 12614 12110 12642
rect 12138 12614 12390 12642
rect 12418 12614 12782 12642
rect 12810 12614 12815 12642
rect 9913 12530 9918 12558
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 10050 12530 10055 12558
rect 0 12474 400 12488
rect 0 12446 966 12474
rect 994 12446 999 12474
rect 7513 12446 7518 12474
rect 7546 12446 8078 12474
rect 8106 12446 8358 12474
rect 8386 12446 8638 12474
rect 8666 12446 8671 12474
rect 0 12432 400 12446
rect 6230 12390 7966 12418
rect 7994 12390 7999 12418
rect 6230 12362 6258 12390
rect 2137 12334 2142 12362
rect 2170 12334 6230 12362
rect 6258 12334 6263 12362
rect 8465 12334 8470 12362
rect 8498 12334 8974 12362
rect 9002 12334 9007 12362
rect 9753 12334 9758 12362
rect 9786 12334 11382 12362
rect 11410 12334 11942 12362
rect 11970 12334 11975 12362
rect 12161 12334 12166 12362
rect 12194 12334 13006 12362
rect 13034 12334 13039 12362
rect 7513 12278 7518 12306
rect 7546 12278 7910 12306
rect 7938 12278 7943 12306
rect 961 12222 966 12250
rect 994 12222 999 12250
rect 0 12138 400 12152
rect 966 12138 994 12222
rect 10537 12166 10542 12194
rect 10570 12166 11830 12194
rect 11858 12166 11863 12194
rect 2233 12138 2238 12166
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2370 12138 2375 12166
rect 17593 12138 17598 12166
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17730 12138 17735 12166
rect 20600 12138 21000 12152
rect 0 12110 994 12138
rect 20001 12110 20006 12138
rect 20034 12110 21000 12138
rect 0 12096 400 12110
rect 20600 12096 21000 12110
rect 9697 12054 9702 12082
rect 9730 12054 10150 12082
rect 10178 12054 10183 12082
rect 7681 11998 7686 12026
rect 7714 11998 8190 12026
rect 8218 11998 8414 12026
rect 8442 11998 8694 12026
rect 8722 11998 8727 12026
rect 12777 11998 12782 12026
rect 12810 11998 18830 12026
rect 18858 11998 18863 12026
rect 13006 11970 13034 11998
rect 7849 11942 7854 11970
rect 7882 11942 9310 11970
rect 9338 11942 10542 11970
rect 10570 11942 10575 11970
rect 13001 11942 13006 11970
rect 13034 11942 13039 11970
rect 9193 11886 9198 11914
rect 9226 11886 9758 11914
rect 9786 11886 9791 11914
rect 7233 11774 7238 11802
rect 7266 11774 8302 11802
rect 8330 11774 8750 11802
rect 8778 11774 8783 11802
rect 9913 11746 9918 11774
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 10050 11746 10055 11774
rect 7177 11662 7182 11690
rect 7210 11662 7350 11690
rect 7378 11662 7686 11690
rect 7714 11662 7966 11690
rect 7994 11662 7999 11690
rect 9361 11662 9366 11690
rect 9394 11662 9926 11690
rect 9954 11662 10710 11690
rect 10738 11662 10743 11690
rect 7401 11606 7406 11634
rect 7434 11606 7798 11634
rect 7826 11606 7831 11634
rect 13057 11606 13062 11634
rect 13090 11606 13846 11634
rect 13874 11606 13879 11634
rect 2137 11550 2142 11578
rect 2170 11550 5670 11578
rect 5698 11550 7294 11578
rect 7322 11550 7327 11578
rect 8857 11550 8862 11578
rect 8890 11550 9310 11578
rect 9338 11550 9343 11578
rect 13785 11550 13790 11578
rect 13818 11550 14294 11578
rect 14322 11550 18830 11578
rect 18858 11550 18863 11578
rect 0 11466 400 11480
rect 20600 11466 21000 11480
rect 0 11438 966 11466
rect 994 11438 999 11466
rect 20001 11438 20006 11466
rect 20034 11438 21000 11466
rect 0 11424 400 11438
rect 20600 11424 21000 11438
rect 2233 11354 2238 11382
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2370 11354 2375 11382
rect 17593 11354 17598 11382
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17730 11354 17735 11382
rect 10985 11270 10990 11298
rect 11018 11270 11662 11298
rect 11690 11270 11695 11298
rect 2137 11158 2142 11186
rect 2170 11158 6734 11186
rect 6762 11158 6767 11186
rect 7009 11158 7014 11186
rect 7042 11158 7406 11186
rect 7434 11158 7439 11186
rect 9641 11158 9646 11186
rect 9674 11158 10766 11186
rect 10794 11158 10799 11186
rect 20600 11130 21000 11144
rect 20001 11102 20006 11130
rect 20034 11102 21000 11130
rect 20600 11088 21000 11102
rect 9913 10962 9918 10990
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 10050 10962 10055 10990
rect 10761 10878 10766 10906
rect 10794 10878 11662 10906
rect 11690 10878 11695 10906
rect 15946 10878 18830 10906
rect 18858 10878 18863 10906
rect 15946 10850 15974 10878
rect 10089 10822 10094 10850
rect 10122 10822 10822 10850
rect 10850 10822 11214 10850
rect 11242 10822 11247 10850
rect 14905 10822 14910 10850
rect 14938 10822 15974 10850
rect 0 10794 400 10808
rect 20600 10794 21000 10808
rect 0 10766 966 10794
rect 994 10766 999 10794
rect 7457 10766 7462 10794
rect 7490 10766 8134 10794
rect 8162 10766 8167 10794
rect 8241 10766 8246 10794
rect 8274 10766 8974 10794
rect 9002 10766 9758 10794
rect 9786 10766 10150 10794
rect 10178 10766 10183 10794
rect 10929 10766 10934 10794
rect 10962 10766 11382 10794
rect 11410 10766 12838 10794
rect 12866 10766 13174 10794
rect 13202 10766 13207 10794
rect 14793 10766 14798 10794
rect 14826 10766 18830 10794
rect 18858 10766 18863 10794
rect 20001 10766 20006 10794
rect 20034 10766 21000 10794
rect 0 10752 400 10766
rect 20600 10752 21000 10766
rect 6785 10710 6790 10738
rect 6818 10710 7574 10738
rect 7602 10710 7607 10738
rect 7737 10710 7742 10738
rect 7770 10710 9422 10738
rect 9450 10710 9455 10738
rect 11825 10710 11830 10738
rect 11858 10710 12334 10738
rect 12362 10710 12367 10738
rect 13841 10710 13846 10738
rect 13874 10710 14574 10738
rect 14602 10710 14607 10738
rect 2233 10570 2238 10598
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2370 10570 2375 10598
rect 17593 10570 17598 10598
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17730 10570 17735 10598
rect 20600 10458 21000 10472
rect 20001 10430 20006 10458
rect 20034 10430 21000 10458
rect 20600 10416 21000 10430
rect 10033 10374 10038 10402
rect 10066 10374 11662 10402
rect 11690 10374 11695 10402
rect 12329 10374 12334 10402
rect 12362 10374 18830 10402
rect 18858 10374 18863 10402
rect 8129 10318 8134 10346
rect 8162 10318 8414 10346
rect 8442 10318 8447 10346
rect 10374 10318 11046 10346
rect 11074 10318 11079 10346
rect 10374 10290 10402 10318
rect 9753 10262 9758 10290
rect 9786 10262 10374 10290
rect 10402 10262 10407 10290
rect 10705 10262 10710 10290
rect 10738 10262 11382 10290
rect 11410 10262 11415 10290
rect 9913 10178 9918 10206
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 10050 10178 10055 10206
rect 20600 10122 21000 10136
rect 9641 10094 9646 10122
rect 9674 10094 10038 10122
rect 10066 10094 10071 10122
rect 20006 10094 21000 10122
rect 20006 10066 20034 10094
rect 20600 10080 21000 10094
rect 12777 10038 12782 10066
rect 12810 10038 13790 10066
rect 13818 10038 13902 10066
rect 13930 10038 13935 10066
rect 20001 10038 20006 10066
rect 20034 10038 20039 10066
rect 7009 9982 7014 10010
rect 7042 9982 8134 10010
rect 8162 9982 8167 10010
rect 9305 9982 9310 10010
rect 9338 9982 9702 10010
rect 9730 9982 9735 10010
rect 10089 9982 10094 10010
rect 10122 9982 13230 10010
rect 13258 9982 13454 10010
rect 13426 9954 13454 9982
rect 7961 9926 7966 9954
rect 7994 9926 11326 9954
rect 11354 9926 13342 9954
rect 13370 9926 13375 9954
rect 13426 9926 13510 9954
rect 13538 9926 13543 9954
rect 8745 9870 8750 9898
rect 8778 9870 9478 9898
rect 9506 9870 9511 9898
rect 2233 9786 2238 9814
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2370 9786 2375 9814
rect 17593 9786 17598 9814
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17730 9786 17735 9814
rect 20600 9786 21000 9800
rect 20001 9758 20006 9786
rect 20034 9758 21000 9786
rect 20600 9744 21000 9758
rect 9529 9702 9534 9730
rect 9562 9702 9814 9730
rect 9842 9702 9847 9730
rect 10257 9702 10262 9730
rect 10290 9702 10990 9730
rect 11018 9702 12054 9730
rect 12082 9702 12087 9730
rect 8409 9646 8414 9674
rect 8442 9646 9422 9674
rect 9450 9646 9455 9674
rect 9697 9590 9702 9618
rect 9730 9590 10094 9618
rect 10122 9590 11998 9618
rect 12026 9590 12138 9618
rect 13673 9590 13678 9618
rect 13706 9590 14574 9618
rect 14602 9590 14854 9618
rect 14882 9590 14887 9618
rect 8913 9534 8918 9562
rect 8946 9534 10822 9562
rect 10850 9534 11102 9562
rect 11130 9534 11135 9562
rect 12110 9506 12138 9590
rect 12217 9534 12222 9562
rect 12250 9534 12894 9562
rect 12922 9534 12927 9562
rect 2081 9478 2086 9506
rect 2114 9478 9310 9506
rect 9338 9478 9343 9506
rect 9473 9478 9478 9506
rect 9506 9478 9926 9506
rect 9954 9478 9959 9506
rect 12110 9478 12334 9506
rect 12362 9478 12670 9506
rect 12698 9478 12703 9506
rect 13057 9478 13062 9506
rect 13090 9478 13454 9506
rect 14737 9478 14742 9506
rect 14770 9478 18774 9506
rect 18802 9478 18807 9506
rect 13426 9450 13454 9478
rect 20600 9450 21000 9464
rect 13426 9422 18830 9450
rect 18858 9422 18863 9450
rect 20001 9422 20006 9450
rect 20034 9422 21000 9450
rect 9913 9394 9918 9422
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 10050 9394 10055 9422
rect 20600 9408 21000 9422
rect 12889 9366 12894 9394
rect 12922 9366 13286 9394
rect 13314 9366 18942 9394
rect 18970 9366 18975 9394
rect 6953 9310 6958 9338
rect 6986 9310 7574 9338
rect 7602 9310 9422 9338
rect 9450 9310 9455 9338
rect 9641 9310 9646 9338
rect 9674 9310 9870 9338
rect 9898 9310 10654 9338
rect 10682 9310 10687 9338
rect 11657 9310 11662 9338
rect 11690 9310 12614 9338
rect 12642 9310 13510 9338
rect 13538 9310 13543 9338
rect 7681 9254 7686 9282
rect 7714 9254 7966 9282
rect 7994 9254 7999 9282
rect 8913 9254 8918 9282
rect 8946 9254 9254 9282
rect 9282 9254 9287 9282
rect 9585 9254 9590 9282
rect 9618 9254 9926 9282
rect 9954 9254 9959 9282
rect 7401 9198 7406 9226
rect 7434 9198 7798 9226
rect 7826 9198 7831 9226
rect 9529 9198 9534 9226
rect 9562 9198 10766 9226
rect 10794 9198 10799 9226
rect 14849 9198 14854 9226
rect 14882 9198 15190 9226
rect 15218 9198 15223 9226
rect 18825 9198 18830 9226
rect 18858 9198 18863 9226
rect 2137 9142 2142 9170
rect 2170 9142 5782 9170
rect 5810 9142 5815 9170
rect 6841 9142 6846 9170
rect 6874 9142 7630 9170
rect 7658 9142 7663 9170
rect 10033 9142 10038 9170
rect 10066 9142 10934 9170
rect 10962 9142 10967 9170
rect 14681 9142 14686 9170
rect 14714 9142 15022 9170
rect 15050 9142 18718 9170
rect 18746 9142 18751 9170
rect 0 9114 400 9128
rect 18830 9114 18858 9198
rect 20600 9114 21000 9128
rect 0 9086 966 9114
rect 994 9086 999 9114
rect 6897 9086 6902 9114
rect 6930 9086 7910 9114
rect 7938 9086 7943 9114
rect 13057 9086 13062 9114
rect 13090 9086 18858 9114
rect 19945 9086 19950 9114
rect 19978 9086 21000 9114
rect 0 9072 400 9086
rect 20600 9072 21000 9086
rect 2233 9002 2238 9030
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2370 9002 2375 9030
rect 17593 9002 17598 9030
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17730 9002 17735 9030
rect 7905 8918 7910 8946
rect 7938 8918 8862 8946
rect 8890 8918 8895 8946
rect 2137 8806 2142 8834
rect 2170 8806 6006 8834
rect 6034 8806 6039 8834
rect 9081 8806 9086 8834
rect 9114 8806 9758 8834
rect 9786 8806 9870 8834
rect 9898 8806 9903 8834
rect 20600 8778 21000 8792
rect 5777 8750 5782 8778
rect 5810 8750 7462 8778
rect 7490 8750 7495 8778
rect 8913 8750 8918 8778
rect 8946 8750 9198 8778
rect 9226 8750 9366 8778
rect 9394 8750 10206 8778
rect 10234 8750 10239 8778
rect 19665 8750 19670 8778
rect 19698 8750 21000 8778
rect 20600 8736 21000 8750
rect 7065 8694 7070 8722
rect 7098 8694 7574 8722
rect 7602 8694 7607 8722
rect 8857 8694 8862 8722
rect 8890 8694 9478 8722
rect 9506 8694 9511 8722
rect 14737 8694 14742 8722
rect 14770 8694 18830 8722
rect 18858 8694 18863 8722
rect 7513 8638 7518 8666
rect 7546 8638 7826 8666
rect 6001 8526 6006 8554
rect 6034 8526 7686 8554
rect 7714 8526 7719 8554
rect 7798 8498 7826 8638
rect 9913 8610 9918 8638
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 10050 8610 10055 8638
rect 10817 8582 10822 8610
rect 10850 8582 11830 8610
rect 11858 8582 13230 8610
rect 13258 8582 13263 8610
rect 7737 8470 7742 8498
rect 7770 8470 8302 8498
rect 8330 8470 10934 8498
rect 10962 8470 10967 8498
rect 0 8442 400 8456
rect 20600 8442 21000 8456
rect 0 8414 966 8442
rect 994 8414 999 8442
rect 8465 8414 8470 8442
rect 8498 8414 8918 8442
rect 8946 8414 8951 8442
rect 9921 8414 9926 8442
rect 9954 8414 10150 8442
rect 10178 8414 10183 8442
rect 11097 8414 11102 8442
rect 11130 8414 11718 8442
rect 11746 8414 12222 8442
rect 12250 8414 12255 8442
rect 19950 8414 21000 8442
rect 0 8400 400 8414
rect 19950 8386 19978 8414
rect 20600 8400 21000 8414
rect 19889 8358 19894 8386
rect 19922 8358 19978 8386
rect 7233 8302 7238 8330
rect 7266 8302 8974 8330
rect 9002 8302 9007 8330
rect 2233 8218 2238 8246
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2370 8218 2375 8246
rect 17593 8218 17598 8246
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17730 8218 17735 8246
rect 20600 8106 21000 8120
rect 8297 8078 8302 8106
rect 8330 8078 8806 8106
rect 8834 8078 8839 8106
rect 20001 8078 20006 8106
rect 20034 8078 21000 8106
rect 20600 8064 21000 8078
rect 6897 8022 6902 8050
rect 6930 8022 7182 8050
rect 7210 8022 7518 8050
rect 7546 8022 8526 8050
rect 8554 8022 8559 8050
rect 15353 8022 15358 8050
rect 15386 8022 18830 8050
rect 18858 8022 18863 8050
rect 9913 7826 9918 7854
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 10050 7826 10055 7854
rect 8521 7630 8526 7658
rect 8554 7630 9422 7658
rect 9450 7630 9455 7658
rect 2233 7434 2238 7462
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2370 7434 2375 7462
rect 17593 7434 17598 7462
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17730 7434 17735 7462
rect 9913 7042 9918 7070
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 10050 7042 10055 7070
rect 2233 6650 2238 6678
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2370 6650 2375 6678
rect 17593 6650 17598 6678
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17730 6650 17735 6678
rect 9913 6258 9918 6286
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 10050 6258 10055 6286
rect 2233 5866 2238 5894
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2370 5866 2375 5894
rect 17593 5866 17598 5894
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17730 5866 17735 5894
rect 9913 5474 9918 5502
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 10050 5474 10055 5502
rect 2233 5082 2238 5110
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2370 5082 2375 5110
rect 17593 5082 17598 5110
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17730 5082 17735 5110
rect 9913 4690 9918 4718
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 10050 4690 10055 4718
rect 2233 4298 2238 4326
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2370 4298 2375 4326
rect 17593 4298 17598 4326
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17730 4298 17735 4326
rect 9913 3906 9918 3934
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 10050 3906 10055 3934
rect 2233 3514 2238 3542
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2370 3514 2375 3542
rect 17593 3514 17598 3542
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17730 3514 17735 3542
rect 9913 3122 9918 3150
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 10050 3122 10055 3150
rect 2233 2730 2238 2758
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2370 2730 2375 2758
rect 17593 2730 17598 2758
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17730 2730 17735 2758
rect 11769 2590 11774 2618
rect 11802 2590 12390 2618
rect 12418 2590 12423 2618
rect 9913 2338 9918 2366
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 10050 2338 10055 2366
rect 2233 1946 2238 1974
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2370 1946 2375 1974
rect 17593 1946 17598 1974
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17730 1946 17735 1974
rect 10425 1806 10430 1834
rect 10458 1806 11046 1834
rect 11074 1806 11079 1834
rect 11433 1806 11438 1834
rect 11466 1806 12782 1834
rect 12810 1806 12815 1834
rect 9913 1554 9918 1582
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 10050 1554 10055 1582
<< via3 >>
rect 2238 19194 2266 19222
rect 2290 19194 2318 19222
rect 2342 19194 2370 19222
rect 17598 19194 17626 19222
rect 17650 19194 17678 19222
rect 17702 19194 17730 19222
rect 9918 18802 9946 18830
rect 9970 18802 9998 18830
rect 10022 18802 10050 18830
rect 2238 18410 2266 18438
rect 2290 18410 2318 18438
rect 2342 18410 2370 18438
rect 17598 18410 17626 18438
rect 17650 18410 17678 18438
rect 17702 18410 17730 18438
rect 9918 18018 9946 18046
rect 9970 18018 9998 18046
rect 10022 18018 10050 18046
rect 2238 17626 2266 17654
rect 2290 17626 2318 17654
rect 2342 17626 2370 17654
rect 17598 17626 17626 17654
rect 17650 17626 17678 17654
rect 17702 17626 17730 17654
rect 9918 17234 9946 17262
rect 9970 17234 9998 17262
rect 10022 17234 10050 17262
rect 2238 16842 2266 16870
rect 2290 16842 2318 16870
rect 2342 16842 2370 16870
rect 17598 16842 17626 16870
rect 17650 16842 17678 16870
rect 17702 16842 17730 16870
rect 9918 16450 9946 16478
rect 9970 16450 9998 16478
rect 10022 16450 10050 16478
rect 2238 16058 2266 16086
rect 2290 16058 2318 16086
rect 2342 16058 2370 16086
rect 17598 16058 17626 16086
rect 17650 16058 17678 16086
rect 17702 16058 17730 16086
rect 9918 15666 9946 15694
rect 9970 15666 9998 15694
rect 10022 15666 10050 15694
rect 2238 15274 2266 15302
rect 2290 15274 2318 15302
rect 2342 15274 2370 15302
rect 17598 15274 17626 15302
rect 17650 15274 17678 15302
rect 17702 15274 17730 15302
rect 9918 14882 9946 14910
rect 9970 14882 9998 14910
rect 10022 14882 10050 14910
rect 2238 14490 2266 14518
rect 2290 14490 2318 14518
rect 2342 14490 2370 14518
rect 17598 14490 17626 14518
rect 17650 14490 17678 14518
rect 17702 14490 17730 14518
rect 9918 14098 9946 14126
rect 9970 14098 9998 14126
rect 10022 14098 10050 14126
rect 2238 13706 2266 13734
rect 2290 13706 2318 13734
rect 2342 13706 2370 13734
rect 17598 13706 17626 13734
rect 17650 13706 17678 13734
rect 17702 13706 17730 13734
rect 9918 13314 9946 13342
rect 9970 13314 9998 13342
rect 10022 13314 10050 13342
rect 2238 12922 2266 12950
rect 2290 12922 2318 12950
rect 2342 12922 2370 12950
rect 17598 12922 17626 12950
rect 17650 12922 17678 12950
rect 17702 12922 17730 12950
rect 9918 12530 9946 12558
rect 9970 12530 9998 12558
rect 10022 12530 10050 12558
rect 2238 12138 2266 12166
rect 2290 12138 2318 12166
rect 2342 12138 2370 12166
rect 17598 12138 17626 12166
rect 17650 12138 17678 12166
rect 17702 12138 17730 12166
rect 9918 11746 9946 11774
rect 9970 11746 9998 11774
rect 10022 11746 10050 11774
rect 2238 11354 2266 11382
rect 2290 11354 2318 11382
rect 2342 11354 2370 11382
rect 17598 11354 17626 11382
rect 17650 11354 17678 11382
rect 17702 11354 17730 11382
rect 9918 10962 9946 10990
rect 9970 10962 9998 10990
rect 10022 10962 10050 10990
rect 2238 10570 2266 10598
rect 2290 10570 2318 10598
rect 2342 10570 2370 10598
rect 17598 10570 17626 10598
rect 17650 10570 17678 10598
rect 17702 10570 17730 10598
rect 9918 10178 9946 10206
rect 9970 10178 9998 10206
rect 10022 10178 10050 10206
rect 2238 9786 2266 9814
rect 2290 9786 2318 9814
rect 2342 9786 2370 9814
rect 17598 9786 17626 9814
rect 17650 9786 17678 9814
rect 17702 9786 17730 9814
rect 9918 9394 9946 9422
rect 9970 9394 9998 9422
rect 10022 9394 10050 9422
rect 2238 9002 2266 9030
rect 2290 9002 2318 9030
rect 2342 9002 2370 9030
rect 17598 9002 17626 9030
rect 17650 9002 17678 9030
rect 17702 9002 17730 9030
rect 9918 8610 9946 8638
rect 9970 8610 9998 8638
rect 10022 8610 10050 8638
rect 2238 8218 2266 8246
rect 2290 8218 2318 8246
rect 2342 8218 2370 8246
rect 17598 8218 17626 8246
rect 17650 8218 17678 8246
rect 17702 8218 17730 8246
rect 9918 7826 9946 7854
rect 9970 7826 9998 7854
rect 10022 7826 10050 7854
rect 2238 7434 2266 7462
rect 2290 7434 2318 7462
rect 2342 7434 2370 7462
rect 17598 7434 17626 7462
rect 17650 7434 17678 7462
rect 17702 7434 17730 7462
rect 9918 7042 9946 7070
rect 9970 7042 9998 7070
rect 10022 7042 10050 7070
rect 2238 6650 2266 6678
rect 2290 6650 2318 6678
rect 2342 6650 2370 6678
rect 17598 6650 17626 6678
rect 17650 6650 17678 6678
rect 17702 6650 17730 6678
rect 9918 6258 9946 6286
rect 9970 6258 9998 6286
rect 10022 6258 10050 6286
rect 2238 5866 2266 5894
rect 2290 5866 2318 5894
rect 2342 5866 2370 5894
rect 17598 5866 17626 5894
rect 17650 5866 17678 5894
rect 17702 5866 17730 5894
rect 9918 5474 9946 5502
rect 9970 5474 9998 5502
rect 10022 5474 10050 5502
rect 2238 5082 2266 5110
rect 2290 5082 2318 5110
rect 2342 5082 2370 5110
rect 17598 5082 17626 5110
rect 17650 5082 17678 5110
rect 17702 5082 17730 5110
rect 9918 4690 9946 4718
rect 9970 4690 9998 4718
rect 10022 4690 10050 4718
rect 2238 4298 2266 4326
rect 2290 4298 2318 4326
rect 2342 4298 2370 4326
rect 17598 4298 17626 4326
rect 17650 4298 17678 4326
rect 17702 4298 17730 4326
rect 9918 3906 9946 3934
rect 9970 3906 9998 3934
rect 10022 3906 10050 3934
rect 2238 3514 2266 3542
rect 2290 3514 2318 3542
rect 2342 3514 2370 3542
rect 17598 3514 17626 3542
rect 17650 3514 17678 3542
rect 17702 3514 17730 3542
rect 9918 3122 9946 3150
rect 9970 3122 9998 3150
rect 10022 3122 10050 3150
rect 2238 2730 2266 2758
rect 2290 2730 2318 2758
rect 2342 2730 2370 2758
rect 17598 2730 17626 2758
rect 17650 2730 17678 2758
rect 17702 2730 17730 2758
rect 9918 2338 9946 2366
rect 9970 2338 9998 2366
rect 10022 2338 10050 2366
rect 2238 1946 2266 1974
rect 2290 1946 2318 1974
rect 2342 1946 2370 1974
rect 17598 1946 17626 1974
rect 17650 1946 17678 1974
rect 17702 1946 17730 1974
rect 9918 1554 9946 1582
rect 9970 1554 9998 1582
rect 10022 1554 10050 1582
<< metal4 >>
rect 2224 19222 2384 19238
rect 2224 19194 2238 19222
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2370 19194 2384 19222
rect 2224 18438 2384 19194
rect 2224 18410 2238 18438
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2370 18410 2384 18438
rect 2224 17654 2384 18410
rect 2224 17626 2238 17654
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2370 17626 2384 17654
rect 2224 16870 2384 17626
rect 2224 16842 2238 16870
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2370 16842 2384 16870
rect 2224 16086 2384 16842
rect 2224 16058 2238 16086
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2370 16058 2384 16086
rect 2224 15302 2384 16058
rect 2224 15274 2238 15302
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2370 15274 2384 15302
rect 2224 14518 2384 15274
rect 2224 14490 2238 14518
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2370 14490 2384 14518
rect 2224 13734 2384 14490
rect 2224 13706 2238 13734
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2370 13706 2384 13734
rect 2224 12950 2384 13706
rect 2224 12922 2238 12950
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2370 12922 2384 12950
rect 2224 12166 2384 12922
rect 2224 12138 2238 12166
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2370 12138 2384 12166
rect 2224 11382 2384 12138
rect 2224 11354 2238 11382
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2370 11354 2384 11382
rect 2224 10598 2384 11354
rect 2224 10570 2238 10598
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2370 10570 2384 10598
rect 2224 9814 2384 10570
rect 2224 9786 2238 9814
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2370 9786 2384 9814
rect 2224 9030 2384 9786
rect 2224 9002 2238 9030
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2370 9002 2384 9030
rect 2224 8246 2384 9002
rect 2224 8218 2238 8246
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2370 8218 2384 8246
rect 2224 7462 2384 8218
rect 2224 7434 2238 7462
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2370 7434 2384 7462
rect 2224 6678 2384 7434
rect 2224 6650 2238 6678
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2370 6650 2384 6678
rect 2224 5894 2384 6650
rect 2224 5866 2238 5894
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2370 5866 2384 5894
rect 2224 5110 2384 5866
rect 2224 5082 2238 5110
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2370 5082 2384 5110
rect 2224 4326 2384 5082
rect 2224 4298 2238 4326
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2370 4298 2384 4326
rect 2224 3542 2384 4298
rect 2224 3514 2238 3542
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2370 3514 2384 3542
rect 2224 2758 2384 3514
rect 2224 2730 2238 2758
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2370 2730 2384 2758
rect 2224 1974 2384 2730
rect 2224 1946 2238 1974
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2370 1946 2384 1974
rect 2224 1538 2384 1946
rect 9904 18830 10064 19238
rect 9904 18802 9918 18830
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 10050 18802 10064 18830
rect 9904 18046 10064 18802
rect 9904 18018 9918 18046
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 10050 18018 10064 18046
rect 9904 17262 10064 18018
rect 9904 17234 9918 17262
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 10050 17234 10064 17262
rect 9904 16478 10064 17234
rect 9904 16450 9918 16478
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 10050 16450 10064 16478
rect 9904 15694 10064 16450
rect 9904 15666 9918 15694
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 10050 15666 10064 15694
rect 9904 14910 10064 15666
rect 9904 14882 9918 14910
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 10050 14882 10064 14910
rect 9904 14126 10064 14882
rect 9904 14098 9918 14126
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 10050 14098 10064 14126
rect 9904 13342 10064 14098
rect 9904 13314 9918 13342
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 10050 13314 10064 13342
rect 9904 12558 10064 13314
rect 9904 12530 9918 12558
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 10050 12530 10064 12558
rect 9904 11774 10064 12530
rect 9904 11746 9918 11774
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 10050 11746 10064 11774
rect 9904 10990 10064 11746
rect 9904 10962 9918 10990
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 10050 10962 10064 10990
rect 9904 10206 10064 10962
rect 9904 10178 9918 10206
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 10050 10178 10064 10206
rect 9904 9422 10064 10178
rect 9904 9394 9918 9422
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 10050 9394 10064 9422
rect 9904 8638 10064 9394
rect 9904 8610 9918 8638
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 10050 8610 10064 8638
rect 9904 7854 10064 8610
rect 9904 7826 9918 7854
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 10050 7826 10064 7854
rect 9904 7070 10064 7826
rect 9904 7042 9918 7070
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 10050 7042 10064 7070
rect 9904 6286 10064 7042
rect 9904 6258 9918 6286
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 10050 6258 10064 6286
rect 9904 5502 10064 6258
rect 9904 5474 9918 5502
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 10050 5474 10064 5502
rect 9904 4718 10064 5474
rect 9904 4690 9918 4718
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 10050 4690 10064 4718
rect 9904 3934 10064 4690
rect 9904 3906 9918 3934
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 10050 3906 10064 3934
rect 9904 3150 10064 3906
rect 9904 3122 9918 3150
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 10050 3122 10064 3150
rect 9904 2366 10064 3122
rect 9904 2338 9918 2366
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 10050 2338 10064 2366
rect 9904 1582 10064 2338
rect 9904 1554 9918 1582
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 10050 1554 10064 1582
rect 9904 1538 10064 1554
rect 17584 19222 17744 19238
rect 17584 19194 17598 19222
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17730 19194 17744 19222
rect 17584 18438 17744 19194
rect 17584 18410 17598 18438
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17730 18410 17744 18438
rect 17584 17654 17744 18410
rect 17584 17626 17598 17654
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17730 17626 17744 17654
rect 17584 16870 17744 17626
rect 17584 16842 17598 16870
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17730 16842 17744 16870
rect 17584 16086 17744 16842
rect 17584 16058 17598 16086
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17730 16058 17744 16086
rect 17584 15302 17744 16058
rect 17584 15274 17598 15302
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17730 15274 17744 15302
rect 17584 14518 17744 15274
rect 17584 14490 17598 14518
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17730 14490 17744 14518
rect 17584 13734 17744 14490
rect 17584 13706 17598 13734
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17730 13706 17744 13734
rect 17584 12950 17744 13706
rect 17584 12922 17598 12950
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17730 12922 17744 12950
rect 17584 12166 17744 12922
rect 17584 12138 17598 12166
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17730 12138 17744 12166
rect 17584 11382 17744 12138
rect 17584 11354 17598 11382
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17730 11354 17744 11382
rect 17584 10598 17744 11354
rect 17584 10570 17598 10598
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17730 10570 17744 10598
rect 17584 9814 17744 10570
rect 17584 9786 17598 9814
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17730 9786 17744 9814
rect 17584 9030 17744 9786
rect 17584 9002 17598 9030
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17730 9002 17744 9030
rect 17584 8246 17744 9002
rect 17584 8218 17598 8246
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17730 8218 17744 8246
rect 17584 7462 17744 8218
rect 17584 7434 17598 7462
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17730 7434 17744 7462
rect 17584 6678 17744 7434
rect 17584 6650 17598 6678
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17730 6650 17744 6678
rect 17584 5894 17744 6650
rect 17584 5866 17598 5894
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17730 5866 17744 5894
rect 17584 5110 17744 5866
rect 17584 5082 17598 5110
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17730 5082 17744 5110
rect 17584 4326 17744 5082
rect 17584 4298 17598 4326
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17730 4298 17744 4326
rect 17584 3542 17744 4298
rect 17584 3514 17598 3542
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17730 3514 17744 3542
rect 17584 2758 17744 3514
rect 17584 2730 17598 2758
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17730 2730 17744 2758
rect 17584 1974 17744 2730
rect 17584 1946 17598 1974
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17730 1946 17744 1974
rect 17584 1538 17744 1946
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _067_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 10360 0 1 9408
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _068_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9688 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _069_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 13720 0 -1 10192
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _070_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 13160 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _071_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 11872 0 -1 9408
box -43 -43 2115 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _072_
timestamp 1698175906
transform -1 0 13888 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _073_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 14224 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _074_
timestamp 1698175906
transform 1 0 10864 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _075_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 11312 0 -1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _076_
timestamp 1698175906
transform -1 0 13944 0 -1 11760
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _077_
timestamp 1698175906
transform -1 0 13608 0 -1 11760
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _078_
timestamp 1698175906
transform -1 0 7840 0 -1 8624
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _079_
timestamp 1698175906
transform 1 0 6776 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _080_
timestamp 1698175906
transform 1 0 7448 0 -1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _081_
timestamp 1698175906
transform 1 0 7616 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _082_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 10808 0 -1 10976
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _083_
timestamp 1698175906
transform 1 0 11312 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _084_
timestamp 1698175906
transform -1 0 11312 0 -1 12544
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _085_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 12432 0 1 9408
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _086_
timestamp 1698175906
transform 1 0 12432 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _087_
timestamp 1698175906
transform -1 0 12040 0 1 10976
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _088_
timestamp 1698175906
transform 1 0 11088 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _089_
timestamp 1698175906
transform -1 0 7616 0 1 8624
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _090_
timestamp 1698175906
transform -1 0 7784 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _091_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 10472 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _092_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 10080 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _093_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 8288 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _094_
timestamp 1698175906
transform 1 0 7560 0 -1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _095_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 9632 0 -1 10192
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _096_
timestamp 1698175906
transform -1 0 9800 0 -1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _097_
timestamp 1698175906
transform -1 0 8960 0 1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _098_
timestamp 1698175906
transform 1 0 7784 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _099_
timestamp 1698175906
transform 1 0 7168 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _100_
timestamp 1698175906
transform 1 0 9576 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _101_
timestamp 1698175906
transform -1 0 9296 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _102_
timestamp 1698175906
transform 1 0 9240 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _103_
timestamp 1698175906
transform -1 0 10024 0 1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _104_
timestamp 1698175906
transform -1 0 10080 0 -1 11760
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _105_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10248 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _106_
timestamp 1698175906
transform 1 0 10584 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _107_
timestamp 1698175906
transform 1 0 8232 0 -1 8624
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _108_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8848 0 -1 8624
box -43 -43 659 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _109_
timestamp 1698175906
transform -1 0 9688 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _110_
timestamp 1698175906
transform -1 0 9016 0 1 8624
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _111_
timestamp 1698175906
transform 1 0 7112 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _112_
timestamp 1698175906
transform 1 0 6776 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _113_
timestamp 1698175906
transform 1 0 9352 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _114_
timestamp 1698175906
transform 1 0 10584 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _115_
timestamp 1698175906
transform 1 0 10976 0 1 10192
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _116_
timestamp 1698175906
transform -1 0 9744 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _117_
timestamp 1698175906
transform 1 0 7392 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _118_
timestamp 1698175906
transform -1 0 7672 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _119_
timestamp 1698175906
transform -1 0 8064 0 -1 9408
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _120_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 10808 0 -1 11760
box -43 -43 771 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _121_
timestamp 1698175906
transform 1 0 8232 0 -1 12544
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _122_
timestamp 1698175906
transform -1 0 9408 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _123_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10584 0 1 10976
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _124_
timestamp 1698175906
transform -1 0 11088 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _125_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8624 0 -1 10976
box -43 -43 715 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _126_
timestamp 1698175906
transform -1 0 9128 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _127_
timestamp 1698175906
transform 1 0 9464 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _128_
timestamp 1698175906
transform 1 0 12544 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _129_
timestamp 1698175906
transform -1 0 13160 0 1 11760
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _130_
timestamp 1698175906
transform 1 0 11760 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _131_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9576 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _132_
timestamp 1698175906
transform 1 0 10024 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _133_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9184 0 1 8624
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _134_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 7784 0 -1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _135_
timestamp 1698175906
transform 1 0 6776 0 1 7840
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _136_
timestamp 1698175906
transform -1 0 7224 0 -1 10976
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _137_
timestamp 1698175906
transform -1 0 8288 0 -1 10192
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _138_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8400 0 1 7840
box -43 -43 1779 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _139_
timestamp 1698175906
transform 1 0 6888 0 1 9408
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _140_
timestamp 1698175906
transform 1 0 8624 0 -1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _141_
timestamp 1698175906
transform 1 0 8568 0 1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _142_
timestamp 1698175906
transform 1 0 11256 0 1 11760
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _143_
timestamp 1698175906
transform 1 0 9352 0 -1 7840
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _144_
timestamp 1698175906
transform 1 0 13048 0 -1 10976
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _145_
timestamp 1698175906
transform 1 0 13160 0 -1 9408
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _146_
timestamp 1698175906
transform 1 0 10696 0 1 7840
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _147_
timestamp 1698175906
transform 1 0 12768 0 1 10976
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _148_
timestamp 1698175906
transform -1 0 7560 0 -1 8624
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _149_
timestamp 1698175906
transform -1 0 8288 0 1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _150_
timestamp 1698175906
transform 1 0 10864 0 1 12544
box -43 -43 1779 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _151_
timestamp 1698175906
transform 1 0 11760 0 1 8624
box -43 -43 1779 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _152_
timestamp 1698175906
transform 1 0 10808 0 -1 10976
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _153_
timestamp 1698175906
transform -1 0 7336 0 -1 9408
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _155_
timestamp 1698175906
transform 1 0 14504 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _156_
timestamp 1698175906
transform -1 0 12936 0 1 12544
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _157_
timestamp 1698175906
transform 1 0 14504 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _158_
timestamp 1698175906
transform 1 0 11648 0 -1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _159_
timestamp 1698175906
transform 1 0 12824 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _160_
timestamp 1698175906
transform 1 0 12824 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _161_
timestamp 1698175906
transform 1 0 15120 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _162_
timestamp 1698175906
transform 1 0 14672 0 -1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _163_
timestamp 1698175906
transform 1 0 11984 0 -1 13328
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 9352 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9632 0 -1 10192
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1698175906
transform -1 0 10472 0 1 10192
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1698175906
transform 1 0 11592 0 1 10192
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout26 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 15120 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 784 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698175906
transform 1 0 2688 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698175906
transform 1 0 4592 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698175906
transform 1 0 6496 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_138 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8400 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_142 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8624 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_172
timestamp 1698175906
transform 1 0 10304 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_174 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10416 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_201
timestamp 1698175906
transform 1 0 11928 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_203
timestamp 1698175906
transform 1 0 12040 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_232
timestamp 1698175906
transform 1 0 13664 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_236
timestamp 1698175906
transform 1 0 13888 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_240
timestamp 1698175906
transform 1 0 14112 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_274
timestamp 1698175906
transform 1 0 16016 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_308
timestamp 1698175906
transform 1 0 17920 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_342
timestamp 1698175906
transform 1 0 19824 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_346
timestamp 1698175906
transform 1 0 20048 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_348
timestamp 1698175906
transform 1 0 20160 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 784 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698175906
transform 1 0 4368 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698175906
transform 1 0 4704 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698175906
transform 1 0 8288 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_142
timestamp 1698175906
transform 1 0 8624 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_206
timestamp 1698175906
transform 1 0 12208 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_212
timestamp 1698175906
transform 1 0 12544 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_276
timestamp 1698175906
transform 1 0 16128 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_282
timestamp 1698175906
transform 1 0 16464 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_346
timestamp 1698175906
transform 1 0 20048 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_348
timestamp 1698175906
transform 1 0 20160 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698175906
transform 1 0 784 0 1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698175906
transform 1 0 2576 0 1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698175906
transform 1 0 2744 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698175906
transform 1 0 6328 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_107
timestamp 1698175906
transform 1 0 6664 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_171
timestamp 1698175906
transform 1 0 10248 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_177 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10584 0 1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_193
timestamp 1698175906
transform 1 0 11480 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_197
timestamp 1698175906
transform 1 0 11704 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_225
timestamp 1698175906
transform 1 0 13272 0 1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_241
timestamp 1698175906
transform 1 0 14168 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698175906
transform 1 0 14504 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698175906
transform 1 0 18088 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_317
timestamp 1698175906
transform 1 0 18424 0 1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698175906
transform 1 0 784 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698175906
transform 1 0 4368 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698175906
transform 1 0 4704 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698175906
transform 1 0 8288 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_142
timestamp 1698175906
transform 1 0 8624 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_206
timestamp 1698175906
transform 1 0 12208 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_212
timestamp 1698175906
transform 1 0 12544 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_276
timestamp 1698175906
transform 1 0 16128 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_282
timestamp 1698175906
transform 1 0 16464 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_346
timestamp 1698175906
transform 1 0 20048 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_348
timestamp 1698175906
transform 1 0 20160 0 -1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698175906
transform 1 0 784 0 1 3136
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698175906
transform 1 0 2576 0 1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698175906
transform 1 0 2744 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698175906
transform 1 0 6328 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_107
timestamp 1698175906
transform 1 0 6664 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698175906
transform 1 0 10248 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_177
timestamp 1698175906
transform 1 0 10584 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_241
timestamp 1698175906
transform 1 0 14168 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698175906
transform 1 0 14504 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698175906
transform 1 0 18088 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_317
timestamp 1698175906
transform 1 0 18424 0 1 3136
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698175906
transform 1 0 784 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698175906
transform 1 0 4368 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698175906
transform 1 0 4704 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698175906
transform 1 0 8288 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_142
timestamp 1698175906
transform 1 0 8624 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_206
timestamp 1698175906
transform 1 0 12208 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_212
timestamp 1698175906
transform 1 0 12544 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698175906
transform 1 0 16128 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_282
timestamp 1698175906
transform 1 0 16464 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_346
timestamp 1698175906
transform 1 0 20048 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_348
timestamp 1698175906
transform 1 0 20160 0 -1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698175906
transform 1 0 784 0 1 3920
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698175906
transform 1 0 2576 0 1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698175906
transform 1 0 2744 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698175906
transform 1 0 6328 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_107
timestamp 1698175906
transform 1 0 6664 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_171
timestamp 1698175906
transform 1 0 10248 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_177
timestamp 1698175906
transform 1 0 10584 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_241
timestamp 1698175906
transform 1 0 14168 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_247
timestamp 1698175906
transform 1 0 14504 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_311
timestamp 1698175906
transform 1 0 18088 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_317
timestamp 1698175906
transform 1 0 18424 0 1 3920
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698175906
transform 1 0 784 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698175906
transform 1 0 4368 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_72
timestamp 1698175906
transform 1 0 4704 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698175906
transform 1 0 8288 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_142
timestamp 1698175906
transform 1 0 8624 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_206
timestamp 1698175906
transform 1 0 12208 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_212
timestamp 1698175906
transform 1 0 12544 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_276
timestamp 1698175906
transform 1 0 16128 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_282
timestamp 1698175906
transform 1 0 16464 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_346
timestamp 1698175906
transform 1 0 20048 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_348
timestamp 1698175906
transform 1 0 20160 0 -1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698175906
transform 1 0 784 0 1 4704
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698175906
transform 1 0 2576 0 1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_37
timestamp 1698175906
transform 1 0 2744 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_101
timestamp 1698175906
transform 1 0 6328 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_107
timestamp 1698175906
transform 1 0 6664 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_171
timestamp 1698175906
transform 1 0 10248 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_177
timestamp 1698175906
transform 1 0 10584 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_241
timestamp 1698175906
transform 1 0 14168 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_247
timestamp 1698175906
transform 1 0 14504 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_311
timestamp 1698175906
transform 1 0 18088 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_317
timestamp 1698175906
transform 1 0 18424 0 1 4704
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698175906
transform 1 0 784 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698175906
transform 1 0 4368 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_72
timestamp 1698175906
transform 1 0 4704 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_136
timestamp 1698175906
transform 1 0 8288 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_142
timestamp 1698175906
transform 1 0 8624 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_206
timestamp 1698175906
transform 1 0 12208 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_212
timestamp 1698175906
transform 1 0 12544 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_276
timestamp 1698175906
transform 1 0 16128 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_282
timestamp 1698175906
transform 1 0 16464 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_346
timestamp 1698175906
transform 1 0 20048 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_348
timestamp 1698175906
transform 1 0 20160 0 -1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698175906
transform 1 0 784 0 1 5488
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698175906
transform 1 0 2576 0 1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_37
timestamp 1698175906
transform 1 0 2744 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698175906
transform 1 0 6328 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_107
timestamp 1698175906
transform 1 0 6664 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_171
timestamp 1698175906
transform 1 0 10248 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_177
timestamp 1698175906
transform 1 0 10584 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_241
timestamp 1698175906
transform 1 0 14168 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_247
timestamp 1698175906
transform 1 0 14504 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_311
timestamp 1698175906
transform 1 0 18088 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_317
timestamp 1698175906
transform 1 0 18424 0 1 5488
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2
timestamp 1698175906
transform 1 0 784 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698175906
transform 1 0 4368 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_72
timestamp 1698175906
transform 1 0 4704 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698175906
transform 1 0 8288 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_142
timestamp 1698175906
transform 1 0 8624 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_206
timestamp 1698175906
transform 1 0 12208 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_212
timestamp 1698175906
transform 1 0 12544 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_276
timestamp 1698175906
transform 1 0 16128 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_282
timestamp 1698175906
transform 1 0 16464 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_346
timestamp 1698175906
transform 1 0 20048 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_348
timestamp 1698175906
transform 1 0 20160 0 -1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698175906
transform 1 0 784 0 1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698175906
transform 1 0 2576 0 1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_37
timestamp 1698175906
transform 1 0 2744 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698175906
transform 1 0 6328 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_107
timestamp 1698175906
transform 1 0 6664 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_171
timestamp 1698175906
transform 1 0 10248 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_177
timestamp 1698175906
transform 1 0 10584 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_241
timestamp 1698175906
transform 1 0 14168 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_247
timestamp 1698175906
transform 1 0 14504 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_311
timestamp 1698175906
transform 1 0 18088 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_317
timestamp 1698175906
transform 1 0 18424 0 1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_2
timestamp 1698175906
transform 1 0 784 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_66
timestamp 1698175906
transform 1 0 4368 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_72
timestamp 1698175906
transform 1 0 4704 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_136
timestamp 1698175906
transform 1 0 8288 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_142
timestamp 1698175906
transform 1 0 8624 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_206
timestamp 1698175906
transform 1 0 12208 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_212
timestamp 1698175906
transform 1 0 12544 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_276
timestamp 1698175906
transform 1 0 16128 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_282
timestamp 1698175906
transform 1 0 16464 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_346
timestamp 1698175906
transform 1 0 20048 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_348
timestamp 1698175906
transform 1 0 20160 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698175906
transform 1 0 784 0 1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698175906
transform 1 0 2576 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_37
timestamp 1698175906
transform 1 0 2744 0 1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_101
timestamp 1698175906
transform 1 0 6328 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_107
timestamp 1698175906
transform 1 0 6664 0 1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_171
timestamp 1698175906
transform 1 0 10248 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_177
timestamp 1698175906
transform 1 0 10584 0 1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_241
timestamp 1698175906
transform 1 0 14168 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_247
timestamp 1698175906
transform 1 0 14504 0 1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_311
timestamp 1698175906
transform 1 0 18088 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_317
timestamp 1698175906
transform 1 0 18424 0 1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_2
timestamp 1698175906
transform 1 0 784 0 -1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_66
timestamp 1698175906
transform 1 0 4368 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_72
timestamp 1698175906
transform 1 0 4704 0 -1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_136
timestamp 1698175906
transform 1 0 8288 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_142 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8624 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_150
timestamp 1698175906
transform 1 0 9072 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_154
timestamp 1698175906
transform 1 0 9296 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_184
timestamp 1698175906
transform 1 0 10976 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_192
timestamp 1698175906
transform 1 0 11424 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_202
timestamp 1698175906
transform 1 0 11984 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_212
timestamp 1698175906
transform 1 0 12544 0 -1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_276
timestamp 1698175906
transform 1 0 16128 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_282
timestamp 1698175906
transform 1 0 16464 0 -1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_314
timestamp 1698175906
transform 1 0 18256 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_322
timestamp 1698175906
transform 1 0 18704 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_2
timestamp 1698175906
transform 1 0 784 0 1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698175906
transform 1 0 2576 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_37
timestamp 1698175906
transform 1 0 2744 0 1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_101
timestamp 1698175906
transform 1 0 6328 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_107
timestamp 1698175906
transform 1 0 6664 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_169
timestamp 1698175906
transform 1 0 10136 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_173
timestamp 1698175906
transform 1 0 10360 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_177
timestamp 1698175906
transform 1 0 10584 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_208
timestamp 1698175906
transform 1 0 12320 0 1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_240
timestamp 1698175906
transform 1 0 14112 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_244
timestamp 1698175906
transform 1 0 14336 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_247
timestamp 1698175906
transform 1 0 14504 0 1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_311
timestamp 1698175906
transform 1 0 18088 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_317
timestamp 1698175906
transform 1 0 18424 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_321
timestamp 1698175906
transform 1 0 18648 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_2
timestamp 1698175906
transform 1 0 784 0 -1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_66
timestamp 1698175906
transform 1 0 4368 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_72
timestamp 1698175906
transform 1 0 4704 0 -1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_88
timestamp 1698175906
transform 1 0 5600 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_92
timestamp 1698175906
transform 1 0 5824 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_128
timestamp 1698175906
transform 1 0 7840 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_132
timestamp 1698175906
transform 1 0 8064 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_134
timestamp 1698175906
transform 1 0 8176 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_142
timestamp 1698175906
transform 1 0 8624 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_169
timestamp 1698175906
transform 1 0 10136 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_177
timestamp 1698175906
transform 1 0 10584 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_181
timestamp 1698175906
transform 1 0 10808 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_196
timestamp 1698175906
transform 1 0 11648 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_204
timestamp 1698175906
transform 1 0 12096 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_208
timestamp 1698175906
transform 1 0 12320 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_212
timestamp 1698175906
transform 1 0 12544 0 -1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_276
timestamp 1698175906
transform 1 0 16128 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_282
timestamp 1698175906
transform 1 0 16464 0 -1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_314
timestamp 1698175906
transform 1 0 18256 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_322
timestamp 1698175906
transform 1 0 18704 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_28
timestamp 1698175906
transform 1 0 2240 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_32
timestamp 1698175906
transform 1 0 2464 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698175906
transform 1 0 2576 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_37
timestamp 1698175906
transform 1 0 2744 0 1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_101
timestamp 1698175906
transform 1 0 6328 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_107
timestamp 1698175906
transform 1 0 6664 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_117
timestamp 1698175906
transform 1 0 7224 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_124
timestamp 1698175906
transform 1 0 7616 0 1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_140
timestamp 1698175906
transform 1 0 8512 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_149
timestamp 1698175906
transform 1 0 9016 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_151
timestamp 1698175906
transform 1 0 9128 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_183
timestamp 1698175906
transform 1 0 10920 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_191
timestamp 1698175906
transform 1 0 11368 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_195
timestamp 1698175906
transform 1 0 11592 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_197
timestamp 1698175906
transform 1 0 11704 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_229
timestamp 1698175906
transform 1 0 13496 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_237
timestamp 1698175906
transform 1 0 13944 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_242
timestamp 1698175906
transform 1 0 14224 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_244
timestamp 1698175906
transform 1 0 14336 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_253
timestamp 1698175906
transform 1 0 14840 0 1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_285
timestamp 1698175906
transform 1 0 16632 0 1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_301
timestamp 1698175906
transform 1 0 17528 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_309
timestamp 1698175906
transform 1 0 17976 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_313
timestamp 1698175906
transform 1 0 18200 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_317
timestamp 1698175906
transform 1 0 18424 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_321
timestamp 1698175906
transform 1 0 18648 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_28
timestamp 1698175906
transform 1 0 2240 0 -1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_60
timestamp 1698175906
transform 1 0 4032 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_68
timestamp 1698175906
transform 1 0 4480 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_72
timestamp 1698175906
transform 1 0 4704 0 -1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_88
timestamp 1698175906
transform 1 0 5600 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_132
timestamp 1698175906
transform 1 0 8064 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_142
timestamp 1698175906
transform 1 0 8624 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_146
timestamp 1698175906
transform 1 0 8848 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_154
timestamp 1698175906
transform 1 0 9296 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_156
timestamp 1698175906
transform 1 0 9408 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_200
timestamp 1698175906
transform 1 0 11872 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_208
timestamp 1698175906
transform 1 0 12320 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_212
timestamp 1698175906
transform 1 0 12544 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_216
timestamp 1698175906
transform 1 0 12768 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_264
timestamp 1698175906
transform 1 0 15456 0 -1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_282
timestamp 1698175906
transform 1 0 16464 0 -1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_314
timestamp 1698175906
transform 1 0 18256 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_322
timestamp 1698175906
transform 1 0 18704 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_2
timestamp 1698175906
transform 1 0 784 0 1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698175906
transform 1 0 2576 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_37
timestamp 1698175906
transform 1 0 2744 0 1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_101
timestamp 1698175906
transform 1 0 6328 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_107
timestamp 1698175906
transform 1 0 6664 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_140
timestamp 1698175906
transform 1 0 8512 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_148
timestamp 1698175906
transform 1 0 8960 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_152
timestamp 1698175906
transform 1 0 9184 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_173
timestamp 1698175906
transform 1 0 10360 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_177
timestamp 1698175906
transform 1 0 10584 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_179
timestamp 1698175906
transform 1 0 10696 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_194
timestamp 1698175906
transform 1 0 11536 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_198
timestamp 1698175906
transform 1 0 11760 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_216
timestamp 1698175906
transform 1 0 12768 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_223
timestamp 1698175906
transform 1 0 13160 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_227
timestamp 1698175906
transform 1 0 13384 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_236
timestamp 1698175906
transform 1 0 13888 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_244
timestamp 1698175906
transform 1 0 14336 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_253
timestamp 1698175906
transform 1 0 14840 0 1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_285
timestamp 1698175906
transform 1 0 16632 0 1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_301
timestamp 1698175906
transform 1 0 17528 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_309
timestamp 1698175906
transform 1 0 17976 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_313
timestamp 1698175906
transform 1 0 18200 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_317
timestamp 1698175906
transform 1 0 18424 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_321
timestamp 1698175906
transform 1 0 18648 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_2
timestamp 1698175906
transform 1 0 784 0 -1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_66
timestamp 1698175906
transform 1 0 4368 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_72
timestamp 1698175906
transform 1 0 4704 0 -1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_104
timestamp 1698175906
transform 1 0 6496 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_106
timestamp 1698175906
transform 1 0 6608 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_136
timestamp 1698175906
transform 1 0 8288 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_142
timestamp 1698175906
transform 1 0 8624 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_144
timestamp 1698175906
transform 1 0 8736 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_218
timestamp 1698175906
transform 1 0 12880 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_222
timestamp 1698175906
transform 1 0 13104 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_231
timestamp 1698175906
transform 1 0 13608 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_238
timestamp 1698175906
transform 1 0 14000 0 -1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_270
timestamp 1698175906
transform 1 0 15792 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_278
timestamp 1698175906
transform 1 0 16240 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_282
timestamp 1698175906
transform 1 0 16464 0 -1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_314
timestamp 1698175906
transform 1 0 18256 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_322
timestamp 1698175906
transform 1 0 18704 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_2
timestamp 1698175906
transform 1 0 784 0 1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698175906
transform 1 0 2576 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_37
timestamp 1698175906
transform 1 0 2744 0 1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_101
timestamp 1698175906
transform 1 0 6328 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_107
timestamp 1698175906
transform 1 0 6664 0 1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_123
timestamp 1698175906
transform 1 0 7560 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_181
timestamp 1698175906
transform 1 0 10808 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_183
timestamp 1698175906
transform 1 0 10920 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_193
timestamp 1698175906
transform 1 0 11480 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_247
timestamp 1698175906
transform 1 0 14504 0 1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_311
timestamp 1698175906
transform 1 0 18088 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_317
timestamp 1698175906
transform 1 0 18424 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_321
timestamp 1698175906
transform 1 0 18648 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_2
timestamp 1698175906
transform 1 0 784 0 -1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_66
timestamp 1698175906
transform 1 0 4368 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_72
timestamp 1698175906
transform 1 0 4704 0 -1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_117
timestamp 1698175906
transform 1 0 7224 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_119
timestamp 1698175906
transform 1 0 7336 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_128
timestamp 1698175906
transform 1 0 7840 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_136
timestamp 1698175906
transform 1 0 8288 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_154
timestamp 1698175906
transform 1 0 9296 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_158
timestamp 1698175906
transform 1 0 9520 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_212
timestamp 1698175906
transform 1 0 12544 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_220
timestamp 1698175906
transform 1 0 12992 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_256
timestamp 1698175906
transform 1 0 15008 0 -1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_272
timestamp 1698175906
transform 1 0 15904 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_282
timestamp 1698175906
transform 1 0 16464 0 -1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_314
timestamp 1698175906
transform 1 0 18256 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_322
timestamp 1698175906
transform 1 0 18704 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_28
timestamp 1698175906
transform 1 0 2240 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_32
timestamp 1698175906
transform 1 0 2464 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698175906
transform 1 0 2576 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_37
timestamp 1698175906
transform 1 0 2744 0 1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_101
timestamp 1698175906
transform 1 0 6328 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_107
timestamp 1698175906
transform 1 0 6664 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_125
timestamp 1698175906
transform 1 0 7672 0 1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_141
timestamp 1698175906
transform 1 0 8568 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_149
timestamp 1698175906
transform 1 0 9016 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_153
timestamp 1698175906
transform 1 0 9240 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_168
timestamp 1698175906
transform 1 0 10080 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_172
timestamp 1698175906
transform 1 0 10304 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_174
timestamp 1698175906
transform 1 0 10416 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_187
timestamp 1698175906
transform 1 0 11144 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_191
timestamp 1698175906
transform 1 0 11368 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_203
timestamp 1698175906
transform 1 0 12040 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_211
timestamp 1698175906
transform 1 0 12488 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_215
timestamp 1698175906
transform 1 0 12712 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_247
timestamp 1698175906
transform 1 0 14504 0 1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_311
timestamp 1698175906
transform 1 0 18088 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_317
timestamp 1698175906
transform 1 0 18424 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_321
timestamp 1698175906
transform 1 0 18648 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_28
timestamp 1698175906
transform 1 0 2240 0 -1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_60
timestamp 1698175906
transform 1 0 4032 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_68
timestamp 1698175906
transform 1 0 4480 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_72
timestamp 1698175906
transform 1 0 4704 0 -1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_104
timestamp 1698175906
transform 1 0 6496 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_112
timestamp 1698175906
transform 1 0 6944 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_114
timestamp 1698175906
transform 1 0 7056 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_129
timestamp 1698175906
transform 1 0 7896 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_137
timestamp 1698175906
transform 1 0 8344 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_139
timestamp 1698175906
transform 1 0 8456 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_142
timestamp 1698175906
transform 1 0 8624 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_150
timestamp 1698175906
transform 1 0 9072 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_152
timestamp 1698175906
transform 1 0 9184 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_181
timestamp 1698175906
transform 1 0 10808 0 -1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_197
timestamp 1698175906
transform 1 0 11704 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_205
timestamp 1698175906
transform 1 0 12152 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_209
timestamp 1698175906
transform 1 0 12376 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_212
timestamp 1698175906
transform 1 0 12544 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_220
timestamp 1698175906
transform 1 0 12992 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_224
timestamp 1698175906
transform 1 0 13216 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_231
timestamp 1698175906
transform 1 0 13608 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_237
timestamp 1698175906
transform 1 0 13944 0 -1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_269
timestamp 1698175906
transform 1 0 15736 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_277
timestamp 1698175906
transform 1 0 16184 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_279
timestamp 1698175906
transform 1 0 16296 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_282
timestamp 1698175906
transform 1 0 16464 0 -1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_314
timestamp 1698175906
transform 1 0 18256 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_322
timestamp 1698175906
transform 1 0 18704 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_2
timestamp 1698175906
transform 1 0 784 0 1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698175906
transform 1 0 2576 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_37
timestamp 1698175906
transform 1 0 2744 0 1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_101
timestamp 1698175906
transform 1 0 6328 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_107
timestamp 1698175906
transform 1 0 6664 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_115
timestamp 1698175906
transform 1 0 7112 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_132
timestamp 1698175906
transform 1 0 8064 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_140
timestamp 1698175906
transform 1 0 8512 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_156
timestamp 1698175906
transform 1 0 9408 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_160
timestamp 1698175906
transform 1 0 9632 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_177
timestamp 1698175906
transform 1 0 10584 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_185
timestamp 1698175906
transform 1 0 11032 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_223
timestamp 1698175906
transform 1 0 13160 0 1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_239
timestamp 1698175906
transform 1 0 14056 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_243
timestamp 1698175906
transform 1 0 14280 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_247
timestamp 1698175906
transform 1 0 14504 0 1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_311
timestamp 1698175906
transform 1 0 18088 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_317
timestamp 1698175906
transform 1 0 18424 0 1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_28
timestamp 1698175906
transform 1 0 2240 0 -1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_60
timestamp 1698175906
transform 1 0 4032 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_68
timestamp 1698175906
transform 1 0 4480 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_72
timestamp 1698175906
transform 1 0 4704 0 -1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_88
timestamp 1698175906
transform 1 0 5600 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_96
timestamp 1698175906
transform 1 0 6048 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_179
timestamp 1698175906
transform 1 0 10696 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_183
timestamp 1698175906
transform 1 0 10920 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_206
timestamp 1698175906
transform 1 0 12208 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_212
timestamp 1698175906
transform 1 0 12544 0 -1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_276
timestamp 1698175906
transform 1 0 16128 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_282
timestamp 1698175906
transform 1 0 16464 0 -1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_314
timestamp 1698175906
transform 1 0 18256 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_322
timestamp 1698175906
transform 1 0 18704 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_28
timestamp 1698175906
transform 1 0 2240 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_32
timestamp 1698175906
transform 1 0 2464 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698175906
transform 1 0 2576 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_37
timestamp 1698175906
transform 1 0 2744 0 1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_101
timestamp 1698175906
transform 1 0 6328 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_136
timestamp 1698175906
transform 1 0 8288 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_140
timestamp 1698175906
transform 1 0 8512 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_170
timestamp 1698175906
transform 1 0 10192 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_174
timestamp 1698175906
transform 1 0 10416 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_177
timestamp 1698175906
transform 1 0 10584 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_181
timestamp 1698175906
transform 1 0 10808 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_219
timestamp 1698175906
transform 1 0 12936 0 1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_235
timestamp 1698175906
transform 1 0 13832 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_243
timestamp 1698175906
transform 1 0 14280 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_247
timestamp 1698175906
transform 1 0 14504 0 1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_311
timestamp 1698175906
transform 1 0 18088 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_317
timestamp 1698175906
transform 1 0 18424 0 1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_2
timestamp 1698175906
transform 1 0 784 0 -1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_66
timestamp 1698175906
transform 1 0 4368 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_72
timestamp 1698175906
transform 1 0 4704 0 -1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_104
timestamp 1698175906
transform 1 0 6496 0 -1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_120
timestamp 1698175906
transform 1 0 7392 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_126
timestamp 1698175906
transform 1 0 7728 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_134
timestamp 1698175906
transform 1 0 8176 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_138
timestamp 1698175906
transform 1 0 8400 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_142
timestamp 1698175906
transform 1 0 8624 0 -1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_174
timestamp 1698175906
transform 1 0 10416 0 -1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_190
timestamp 1698175906
transform 1 0 11312 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_198
timestamp 1698175906
transform 1 0 11760 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_208
timestamp 1698175906
transform 1 0 12320 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_212
timestamp 1698175906
transform 1 0 12544 0 -1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_276
timestamp 1698175906
transform 1 0 16128 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_282
timestamp 1698175906
transform 1 0 16464 0 -1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_346
timestamp 1698175906
transform 1 0 20048 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_348
timestamp 1698175906
transform 1 0 20160 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_2
timestamp 1698175906
transform 1 0 784 0 1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698175906
transform 1 0 2576 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_37
timestamp 1698175906
transform 1 0 2744 0 1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_101
timestamp 1698175906
transform 1 0 6328 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_107
timestamp 1698175906
transform 1 0 6664 0 1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_171
timestamp 1698175906
transform 1 0 10248 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_177
timestamp 1698175906
transform 1 0 10584 0 1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_241
timestamp 1698175906
transform 1 0 14168 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_247
timestamp 1698175906
transform 1 0 14504 0 1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_311
timestamp 1698175906
transform 1 0 18088 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_317
timestamp 1698175906
transform 1 0 18424 0 1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_2
timestamp 1698175906
transform 1 0 784 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_66
timestamp 1698175906
transform 1 0 4368 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_72
timestamp 1698175906
transform 1 0 4704 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_136
timestamp 1698175906
transform 1 0 8288 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_142
timestamp 1698175906
transform 1 0 8624 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_206
timestamp 1698175906
transform 1 0 12208 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_212
timestamp 1698175906
transform 1 0 12544 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_276
timestamp 1698175906
transform 1 0 16128 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_282
timestamp 1698175906
transform 1 0 16464 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_346
timestamp 1698175906
transform 1 0 20048 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_348
timestamp 1698175906
transform 1 0 20160 0 -1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_2
timestamp 1698175906
transform 1 0 784 0 1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698175906
transform 1 0 2576 0 1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_37
timestamp 1698175906
transform 1 0 2744 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_101
timestamp 1698175906
transform 1 0 6328 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_107
timestamp 1698175906
transform 1 0 6664 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_171
timestamp 1698175906
transform 1 0 10248 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_177
timestamp 1698175906
transform 1 0 10584 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_241
timestamp 1698175906
transform 1 0 14168 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_247
timestamp 1698175906
transform 1 0 14504 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_311
timestamp 1698175906
transform 1 0 18088 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_317
timestamp 1698175906
transform 1 0 18424 0 1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_2
timestamp 1698175906
transform 1 0 784 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_66
timestamp 1698175906
transform 1 0 4368 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_72
timestamp 1698175906
transform 1 0 4704 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_136
timestamp 1698175906
transform 1 0 8288 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_142
timestamp 1698175906
transform 1 0 8624 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_206
timestamp 1698175906
transform 1 0 12208 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_212
timestamp 1698175906
transform 1 0 12544 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_276
timestamp 1698175906
transform 1 0 16128 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_282
timestamp 1698175906
transform 1 0 16464 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_346
timestamp 1698175906
transform 1 0 20048 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_348
timestamp 1698175906
transform 1 0 20160 0 -1 14896
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698175906
transform 1 0 784 0 1 14896
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698175906
transform 1 0 2576 0 1 14896
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_37
timestamp 1698175906
transform 1 0 2744 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_101
timestamp 1698175906
transform 1 0 6328 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_107
timestamp 1698175906
transform 1 0 6664 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_171
timestamp 1698175906
transform 1 0 10248 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_177
timestamp 1698175906
transform 1 0 10584 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_241
timestamp 1698175906
transform 1 0 14168 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_247
timestamp 1698175906
transform 1 0 14504 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_311
timestamp 1698175906
transform 1 0 18088 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_317
timestamp 1698175906
transform 1 0 18424 0 1 14896
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2
timestamp 1698175906
transform 1 0 784 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_66
timestamp 1698175906
transform 1 0 4368 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_72
timestamp 1698175906
transform 1 0 4704 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_136
timestamp 1698175906
transform 1 0 8288 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_142
timestamp 1698175906
transform 1 0 8624 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_206
timestamp 1698175906
transform 1 0 12208 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_212
timestamp 1698175906
transform 1 0 12544 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_276
timestamp 1698175906
transform 1 0 16128 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_282
timestamp 1698175906
transform 1 0 16464 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_346
timestamp 1698175906
transform 1 0 20048 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_348
timestamp 1698175906
transform 1 0 20160 0 -1 15680
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_2
timestamp 1698175906
transform 1 0 784 0 1 15680
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698175906
transform 1 0 2576 0 1 15680
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_37
timestamp 1698175906
transform 1 0 2744 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_101
timestamp 1698175906
transform 1 0 6328 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_107
timestamp 1698175906
transform 1 0 6664 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_171
timestamp 1698175906
transform 1 0 10248 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_177
timestamp 1698175906
transform 1 0 10584 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_241
timestamp 1698175906
transform 1 0 14168 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_247
timestamp 1698175906
transform 1 0 14504 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_311
timestamp 1698175906
transform 1 0 18088 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_317
timestamp 1698175906
transform 1 0 18424 0 1 15680
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2
timestamp 1698175906
transform 1 0 784 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_66
timestamp 1698175906
transform 1 0 4368 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_72
timestamp 1698175906
transform 1 0 4704 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_136
timestamp 1698175906
transform 1 0 8288 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_142
timestamp 1698175906
transform 1 0 8624 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_206
timestamp 1698175906
transform 1 0 12208 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_212
timestamp 1698175906
transform 1 0 12544 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_276
timestamp 1698175906
transform 1 0 16128 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_282
timestamp 1698175906
transform 1 0 16464 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_346
timestamp 1698175906
transform 1 0 20048 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_348
timestamp 1698175906
transform 1 0 20160 0 -1 16464
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698175906
transform 1 0 784 0 1 16464
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698175906
transform 1 0 2576 0 1 16464
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_37
timestamp 1698175906
transform 1 0 2744 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_101
timestamp 1698175906
transform 1 0 6328 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_107
timestamp 1698175906
transform 1 0 6664 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_171
timestamp 1698175906
transform 1 0 10248 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_177
timestamp 1698175906
transform 1 0 10584 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_241
timestamp 1698175906
transform 1 0 14168 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_247
timestamp 1698175906
transform 1 0 14504 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_311
timestamp 1698175906
transform 1 0 18088 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_317
timestamp 1698175906
transform 1 0 18424 0 1 16464
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_2
timestamp 1698175906
transform 1 0 784 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_66
timestamp 1698175906
transform 1 0 4368 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_72
timestamp 1698175906
transform 1 0 4704 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_136
timestamp 1698175906
transform 1 0 8288 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_142
timestamp 1698175906
transform 1 0 8624 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_206
timestamp 1698175906
transform 1 0 12208 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_212
timestamp 1698175906
transform 1 0 12544 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_276
timestamp 1698175906
transform 1 0 16128 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_282
timestamp 1698175906
transform 1 0 16464 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_346
timestamp 1698175906
transform 1 0 20048 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_348
timestamp 1698175906
transform 1 0 20160 0 -1 17248
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698175906
transform 1 0 784 0 1 17248
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698175906
transform 1 0 2576 0 1 17248
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_37
timestamp 1698175906
transform 1 0 2744 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_101
timestamp 1698175906
transform 1 0 6328 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_107
timestamp 1698175906
transform 1 0 6664 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_171
timestamp 1698175906
transform 1 0 10248 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_177
timestamp 1698175906
transform 1 0 10584 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_241
timestamp 1698175906
transform 1 0 14168 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_247
timestamp 1698175906
transform 1 0 14504 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_311
timestamp 1698175906
transform 1 0 18088 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_317
timestamp 1698175906
transform 1 0 18424 0 1 17248
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2
timestamp 1698175906
transform 1 0 784 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1698175906
transform 1 0 4368 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_72
timestamp 1698175906
transform 1 0 4704 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_136
timestamp 1698175906
transform 1 0 8288 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_142
timestamp 1698175906
transform 1 0 8624 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_206
timestamp 1698175906
transform 1 0 12208 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_212
timestamp 1698175906
transform 1 0 12544 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_276
timestamp 1698175906
transform 1 0 16128 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_282
timestamp 1698175906
transform 1 0 16464 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_346
timestamp 1698175906
transform 1 0 20048 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_348
timestamp 1698175906
transform 1 0 20160 0 -1 18032
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_2
timestamp 1698175906
transform 1 0 784 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698175906
transform 1 0 2576 0 1 18032
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_37
timestamp 1698175906
transform 1 0 2744 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_101
timestamp 1698175906
transform 1 0 6328 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_107
timestamp 1698175906
transform 1 0 6664 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_171
timestamp 1698175906
transform 1 0 10248 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_177
timestamp 1698175906
transform 1 0 10584 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_209
timestamp 1698175906
transform 1 0 12376 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_237
timestamp 1698175906
transform 1 0 13944 0 1 18032
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_247
timestamp 1698175906
transform 1 0 14504 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_311
timestamp 1698175906
transform 1 0 18088 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_317
timestamp 1698175906
transform 1 0 18424 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_2
timestamp 1698175906
transform 1 0 784 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_66
timestamp 1698175906
transform 1 0 4368 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_72
timestamp 1698175906
transform 1 0 4704 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_136
timestamp 1698175906
transform 1 0 8288 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_142
timestamp 1698175906
transform 1 0 8624 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_206
timestamp 1698175906
transform 1 0 12208 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_238
timestamp 1698175906
transform 1 0 14000 0 -1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_270
timestamp 1698175906
transform 1 0 15792 0 -1 18816
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_278
timestamp 1698175906
transform 1 0 16240 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_282
timestamp 1698175906
transform 1 0 16464 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_346
timestamp 1698175906
transform 1 0 20048 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_348
timestamp 1698175906
transform 1 0 20160 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_2
timestamp 1698175906
transform 1 0 784 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_36
timestamp 1698175906
transform 1 0 2688 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_70
timestamp 1698175906
transform 1 0 4592 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_104
timestamp 1698175906
transform 1 0 6496 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_138
timestamp 1698175906
transform 1 0 8400 0 1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_143
timestamp 1698175906
transform 1 0 8680 0 1 18816
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_159
timestamp 1698175906
transform 1 0 9576 0 1 18816
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_167
timestamp 1698175906
transform 1 0 10024 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_169
timestamp 1698175906
transform 1 0 10136 0 1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_172
timestamp 1698175906
transform 1 0 10304 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_232
timestamp 1698175906
transform 1 0 13664 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_236
timestamp 1698175906
transform 1 0 13888 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_240
timestamp 1698175906
transform 1 0 14112 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_274
timestamp 1698175906
transform 1 0 16016 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_308
timestamp 1698175906
transform 1 0 17920 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_342
timestamp 1698175906
transform 1 0 19824 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_346
timestamp 1698175906
transform 1 0 20048 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_348
timestamp 1698175906
transform 1 0 20160 0 1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita29_27 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 8680 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18760 0 -1 7840
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output2
timestamp 1698175906
transform 1 0 18760 0 1 10192
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output3
timestamp 1698175906
transform 1 0 18760 0 -1 10192
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output4
timestamp 1698175906
transform 1 0 18760 0 -1 11760
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output5
timestamp 1698175906
transform 1 0 18760 0 -1 8624
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output6
timestamp 1698175906
transform 1 0 18760 0 -1 10976
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output7
timestamp 1698175906
transform 1 0 12488 0 1 18032
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output8
timestamp 1698175906
transform 1 0 18760 0 1 8624
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output9
timestamp 1698175906
transform 1 0 12208 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output10
timestamp 1698175906
transform 1 0 11816 0 1 2352
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output11
timestamp 1698175906
transform 1 0 12208 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output12
timestamp 1698175906
transform 1 0 18760 0 1 9408
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output13
timestamp 1698175906
transform 1 0 18760 0 -1 9408
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output14
timestamp 1698175906
transform 1 0 18760 0 1 7840
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output15
timestamp 1698175906
transform -1 0 2240 0 1 8624
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output16
timestamp 1698175906
transform -1 0 2240 0 1 12544
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output17
timestamp 1698175906
transform 1 0 18760 0 1 10976
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output18
timestamp 1698175906
transform 1 0 10472 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output19
timestamp 1698175906
transform 1 0 18760 0 -1 12544
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output20
timestamp 1698175906
transform 1 0 12544 0 -1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output21
timestamp 1698175906
transform -1 0 2240 0 1 10976
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output22
timestamp 1698175906
transform -1 0 2240 0 -1 11760
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output23
timestamp 1698175906
transform -1 0 2240 0 -1 12544
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output24
timestamp 1698175906
transform 1 0 8736 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output25
timestamp 1698175906
transform -1 0 2240 0 -1 9408
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_45 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 672 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698175906
transform -1 0 20328 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_46
timestamp 1698175906
transform 1 0 672 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698175906
transform -1 0 20328 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_47
timestamp 1698175906
transform 1 0 672 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698175906
transform -1 0 20328 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_48
timestamp 1698175906
transform 1 0 672 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698175906
transform -1 0 20328 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_49
timestamp 1698175906
transform 1 0 672 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698175906
transform -1 0 20328 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_50
timestamp 1698175906
transform 1 0 672 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698175906
transform -1 0 20328 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_51
timestamp 1698175906
transform 1 0 672 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698175906
transform -1 0 20328 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_52
timestamp 1698175906
transform 1 0 672 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698175906
transform -1 0 20328 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_53
timestamp 1698175906
transform 1 0 672 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698175906
transform -1 0 20328 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_54
timestamp 1698175906
transform 1 0 672 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698175906
transform -1 0 20328 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_55
timestamp 1698175906
transform 1 0 672 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698175906
transform -1 0 20328 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_56
timestamp 1698175906
transform 1 0 672 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698175906
transform -1 0 20328 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_57
timestamp 1698175906
transform 1 0 672 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698175906
transform -1 0 20328 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_58
timestamp 1698175906
transform 1 0 672 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698175906
transform -1 0 20328 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_59
timestamp 1698175906
transform 1 0 672 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698175906
transform -1 0 20328 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_60
timestamp 1698175906
transform 1 0 672 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698175906
transform -1 0 20328 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_61
timestamp 1698175906
transform 1 0 672 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698175906
transform -1 0 20328 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_62
timestamp 1698175906
transform 1 0 672 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698175906
transform -1 0 20328 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_63
timestamp 1698175906
transform 1 0 672 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698175906
transform -1 0 20328 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_64
timestamp 1698175906
transform 1 0 672 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698175906
transform -1 0 20328 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_65
timestamp 1698175906
transform 1 0 672 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698175906
transform -1 0 20328 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_66
timestamp 1698175906
transform 1 0 672 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698175906
transform -1 0 20328 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_67
timestamp 1698175906
transform 1 0 672 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698175906
transform -1 0 20328 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_68
timestamp 1698175906
transform 1 0 672 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698175906
transform -1 0 20328 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_69
timestamp 1698175906
transform 1 0 672 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698175906
transform -1 0 20328 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_70
timestamp 1698175906
transform 1 0 672 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698175906
transform -1 0 20328 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_71
timestamp 1698175906
transform 1 0 672 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698175906
transform -1 0 20328 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_72
timestamp 1698175906
transform 1 0 672 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698175906
transform -1 0 20328 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_73
timestamp 1698175906
transform 1 0 672 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698175906
transform -1 0 20328 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_74
timestamp 1698175906
transform 1 0 672 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698175906
transform -1 0 20328 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_75
timestamp 1698175906
transform 1 0 672 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698175906
transform -1 0 20328 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_76
timestamp 1698175906
transform 1 0 672 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698175906
transform -1 0 20328 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_77
timestamp 1698175906
transform 1 0 672 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698175906
transform -1 0 20328 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_78
timestamp 1698175906
transform 1 0 672 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698175906
transform -1 0 20328 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_79
timestamp 1698175906
transform 1 0 672 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698175906
transform -1 0 20328 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_80
timestamp 1698175906
transform 1 0 672 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698175906
transform -1 0 20328 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_81
timestamp 1698175906
transform 1 0 672 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698175906
transform -1 0 20328 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_82
timestamp 1698175906
transform 1 0 672 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698175906
transform -1 0 20328 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_83
timestamp 1698175906
transform 1 0 672 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698175906
transform -1 0 20328 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_84
timestamp 1698175906
transform 1 0 672 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698175906
transform -1 0 20328 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_85
timestamp 1698175906
transform 1 0 672 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698175906
transform -1 0 20328 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_86
timestamp 1698175906
transform 1 0 672 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698175906
transform -1 0 20328 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_87
timestamp 1698175906
transform 1 0 672 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698175906
transform -1 0 20328 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_88
timestamp 1698175906
transform 1 0 672 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698175906
transform -1 0 20328 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_89
timestamp 1698175906
transform 1 0 672 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698175906
transform -1 0 20328 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_90 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 2576 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_91
timestamp 1698175906
transform 1 0 4480 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_92
timestamp 1698175906
transform 1 0 6384 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_93
timestamp 1698175906
transform 1 0 8288 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_94
timestamp 1698175906
transform 1 0 10192 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_95
timestamp 1698175906
transform 1 0 12096 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_96
timestamp 1698175906
transform 1 0 14000 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_97
timestamp 1698175906
transform 1 0 15904 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_98
timestamp 1698175906
transform 1 0 17808 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_99
timestamp 1698175906
transform 1 0 19712 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_100
timestamp 1698175906
transform 1 0 4592 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_101
timestamp 1698175906
transform 1 0 8512 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_102
timestamp 1698175906
transform 1 0 12432 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_103
timestamp 1698175906
transform 1 0 16352 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_104
timestamp 1698175906
transform 1 0 2632 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_105
timestamp 1698175906
transform 1 0 6552 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_106
timestamp 1698175906
transform 1 0 10472 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_107
timestamp 1698175906
transform 1 0 14392 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_108
timestamp 1698175906
transform 1 0 18312 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_109
timestamp 1698175906
transform 1 0 4592 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_110
timestamp 1698175906
transform 1 0 8512 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_111
timestamp 1698175906
transform 1 0 12432 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_112
timestamp 1698175906
transform 1 0 16352 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_113
timestamp 1698175906
transform 1 0 2632 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_114
timestamp 1698175906
transform 1 0 6552 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_115
timestamp 1698175906
transform 1 0 10472 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_116
timestamp 1698175906
transform 1 0 14392 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_117
timestamp 1698175906
transform 1 0 18312 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_118
timestamp 1698175906
transform 1 0 4592 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_119
timestamp 1698175906
transform 1 0 8512 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_120
timestamp 1698175906
transform 1 0 12432 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_121
timestamp 1698175906
transform 1 0 16352 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_122
timestamp 1698175906
transform 1 0 2632 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_123
timestamp 1698175906
transform 1 0 6552 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_124
timestamp 1698175906
transform 1 0 10472 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_125
timestamp 1698175906
transform 1 0 14392 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_126
timestamp 1698175906
transform 1 0 18312 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_127
timestamp 1698175906
transform 1 0 4592 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_128
timestamp 1698175906
transform 1 0 8512 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_129
timestamp 1698175906
transform 1 0 12432 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_130
timestamp 1698175906
transform 1 0 16352 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_131
timestamp 1698175906
transform 1 0 2632 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_132
timestamp 1698175906
transform 1 0 6552 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_133
timestamp 1698175906
transform 1 0 10472 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_134
timestamp 1698175906
transform 1 0 14392 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_135
timestamp 1698175906
transform 1 0 18312 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_136
timestamp 1698175906
transform 1 0 4592 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_137
timestamp 1698175906
transform 1 0 8512 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_138
timestamp 1698175906
transform 1 0 12432 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_139
timestamp 1698175906
transform 1 0 16352 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_140
timestamp 1698175906
transform 1 0 2632 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_141
timestamp 1698175906
transform 1 0 6552 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_142
timestamp 1698175906
transform 1 0 10472 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_143
timestamp 1698175906
transform 1 0 14392 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_144
timestamp 1698175906
transform 1 0 18312 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_145
timestamp 1698175906
transform 1 0 4592 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_146
timestamp 1698175906
transform 1 0 8512 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_147
timestamp 1698175906
transform 1 0 12432 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_148
timestamp 1698175906
transform 1 0 16352 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_149
timestamp 1698175906
transform 1 0 2632 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_150
timestamp 1698175906
transform 1 0 6552 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_151
timestamp 1698175906
transform 1 0 10472 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_152
timestamp 1698175906
transform 1 0 14392 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_153
timestamp 1698175906
transform 1 0 18312 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_154
timestamp 1698175906
transform 1 0 4592 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_155
timestamp 1698175906
transform 1 0 8512 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_156
timestamp 1698175906
transform 1 0 12432 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_157
timestamp 1698175906
transform 1 0 16352 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_158
timestamp 1698175906
transform 1 0 2632 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_159
timestamp 1698175906
transform 1 0 6552 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_160
timestamp 1698175906
transform 1 0 10472 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_161
timestamp 1698175906
transform 1 0 14392 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_162
timestamp 1698175906
transform 1 0 18312 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_163
timestamp 1698175906
transform 1 0 4592 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_164
timestamp 1698175906
transform 1 0 8512 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_165
timestamp 1698175906
transform 1 0 12432 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_166
timestamp 1698175906
transform 1 0 16352 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_167
timestamp 1698175906
transform 1 0 2632 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_168
timestamp 1698175906
transform 1 0 6552 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_169
timestamp 1698175906
transform 1 0 10472 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_170
timestamp 1698175906
transform 1 0 14392 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_171
timestamp 1698175906
transform 1 0 18312 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_172
timestamp 1698175906
transform 1 0 4592 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_173
timestamp 1698175906
transform 1 0 8512 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_174
timestamp 1698175906
transform 1 0 12432 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_175
timestamp 1698175906
transform 1 0 16352 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_176
timestamp 1698175906
transform 1 0 2632 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_177
timestamp 1698175906
transform 1 0 6552 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_178
timestamp 1698175906
transform 1 0 10472 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_179
timestamp 1698175906
transform 1 0 14392 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_180
timestamp 1698175906
transform 1 0 18312 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_181
timestamp 1698175906
transform 1 0 4592 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_182
timestamp 1698175906
transform 1 0 8512 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_183
timestamp 1698175906
transform 1 0 12432 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_184
timestamp 1698175906
transform 1 0 16352 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_185
timestamp 1698175906
transform 1 0 2632 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_186
timestamp 1698175906
transform 1 0 6552 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_187
timestamp 1698175906
transform 1 0 10472 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_188
timestamp 1698175906
transform 1 0 14392 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_189
timestamp 1698175906
transform 1 0 18312 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_190
timestamp 1698175906
transform 1 0 4592 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_191
timestamp 1698175906
transform 1 0 8512 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_192
timestamp 1698175906
transform 1 0 12432 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_193
timestamp 1698175906
transform 1 0 16352 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_194
timestamp 1698175906
transform 1 0 2632 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_195
timestamp 1698175906
transform 1 0 6552 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_196
timestamp 1698175906
transform 1 0 10472 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_197
timestamp 1698175906
transform 1 0 14392 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_198
timestamp 1698175906
transform 1 0 18312 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_199
timestamp 1698175906
transform 1 0 4592 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_200
timestamp 1698175906
transform 1 0 8512 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_201
timestamp 1698175906
transform 1 0 12432 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_202
timestamp 1698175906
transform 1 0 16352 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_203
timestamp 1698175906
transform 1 0 2632 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_204
timestamp 1698175906
transform 1 0 6552 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_205
timestamp 1698175906
transform 1 0 10472 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_206
timestamp 1698175906
transform 1 0 14392 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_207
timestamp 1698175906
transform 1 0 18312 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_208
timestamp 1698175906
transform 1 0 4592 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_209
timestamp 1698175906
transform 1 0 8512 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_210
timestamp 1698175906
transform 1 0 12432 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_211
timestamp 1698175906
transform 1 0 16352 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_212
timestamp 1698175906
transform 1 0 2632 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_213
timestamp 1698175906
transform 1 0 6552 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_214
timestamp 1698175906
transform 1 0 10472 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_215
timestamp 1698175906
transform 1 0 14392 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_216
timestamp 1698175906
transform 1 0 18312 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_217
timestamp 1698175906
transform 1 0 4592 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_218
timestamp 1698175906
transform 1 0 8512 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_219
timestamp 1698175906
transform 1 0 12432 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_220
timestamp 1698175906
transform 1 0 16352 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_221
timestamp 1698175906
transform 1 0 2632 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_222
timestamp 1698175906
transform 1 0 6552 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_223
timestamp 1698175906
transform 1 0 10472 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_224
timestamp 1698175906
transform 1 0 14392 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_225
timestamp 1698175906
transform 1 0 18312 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_226
timestamp 1698175906
transform 1 0 4592 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_227
timestamp 1698175906
transform 1 0 8512 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_228
timestamp 1698175906
transform 1 0 12432 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_229
timestamp 1698175906
transform 1 0 16352 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_230
timestamp 1698175906
transform 1 0 2632 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_231
timestamp 1698175906
transform 1 0 6552 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_232
timestamp 1698175906
transform 1 0 10472 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_233
timestamp 1698175906
transform 1 0 14392 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_234
timestamp 1698175906
transform 1 0 18312 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_235
timestamp 1698175906
transform 1 0 4592 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_236
timestamp 1698175906
transform 1 0 8512 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_237
timestamp 1698175906
transform 1 0 12432 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_238
timestamp 1698175906
transform 1 0 16352 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_239
timestamp 1698175906
transform 1 0 2632 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_240
timestamp 1698175906
transform 1 0 6552 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_241
timestamp 1698175906
transform 1 0 10472 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_242
timestamp 1698175906
transform 1 0 14392 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_243
timestamp 1698175906
transform 1 0 18312 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_244
timestamp 1698175906
transform 1 0 4592 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_245
timestamp 1698175906
transform 1 0 8512 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_246
timestamp 1698175906
transform 1 0 12432 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_247
timestamp 1698175906
transform 1 0 16352 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_248
timestamp 1698175906
transform 1 0 2632 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_249
timestamp 1698175906
transform 1 0 6552 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_250
timestamp 1698175906
transform 1 0 10472 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_251
timestamp 1698175906
transform 1 0 14392 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_252
timestamp 1698175906
transform 1 0 18312 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_253
timestamp 1698175906
transform 1 0 4592 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_254
timestamp 1698175906
transform 1 0 8512 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_255
timestamp 1698175906
transform 1 0 12432 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_256
timestamp 1698175906
transform 1 0 16352 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_257
timestamp 1698175906
transform 1 0 2632 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_258
timestamp 1698175906
transform 1 0 6552 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_259
timestamp 1698175906
transform 1 0 10472 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_260
timestamp 1698175906
transform 1 0 14392 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_261
timestamp 1698175906
transform 1 0 18312 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_262
timestamp 1698175906
transform 1 0 4592 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_263
timestamp 1698175906
transform 1 0 8512 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_264
timestamp 1698175906
transform 1 0 12432 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_265
timestamp 1698175906
transform 1 0 16352 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_266
timestamp 1698175906
transform 1 0 2632 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_267
timestamp 1698175906
transform 1 0 6552 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_268
timestamp 1698175906
transform 1 0 10472 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_269
timestamp 1698175906
transform 1 0 14392 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_270
timestamp 1698175906
transform 1 0 18312 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_271
timestamp 1698175906
transform 1 0 4592 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_272
timestamp 1698175906
transform 1 0 8512 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_273
timestamp 1698175906
transform 1 0 12432 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_274
timestamp 1698175906
transform 1 0 16352 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_275
timestamp 1698175906
transform 1 0 2632 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_276
timestamp 1698175906
transform 1 0 6552 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_277
timestamp 1698175906
transform 1 0 10472 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_278
timestamp 1698175906
transform 1 0 14392 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_279
timestamp 1698175906
transform 1 0 18312 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_280
timestamp 1698175906
transform 1 0 4592 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_281
timestamp 1698175906
transform 1 0 8512 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_282
timestamp 1698175906
transform 1 0 12432 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_283
timestamp 1698175906
transform 1 0 16352 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_284
timestamp 1698175906
transform 1 0 2632 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_285
timestamp 1698175906
transform 1 0 6552 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_286
timestamp 1698175906
transform 1 0 10472 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_287
timestamp 1698175906
transform 1 0 14392 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_288
timestamp 1698175906
transform 1 0 18312 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_289
timestamp 1698175906
transform 1 0 4592 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_290
timestamp 1698175906
transform 1 0 8512 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_291
timestamp 1698175906
transform 1 0 12432 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_292
timestamp 1698175906
transform 1 0 16352 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_293
timestamp 1698175906
transform 1 0 2576 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_294
timestamp 1698175906
transform 1 0 4480 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_295
timestamp 1698175906
transform 1 0 6384 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_296
timestamp 1698175906
transform 1 0 8288 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_297
timestamp 1698175906
transform 1 0 10192 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_298
timestamp 1698175906
transform 1 0 12096 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_299
timestamp 1698175906
transform 1 0 14000 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_300
timestamp 1698175906
transform 1 0 15904 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_301
timestamp 1698175906
transform 1 0 17808 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_302
timestamp 1698175906
transform 1 0 19712 0 1 18816
box -43 -43 155 435
<< labels >>
flabel metal3 s 0 12768 400 12824 0 FreeSans 224 0 0 0 clk
port 0 nsew signal input
flabel metal2 s 8400 20600 8456 21000 0 FreeSans 224 90 0 0 segm[0]
port 1 nsew signal tristate
flabel metal3 s 20600 8064 21000 8120 0 FreeSans 224 0 0 0 segm[10]
port 2 nsew signal tristate
flabel metal3 s 20600 10416 21000 10472 0 FreeSans 224 0 0 0 segm[11]
port 3 nsew signal tristate
flabel metal3 s 20600 10080 21000 10136 0 FreeSans 224 0 0 0 segm[12]
port 4 nsew signal tristate
flabel metal3 s 20600 11424 21000 11480 0 FreeSans 224 0 0 0 segm[13]
port 5 nsew signal tristate
flabel metal3 s 20600 8736 21000 8792 0 FreeSans 224 0 0 0 segm[1]
port 6 nsew signal tristate
flabel metal3 s 20600 10752 21000 10808 0 FreeSans 224 0 0 0 segm[2]
port 7 nsew signal tristate
flabel metal2 s 12432 20600 12488 21000 0 FreeSans 224 90 0 0 segm[3]
port 8 nsew signal tristate
flabel metal3 s 20600 9072 21000 9128 0 FreeSans 224 0 0 0 segm[4]
port 9 nsew signal tristate
flabel metal2 s 11760 20600 11816 21000 0 FreeSans 224 90 0 0 segm[5]
port 10 nsew signal tristate
flabel metal2 s 11760 0 11816 400 0 FreeSans 224 90 0 0 segm[6]
port 11 nsew signal tristate
flabel metal2 s 11424 0 11480 400 0 FreeSans 224 90 0 0 segm[7]
port 12 nsew signal tristate
flabel metal3 s 20600 9744 21000 9800 0 FreeSans 224 0 0 0 segm[8]
port 13 nsew signal tristate
flabel metal3 s 20600 9408 21000 9464 0 FreeSans 224 0 0 0 segm[9]
port 14 nsew signal tristate
flabel metal3 s 20600 8400 21000 8456 0 FreeSans 224 0 0 0 sel[0]
port 15 nsew signal tristate
flabel metal3 s 0 8400 400 8456 0 FreeSans 224 0 0 0 sel[10]
port 16 nsew signal tristate
flabel metal3 s 0 12432 400 12488 0 FreeSans 224 0 0 0 sel[11]
port 17 nsew signal tristate
flabel metal3 s 20600 11088 21000 11144 0 FreeSans 224 0 0 0 sel[1]
port 18 nsew signal tristate
flabel metal2 s 10416 0 10472 400 0 FreeSans 224 90 0 0 sel[2]
port 19 nsew signal tristate
flabel metal3 s 20600 12096 21000 12152 0 FreeSans 224 0 0 0 sel[3]
port 20 nsew signal tristate
flabel metal2 s 12096 20600 12152 21000 0 FreeSans 224 90 0 0 sel[4]
port 21 nsew signal tristate
flabel metal3 s 0 10752 400 10808 0 FreeSans 224 0 0 0 sel[5]
port 22 nsew signal tristate
flabel metal3 s 0 11424 400 11480 0 FreeSans 224 0 0 0 sel[6]
port 23 nsew signal tristate
flabel metal3 s 0 12096 400 12152 0 FreeSans 224 0 0 0 sel[7]
port 24 nsew signal tristate
flabel metal2 s 9072 0 9128 400 0 FreeSans 224 90 0 0 sel[8]
port 25 nsew signal tristate
flabel metal3 s 0 9072 400 9128 0 FreeSans 224 0 0 0 sel[9]
port 26 nsew signal tristate
flabel metal4 s 2224 1538 2384 19238 0 FreeSans 640 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 17584 1538 17744 19238 0 FreeSans 640 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 9904 1538 10064 19238 0 FreeSans 640 90 0 0 vss
port 28 nsew ground bidirectional
rlabel metal1 10500 19208 10500 19208 0 vdd
rlabel metal1 10500 18816 10500 18816 0 vss
rlabel metal2 7308 12152 7308 12152 0 _000_
rlabel metal2 7252 8204 7252 8204 0 _001_
rlabel metal2 6748 10864 6748 10864 0 _002_
rlabel metal2 7532 11032 7532 11032 0 _003_
rlabel metal2 8876 8400 8876 8400 0 _004_
rlabel metal2 7420 9380 7420 9380 0 _005_
rlabel metal2 9240 12012 9240 12012 0 _006_
rlabel metal2 8988 10276 8988 10276 0 _007_
rlabel metal2 11732 12040 11732 12040 0 _008_
rlabel metal2 9828 8036 9828 8036 0 _009_
rlabel metal2 13300 10388 13300 10388 0 _010_
rlabel metal2 14084 9044 14084 9044 0 _011_
rlabel metal2 11172 8120 11172 8120 0 _012_
rlabel metal2 13244 11396 13244 11396 0 _013_
rlabel metal2 7084 8512 7084 8512 0 _014_
rlabel metal2 7812 11928 7812 11928 0 _015_
rlabel metal2 11172 12572 11172 12572 0 _016_
rlabel metal2 12236 9016 12236 9016 0 _017_
rlabel metal2 11284 10108 11284 10108 0 _018_
rlabel metal3 7252 9156 7252 9156 0 _019_
rlabel metal2 11340 12236 11340 12236 0 _020_
rlabel metal2 12404 9660 12404 9660 0 _021_
rlabel metal2 11452 10332 11452 10332 0 _022_
rlabel metal2 7364 9016 7364 9016 0 _023_
rlabel metal2 10836 11032 10836 11032 0 _024_
rlabel metal3 9968 10780 9968 10780 0 _025_
rlabel metal2 7392 10836 7392 10836 0 _026_
rlabel metal3 7224 11172 7224 11172 0 _027_
rlabel metal2 7252 11844 7252 11844 0 _028_
rlabel metal3 10220 11172 10220 11172 0 _029_
rlabel metal2 7532 12796 7532 12796 0 _030_
rlabel metal2 7532 12124 7532 12124 0 _031_
rlabel metal2 9884 8848 9884 8848 0 _032_
rlabel metal3 9800 8764 9800 8764 0 _033_
rlabel metal2 10724 11648 10724 11648 0 _034_
rlabel metal3 11676 12348 11676 12348 0 _035_
rlabel metal2 6972 9072 6972 9072 0 _036_
rlabel metal2 10752 8820 10752 8820 0 _037_
rlabel metal2 7532 8708 7532 8708 0 _038_
rlabel metal3 8708 8428 8708 8428 0 _039_
rlabel metal2 6916 11172 6916 11172 0 _040_
rlabel metal2 7196 11172 7196 11172 0 _041_
rlabel metal2 9660 9492 9660 9492 0 _042_
rlabel metal2 11368 10388 11368 10388 0 _043_
rlabel metal2 11340 10108 11340 10108 0 _044_
rlabel metal2 10080 9492 10080 9492 0 _045_
rlabel metal2 7532 10920 7532 10920 0 _046_
rlabel metal2 10556 11928 10556 11928 0 _047_
rlabel metal2 9044 12152 9044 12152 0 _048_
rlabel metal3 11340 11284 11340 11284 0 _049_
rlabel metal2 9268 9044 9268 9044 0 _050_
rlabel metal2 9044 10388 9044 10388 0 _051_
rlabel metal3 9912 9604 9912 9604 0 _052_
rlabel metal2 13860 11368 13860 11368 0 _053_
rlabel metal2 13020 12208 13020 12208 0 _054_
rlabel metal2 13524 10836 13524 10836 0 _055_
rlabel metal3 10052 8428 10052 8428 0 _056_
rlabel metal2 9716 8512 9716 8512 0 _057_
rlabel metal2 9996 8484 9996 8484 0 _058_
rlabel metal2 13580 9940 13580 9940 0 _059_
rlabel metal2 13524 9436 13524 9436 0 _060_
rlabel metal2 14140 9072 14140 9072 0 _061_
rlabel metal2 11396 8456 11396 8456 0 _062_
rlabel metal2 13608 11564 13608 11564 0 _063_
rlabel metal2 7588 8624 7588 8624 0 _064_
rlabel metal2 7644 12488 7644 12488 0 _065_
rlabel metal2 11676 11032 11676 11032 0 _066_
rlabel metal3 1239 12796 1239 12796 0 clk
rlabel metal2 11676 10220 11676 10220 0 clknet_0_clk
rlabel metal2 7084 10430 7084 10430 0 clknet_1_0__leaf_clk
rlabel metal2 11844 8708 11844 8708 0 clknet_1_1__leaf_clk
rlabel metal3 9772 9268 9772 9268 0 dut29.count\[0\]
rlabel metal2 9436 9800 9436 9800 0 dut29.count\[1\]
rlabel metal2 10164 12180 10164 12180 0 dut29.count\[2\]
rlabel metal2 10444 12572 10444 12572 0 dut29.count\[3\]
rlabel metal2 15036 9184 15036 9184 0 net1
rlabel metal2 11900 5124 11900 5124 0 net10
rlabel metal2 12292 4662 12292 4662 0 net11
rlabel metal2 18844 9520 18844 9520 0 net12
rlabel metal3 18844 9156 18844 9156 0 net13
rlabel metal2 15372 8652 15372 8652 0 net14
rlabel metal2 6020 8596 6020 8596 0 net15
rlabel metal2 6748 12768 6748 12768 0 net16
rlabel metal3 15442 10836 15442 10836 0 net17
rlabel metal2 10556 2982 10556 2982 0 net18
rlabel metal2 18844 12180 18844 12180 0 net19
rlabel metal2 12348 10556 12348 10556 0 net2
rlabel metal3 12432 13244 12432 13244 0 net20
rlabel metal2 6748 10724 6748 10724 0 net21
rlabel metal2 5684 11144 5684 11144 0 net22
rlabel metal2 6244 12320 6244 12320 0 net23
rlabel metal3 8568 8092 8568 8092 0 net24
rlabel metal2 2156 9184 2156 9184 0 net25
rlabel metal3 14140 9604 14140 9604 0 net26
rlabel metal2 8484 18956 8484 18956 0 net27
rlabel metal2 18956 9688 18956 9688 0 net3
rlabel metal2 14308 11396 14308 11396 0 net4
rlabel metal2 18844 8568 18844 8568 0 net5
rlabel metal2 14588 10752 14588 10752 0 net6
rlabel metal2 12684 15456 12684 15456 0 net7
rlabel metal2 18788 9156 18788 9156 0 net8
rlabel metal2 12460 16226 12460 16226 0 net9
rlabel metal2 20020 7840 20020 7840 0 segm[10]
rlabel metal3 20321 10444 20321 10444 0 segm[11]
rlabel metal3 20321 10108 20321 10108 0 segm[12]
rlabel metal3 20321 11452 20321 11452 0 segm[13]
rlabel metal2 19684 8624 19684 8624 0 segm[1]
rlabel metal2 20020 10752 20020 10752 0 segm[2]
rlabel metal2 12460 20265 12460 20265 0 segm[3]
rlabel metal2 19964 8988 19964 8988 0 segm[4]
rlabel metal2 11788 19873 11788 19873 0 segm[5]
rlabel metal2 11788 1491 11788 1491 0 segm[6]
rlabel metal2 11452 1099 11452 1099 0 segm[7]
rlabel metal2 20020 9744 20020 9744 0 segm[8]
rlabel metal2 20020 9296 20020 9296 0 segm[9]
rlabel metal2 19908 8232 19908 8232 0 sel[0]
rlabel metal3 679 8428 679 8428 0 sel[10]
rlabel metal3 679 12460 679 12460 0 sel[11]
rlabel metal2 20020 11172 20020 11172 0 sel[1]
rlabel metal2 10444 1099 10444 1099 0 sel[2]
rlabel metal2 20020 12180 20020 12180 0 sel[3]
rlabel metal2 12124 19677 12124 19677 0 sel[4]
rlabel metal3 679 10780 679 10780 0 sel[5]
rlabel metal3 679 11452 679 11452 0 sel[6]
rlabel metal3 679 12124 679 12124 0 sel[7]
rlabel metal2 9100 1099 9100 1099 0 sel[8]
rlabel metal3 679 9100 679 9100 0 sel[9]
<< properties >>
string FIXED_BBOX 0 0 21000 21000
<< end >>
