magic
tech gf180mcuD
magscale 1 5
timestamp 1699644639
<< metal1 >>
rect 672 19221 20328 19238
rect 672 19195 2239 19221
rect 2265 19195 2291 19221
rect 2317 19195 2343 19221
rect 2369 19195 17599 19221
rect 17625 19195 17651 19221
rect 17677 19195 17703 19221
rect 17729 19195 20328 19221
rect 672 19178 20328 19195
rect 9031 19137 9057 19143
rect 9031 19105 9057 19111
rect 10879 19137 10905 19143
rect 10879 19105 10905 19111
rect 12783 19137 12809 19143
rect 12783 19105 12809 19111
rect 14687 19137 14713 19143
rect 14687 19105 14713 19111
rect 8521 18999 8527 19025
rect 8553 18999 8559 19025
rect 10369 18999 10375 19025
rect 10401 18999 10407 19025
rect 12273 18999 12279 19025
rect 12305 18999 12311 19025
rect 14289 18999 14295 19025
rect 14321 18999 14327 19025
rect 672 18829 20328 18846
rect 672 18803 9919 18829
rect 9945 18803 9971 18829
rect 9997 18803 10023 18829
rect 10049 18803 20328 18829
rect 672 18786 20328 18803
rect 10039 18745 10065 18751
rect 10039 18713 10065 18719
rect 12615 18745 12641 18751
rect 12615 18713 12641 18719
rect 13399 18745 13425 18751
rect 13399 18713 13425 18719
rect 9529 18607 9535 18633
rect 9561 18607 9567 18633
rect 12889 18607 12895 18633
rect 12921 18607 12927 18633
rect 672 18437 20328 18454
rect 672 18411 2239 18437
rect 2265 18411 2291 18437
rect 2317 18411 2343 18437
rect 2369 18411 17599 18437
rect 17625 18411 17651 18437
rect 17677 18411 17703 18437
rect 17729 18411 20328 18437
rect 672 18394 20328 18411
rect 672 18045 20328 18062
rect 672 18019 9919 18045
rect 9945 18019 9971 18045
rect 9997 18019 10023 18045
rect 10049 18019 20328 18045
rect 672 18002 20328 18019
rect 672 17653 20328 17670
rect 672 17627 2239 17653
rect 2265 17627 2291 17653
rect 2317 17627 2343 17653
rect 2369 17627 17599 17653
rect 17625 17627 17651 17653
rect 17677 17627 17703 17653
rect 17729 17627 20328 17653
rect 672 17610 20328 17627
rect 672 17261 20328 17278
rect 672 17235 9919 17261
rect 9945 17235 9971 17261
rect 9997 17235 10023 17261
rect 10049 17235 20328 17261
rect 672 17218 20328 17235
rect 672 16869 20328 16886
rect 672 16843 2239 16869
rect 2265 16843 2291 16869
rect 2317 16843 2343 16869
rect 2369 16843 17599 16869
rect 17625 16843 17651 16869
rect 17677 16843 17703 16869
rect 17729 16843 20328 16869
rect 672 16826 20328 16843
rect 672 16477 20328 16494
rect 672 16451 9919 16477
rect 9945 16451 9971 16477
rect 9997 16451 10023 16477
rect 10049 16451 20328 16477
rect 672 16434 20328 16451
rect 672 16085 20328 16102
rect 672 16059 2239 16085
rect 2265 16059 2291 16085
rect 2317 16059 2343 16085
rect 2369 16059 17599 16085
rect 17625 16059 17651 16085
rect 17677 16059 17703 16085
rect 17729 16059 20328 16085
rect 672 16042 20328 16059
rect 672 15693 20328 15710
rect 672 15667 9919 15693
rect 9945 15667 9971 15693
rect 9997 15667 10023 15693
rect 10049 15667 20328 15693
rect 672 15650 20328 15667
rect 672 15301 20328 15318
rect 672 15275 2239 15301
rect 2265 15275 2291 15301
rect 2317 15275 2343 15301
rect 2369 15275 17599 15301
rect 17625 15275 17651 15301
rect 17677 15275 17703 15301
rect 17729 15275 20328 15301
rect 672 15258 20328 15275
rect 672 14909 20328 14926
rect 672 14883 9919 14909
rect 9945 14883 9971 14909
rect 9997 14883 10023 14909
rect 10049 14883 20328 14909
rect 672 14866 20328 14883
rect 672 14517 20328 14534
rect 672 14491 2239 14517
rect 2265 14491 2291 14517
rect 2317 14491 2343 14517
rect 2369 14491 17599 14517
rect 17625 14491 17651 14517
rect 17677 14491 17703 14517
rect 17729 14491 20328 14517
rect 672 14474 20328 14491
rect 9529 14351 9535 14377
rect 9561 14351 9567 14377
rect 12105 14351 12111 14377
rect 12137 14351 12143 14377
rect 9759 14321 9785 14327
rect 12335 14321 12361 14327
rect 8129 14295 8135 14321
rect 8161 14295 8167 14321
rect 10705 14295 10711 14321
rect 10737 14295 10743 14321
rect 11041 14295 11047 14321
rect 11073 14295 11079 14321
rect 9759 14289 9785 14295
rect 12335 14289 12361 14295
rect 8465 14239 8471 14265
rect 8497 14239 8503 14265
rect 672 14125 20328 14142
rect 672 14099 9919 14125
rect 9945 14099 9971 14125
rect 9997 14099 10023 14125
rect 10049 14099 20328 14125
rect 672 14082 20328 14099
rect 8415 14041 8441 14047
rect 8415 14009 8441 14015
rect 10879 14041 10905 14047
rect 10879 14009 10905 14015
rect 11271 14041 11297 14047
rect 11271 14009 11297 14015
rect 10767 13985 10793 13991
rect 10767 13953 10793 13959
rect 11159 13985 11185 13991
rect 11159 13953 11185 13959
rect 10711 13929 10737 13935
rect 8913 13903 8919 13929
rect 8945 13903 8951 13929
rect 10711 13897 10737 13903
rect 11327 13929 11353 13935
rect 11327 13897 11353 13903
rect 9249 13847 9255 13873
rect 9281 13847 9287 13873
rect 10313 13847 10319 13873
rect 10345 13847 10351 13873
rect 672 13733 20328 13750
rect 672 13707 2239 13733
rect 2265 13707 2291 13733
rect 2317 13707 2343 13733
rect 2369 13707 17599 13733
rect 17625 13707 17651 13733
rect 17677 13707 17703 13733
rect 17729 13707 20328 13733
rect 672 13690 20328 13707
rect 9647 13649 9673 13655
rect 9647 13617 9673 13623
rect 8695 13593 8721 13599
rect 8465 13567 8471 13593
rect 8497 13567 8503 13593
rect 13225 13567 13231 13593
rect 13257 13567 13263 13593
rect 8695 13561 8721 13567
rect 9031 13537 9057 13543
rect 7065 13511 7071 13537
rect 7097 13511 7103 13537
rect 9031 13505 9057 13511
rect 9311 13537 9337 13543
rect 9311 13505 9337 13511
rect 9479 13537 9505 13543
rect 11825 13511 11831 13537
rect 11857 13511 11863 13537
rect 9479 13505 9505 13511
rect 9143 13481 9169 13487
rect 7401 13455 7407 13481
rect 7433 13455 7439 13481
rect 9143 13449 9169 13455
rect 9199 13481 9225 13487
rect 9199 13449 9225 13455
rect 9423 13481 9449 13487
rect 9423 13449 9449 13455
rect 9703 13481 9729 13487
rect 13455 13481 13481 13487
rect 12161 13455 12167 13481
rect 12193 13455 12199 13481
rect 9703 13449 9729 13455
rect 13455 13449 13481 13455
rect 672 13341 20328 13358
rect 672 13315 9919 13341
rect 9945 13315 9971 13341
rect 9997 13315 10023 13341
rect 10049 13315 20328 13341
rect 672 13298 20328 13315
rect 7463 13257 7489 13263
rect 7463 13225 7489 13231
rect 7911 13257 7937 13263
rect 7911 13225 7937 13231
rect 8807 13257 8833 13263
rect 9927 13257 9953 13263
rect 9361 13231 9367 13257
rect 9393 13231 9399 13257
rect 8807 13225 8833 13231
rect 9927 13225 9953 13231
rect 9983 13257 10009 13263
rect 9983 13225 10009 13231
rect 12167 13257 12193 13263
rect 12167 13225 12193 13231
rect 7183 13201 7209 13207
rect 7183 13169 7209 13175
rect 8695 13201 8721 13207
rect 8695 13169 8721 13175
rect 12839 13201 12865 13207
rect 12839 13169 12865 13175
rect 7127 13145 7153 13151
rect 2137 13119 2143 13145
rect 2169 13119 2175 13145
rect 6953 13119 6959 13145
rect 6985 13119 6991 13145
rect 7127 13113 7153 13119
rect 8919 13145 8945 13151
rect 9535 13145 9561 13151
rect 9871 13145 9897 13151
rect 11383 13145 11409 13151
rect 9025 13119 9031 13145
rect 9057 13119 9063 13145
rect 9753 13119 9759 13145
rect 9785 13119 9791 13145
rect 10089 13119 10095 13145
rect 10121 13119 10127 13145
rect 8919 13113 8945 13119
rect 9535 13113 9561 13119
rect 9871 13113 9897 13119
rect 11383 13113 11409 13119
rect 11439 13145 11465 13151
rect 11439 13113 11465 13119
rect 11663 13145 11689 13151
rect 12111 13145 12137 13151
rect 11769 13119 11775 13145
rect 11801 13119 11807 13145
rect 11881 13119 11887 13145
rect 11913 13119 11919 13145
rect 11663 13113 11689 13119
rect 12111 13113 12137 13119
rect 12223 13145 12249 13151
rect 12223 13113 12249 13119
rect 12783 13145 12809 13151
rect 18825 13119 18831 13145
rect 18857 13119 18863 13145
rect 12783 13113 12809 13119
rect 7967 13089 7993 13095
rect 5497 13063 5503 13089
rect 5529 13063 5535 13089
rect 6561 13063 6567 13089
rect 6593 13063 6599 13089
rect 7967 13057 7993 13063
rect 8863 13089 8889 13095
rect 8863 13057 8889 13063
rect 11551 13089 11577 13095
rect 11551 13057 11577 13063
rect 11999 13089 12025 13095
rect 19945 13063 19951 13089
rect 19977 13063 19983 13089
rect 11999 13057 12025 13063
rect 967 13033 993 13039
rect 967 13001 993 13007
rect 7183 13033 7209 13039
rect 7183 13001 7209 13007
rect 672 12949 20328 12966
rect 672 12923 2239 12949
rect 2265 12923 2291 12949
rect 2317 12923 2343 12949
rect 2369 12923 17599 12949
rect 17625 12923 17651 12949
rect 17677 12923 17703 12949
rect 17729 12923 20328 12949
rect 672 12906 20328 12923
rect 10929 12839 10935 12865
rect 10961 12839 10967 12865
rect 20007 12809 20033 12815
rect 11713 12783 11719 12809
rect 11745 12783 11751 12809
rect 12777 12783 12783 12809
rect 12809 12783 12815 12809
rect 20007 12777 20033 12783
rect 6903 12753 6929 12759
rect 10655 12753 10681 12759
rect 9753 12727 9759 12753
rect 9785 12727 9791 12753
rect 6903 12721 6929 12727
rect 10655 12721 10681 12727
rect 10767 12753 10793 12759
rect 11377 12727 11383 12753
rect 11409 12727 11415 12753
rect 14625 12727 14631 12753
rect 14657 12727 14663 12753
rect 18825 12727 18831 12753
rect 18857 12727 18863 12753
rect 10767 12721 10793 12727
rect 6735 12697 6761 12703
rect 6735 12665 6761 12671
rect 6791 12697 6817 12703
rect 13903 12697 13929 12703
rect 9865 12671 9871 12697
rect 9897 12671 9903 12697
rect 14737 12671 14743 12697
rect 14769 12671 14775 12697
rect 6791 12665 6817 12671
rect 13903 12665 13929 12671
rect 7127 12641 7153 12647
rect 7127 12609 7153 12615
rect 13007 12641 13033 12647
rect 13007 12609 13033 12615
rect 13231 12641 13257 12647
rect 13231 12609 13257 12615
rect 13847 12641 13873 12647
rect 13847 12609 13873 12615
rect 672 12557 20328 12574
rect 672 12531 9919 12557
rect 9945 12531 9971 12557
rect 9997 12531 10023 12557
rect 10049 12531 20328 12557
rect 672 12514 20328 12531
rect 6511 12473 6537 12479
rect 6511 12441 6537 12447
rect 11999 12473 12025 12479
rect 11999 12441 12025 12447
rect 13063 12473 13089 12479
rect 13063 12441 13089 12447
rect 13119 12473 13145 12479
rect 13119 12441 13145 12447
rect 9479 12417 9505 12423
rect 9479 12385 9505 12391
rect 9703 12417 9729 12423
rect 9703 12385 9729 12391
rect 10039 12417 10065 12423
rect 12111 12417 12137 12423
rect 11657 12391 11663 12417
rect 11689 12391 11695 12417
rect 13785 12391 13791 12417
rect 13817 12391 13823 12417
rect 10039 12385 10065 12391
rect 12111 12385 12137 12391
rect 9311 12361 9337 12367
rect 11943 12361 11969 12367
rect 11545 12335 11551 12361
rect 11577 12335 11583 12361
rect 9311 12329 9337 12335
rect 11943 12329 11969 12335
rect 12223 12361 12249 12367
rect 12223 12329 12249 12335
rect 12951 12361 12977 12367
rect 12951 12329 12977 12335
rect 13007 12361 13033 12367
rect 13225 12335 13231 12361
rect 13257 12335 13263 12361
rect 13393 12335 13399 12361
rect 13425 12335 13431 12361
rect 13007 12329 13033 12335
rect 9977 12279 9983 12305
rect 10009 12279 10015 12305
rect 14849 12279 14855 12305
rect 14881 12279 14887 12305
rect 9647 12249 9673 12255
rect 9647 12217 9673 12223
rect 9815 12249 9841 12255
rect 9815 12217 9841 12223
rect 10151 12249 10177 12255
rect 10151 12217 10177 12223
rect 672 12165 20328 12182
rect 672 12139 2239 12165
rect 2265 12139 2291 12165
rect 2317 12139 2343 12165
rect 2369 12139 17599 12165
rect 17625 12139 17651 12165
rect 17677 12139 17703 12165
rect 17729 12139 20328 12165
rect 672 12122 20328 12139
rect 10431 12081 10457 12087
rect 10431 12049 10457 12055
rect 967 12025 993 12031
rect 7071 12025 7097 12031
rect 8919 12025 8945 12031
rect 20007 12025 20033 12031
rect 4937 11999 4943 12025
rect 4969 11999 4975 12025
rect 8689 11999 8695 12025
rect 8721 11999 8727 12025
rect 11601 11999 11607 12025
rect 11633 11999 11639 12025
rect 967 11993 993 11999
rect 7071 11993 7097 11999
rect 8919 11993 8945 11999
rect 20007 11993 20033 11999
rect 6847 11969 6873 11975
rect 9423 11969 9449 11975
rect 2137 11943 2143 11969
rect 2169 11943 2175 11969
rect 6393 11943 6399 11969
rect 6425 11943 6431 11969
rect 7233 11943 7239 11969
rect 7265 11943 7271 11969
rect 6847 11937 6873 11943
rect 9423 11937 9449 11943
rect 10095 11969 10121 11975
rect 13847 11969 13873 11975
rect 10705 11943 10711 11969
rect 10737 11943 10743 11969
rect 13001 11943 13007 11969
rect 13033 11943 13039 11969
rect 18825 11943 18831 11969
rect 18857 11943 18863 11969
rect 10095 11937 10121 11943
rect 13847 11937 13873 11943
rect 6791 11913 6817 11919
rect 13903 11913 13929 11919
rect 6001 11887 6007 11913
rect 6033 11887 6039 11913
rect 7625 11887 7631 11913
rect 7657 11887 7663 11913
rect 9249 11887 9255 11913
rect 9281 11887 9287 11913
rect 9529 11887 9535 11913
rect 9561 11887 9567 11913
rect 9809 11887 9815 11913
rect 9841 11887 9847 11913
rect 12665 11887 12671 11913
rect 12697 11887 12703 11913
rect 6791 11881 6817 11887
rect 13903 11881 13929 11887
rect 6679 11857 6705 11863
rect 6679 11825 6705 11831
rect 9087 11857 9113 11863
rect 10263 11857 10289 11863
rect 9641 11831 9647 11857
rect 9673 11831 9679 11857
rect 9087 11825 9113 11831
rect 10263 11825 10289 11831
rect 10375 11857 10401 11863
rect 13287 11857 13313 11863
rect 10817 11831 10823 11857
rect 10849 11831 10855 11857
rect 10375 11825 10401 11831
rect 13287 11825 13313 11831
rect 14015 11857 14041 11863
rect 14015 11825 14041 11831
rect 672 11773 20328 11790
rect 672 11747 9919 11773
rect 9945 11747 9971 11773
rect 9997 11747 10023 11773
rect 10049 11747 20328 11773
rect 672 11730 20328 11747
rect 6175 11689 6201 11695
rect 6175 11657 6201 11663
rect 9479 11689 9505 11695
rect 9479 11657 9505 11663
rect 12671 11689 12697 11695
rect 12671 11657 12697 11663
rect 13063 11689 13089 11695
rect 13063 11657 13089 11663
rect 6287 11633 6313 11639
rect 6287 11601 6313 11607
rect 6343 11633 6369 11639
rect 6343 11601 6369 11607
rect 7743 11633 7769 11639
rect 9255 11633 9281 11639
rect 8017 11607 8023 11633
rect 8049 11607 8055 11633
rect 7743 11601 7769 11607
rect 9255 11601 9281 11607
rect 9311 11633 9337 11639
rect 9311 11601 9337 11607
rect 11887 11633 11913 11639
rect 11887 11601 11913 11607
rect 9031 11577 9057 11583
rect 8129 11551 8135 11577
rect 8161 11551 8167 11577
rect 9031 11545 9057 11551
rect 9143 11577 9169 11583
rect 9143 11545 9169 11551
rect 10039 11577 10065 11583
rect 11047 11577 11073 11583
rect 10649 11551 10655 11577
rect 10681 11551 10687 11577
rect 10039 11545 10065 11551
rect 11047 11545 11073 11551
rect 11663 11577 11689 11583
rect 11663 11545 11689 11551
rect 12839 11577 12865 11583
rect 12839 11545 12865 11551
rect 12951 11577 12977 11583
rect 13281 11551 13287 11577
rect 13313 11551 13319 11577
rect 12951 11545 12977 11551
rect 7855 11521 7881 11527
rect 7681 11495 7687 11521
rect 7713 11495 7719 11521
rect 7855 11489 7881 11495
rect 9759 11521 9785 11527
rect 9759 11489 9785 11495
rect 9927 11521 9953 11527
rect 9927 11489 9953 11495
rect 10879 11521 10905 11527
rect 10879 11489 10905 11495
rect 11327 11521 11353 11527
rect 11327 11489 11353 11495
rect 11719 11521 11745 11527
rect 11719 11489 11745 11495
rect 12895 11521 12921 11527
rect 13673 11495 13679 11521
rect 13705 11495 13711 11521
rect 14737 11495 14743 11521
rect 14769 11495 14775 11521
rect 12895 11489 12921 11495
rect 8975 11465 9001 11471
rect 8975 11433 9001 11439
rect 10207 11465 10233 11471
rect 10207 11433 10233 11439
rect 11831 11465 11857 11471
rect 11831 11433 11857 11439
rect 672 11381 20328 11398
rect 672 11355 2239 11381
rect 2265 11355 2291 11381
rect 2317 11355 2343 11381
rect 2369 11355 17599 11381
rect 17625 11355 17651 11381
rect 17677 11355 17703 11381
rect 17729 11355 20328 11381
rect 672 11338 20328 11355
rect 12721 11271 12727 11297
rect 12753 11271 12759 11297
rect 967 11241 993 11247
rect 8913 11215 8919 11241
rect 8945 11215 8951 11241
rect 11153 11215 11159 11241
rect 11185 11215 11191 11241
rect 967 11209 993 11215
rect 7015 11185 7041 11191
rect 2137 11159 2143 11185
rect 2169 11159 2175 11185
rect 7015 11153 7041 11159
rect 7127 11185 7153 11191
rect 12223 11185 12249 11191
rect 9697 11159 9703 11185
rect 9729 11159 9735 11185
rect 10929 11159 10935 11185
rect 10961 11159 10967 11185
rect 7127 11153 7153 11159
rect 12223 11153 12249 11159
rect 12447 11185 12473 11191
rect 12447 11153 12473 11159
rect 12559 11185 12585 11191
rect 12945 11159 12951 11185
rect 12977 11159 12983 11185
rect 12559 11153 12585 11159
rect 7351 11129 7377 11135
rect 10985 11103 10991 11129
rect 11017 11103 11023 11129
rect 11433 11103 11439 11129
rect 11465 11103 11471 11129
rect 7351 11097 7377 11103
rect 6959 11073 6985 11079
rect 6959 11041 6985 11047
rect 7239 11073 7265 11079
rect 13057 11047 13063 11073
rect 13089 11047 13095 11073
rect 7239 11041 7265 11047
rect 672 10989 20328 11006
rect 672 10963 9919 10989
rect 9945 10963 9971 10989
rect 9997 10963 10023 10989
rect 10049 10963 20328 10989
rect 672 10946 20328 10963
rect 7743 10905 7769 10911
rect 7743 10873 7769 10879
rect 12671 10905 12697 10911
rect 12671 10873 12697 10879
rect 7687 10849 7713 10855
rect 6729 10823 6735 10849
rect 6761 10823 6767 10849
rect 8969 10823 8975 10849
rect 9001 10823 9007 10849
rect 7687 10817 7713 10823
rect 7799 10793 7825 10799
rect 2137 10767 2143 10793
rect 2169 10767 2175 10793
rect 7121 10767 7127 10793
rect 7153 10767 7159 10793
rect 7513 10767 7519 10793
rect 7545 10767 7551 10793
rect 7799 10761 7825 10767
rect 7911 10793 7937 10799
rect 7911 10761 7937 10767
rect 8135 10793 8161 10799
rect 8135 10761 8161 10767
rect 8247 10793 8273 10799
rect 9255 10793 9281 10799
rect 8857 10767 8863 10793
rect 8889 10767 8895 10793
rect 9585 10767 9591 10793
rect 9617 10767 9623 10793
rect 18825 10767 18831 10793
rect 18857 10767 18863 10793
rect 8247 10761 8273 10767
rect 9255 10761 9281 10767
rect 7351 10737 7377 10743
rect 5665 10711 5671 10737
rect 5697 10711 5703 10737
rect 7351 10705 7377 10711
rect 8191 10737 8217 10743
rect 8191 10705 8217 10711
rect 9143 10737 9169 10743
rect 13287 10737 13313 10743
rect 11321 10711 11327 10737
rect 11353 10711 11359 10737
rect 9143 10705 9169 10711
rect 13287 10705 13313 10711
rect 14575 10737 14601 10743
rect 14575 10705 14601 10711
rect 967 10681 993 10687
rect 14519 10681 14545 10687
rect 9417 10655 9423 10681
rect 9449 10655 9455 10681
rect 967 10649 993 10655
rect 14519 10649 14545 10655
rect 20007 10681 20033 10687
rect 20007 10649 20033 10655
rect 672 10597 20328 10614
rect 672 10571 2239 10597
rect 2265 10571 2291 10597
rect 2317 10571 2343 10597
rect 2369 10571 17599 10597
rect 17625 10571 17651 10597
rect 17677 10571 17703 10597
rect 17729 10571 20328 10597
rect 672 10554 20328 10571
rect 6063 10513 6089 10519
rect 6063 10481 6089 10487
rect 9199 10513 9225 10519
rect 9199 10481 9225 10487
rect 10711 10457 10737 10463
rect 7121 10431 7127 10457
rect 7153 10431 7159 10457
rect 8185 10431 8191 10457
rect 8217 10431 8223 10457
rect 10711 10425 10737 10431
rect 11103 10457 11129 10463
rect 11103 10425 11129 10431
rect 6119 10401 6145 10407
rect 6119 10369 6145 10375
rect 6343 10401 6369 10407
rect 8359 10401 8385 10407
rect 10823 10401 10849 10407
rect 6785 10375 6791 10401
rect 6817 10375 6823 10401
rect 8745 10375 8751 10401
rect 8777 10375 8783 10401
rect 9473 10375 9479 10401
rect 9505 10375 9511 10401
rect 9641 10375 9647 10401
rect 9673 10375 9679 10401
rect 10089 10375 10095 10401
rect 10121 10375 10127 10401
rect 10313 10375 10319 10401
rect 10345 10375 10351 10401
rect 6343 10369 6369 10375
rect 8359 10369 8385 10375
rect 10823 10369 10849 10375
rect 11047 10401 11073 10407
rect 11321 10375 11327 10401
rect 11353 10375 11359 10401
rect 11047 10369 11073 10375
rect 9031 10345 9057 10351
rect 8857 10319 8863 10345
rect 8889 10319 8895 10345
rect 10257 10319 10263 10345
rect 10289 10319 10295 10345
rect 13337 10319 13343 10345
rect 13369 10319 13375 10345
rect 9031 10313 9057 10319
rect 6063 10289 6089 10295
rect 9143 10289 9169 10295
rect 11159 10289 11185 10295
rect 8521 10263 8527 10289
rect 8553 10263 8559 10289
rect 9361 10263 9367 10289
rect 9393 10263 9399 10289
rect 6063 10257 6089 10263
rect 9143 10257 9169 10263
rect 11159 10257 11185 10263
rect 20119 10289 20145 10295
rect 20119 10257 20145 10263
rect 672 10205 20328 10222
rect 672 10179 9919 10205
rect 9945 10179 9971 10205
rect 9997 10179 10023 10205
rect 10049 10179 20328 10205
rect 672 10162 20328 10179
rect 8303 10121 8329 10127
rect 7849 10095 7855 10121
rect 7881 10095 7887 10121
rect 8303 10089 8329 10095
rect 11383 10121 11409 10127
rect 11383 10089 11409 10095
rect 6455 10065 6481 10071
rect 6455 10033 6481 10039
rect 6511 10065 6537 10071
rect 6511 10033 6537 10039
rect 6791 10065 6817 10071
rect 8247 10065 8273 10071
rect 11719 10065 11745 10071
rect 12279 10065 12305 10071
rect 7457 10039 7463 10065
rect 7489 10039 7495 10065
rect 7737 10039 7743 10065
rect 7769 10039 7775 10065
rect 9585 10039 9591 10065
rect 9617 10039 9623 10065
rect 10089 10039 10095 10065
rect 10121 10039 10127 10065
rect 11881 10039 11887 10065
rect 11913 10039 11919 10065
rect 6791 10033 6817 10039
rect 8247 10033 8273 10039
rect 11719 10033 11745 10039
rect 12279 10033 12305 10039
rect 12391 10065 12417 10071
rect 12391 10033 12417 10039
rect 13063 10065 13089 10071
rect 13063 10033 13089 10039
rect 7911 10009 7937 10015
rect 11271 10009 11297 10015
rect 6281 9983 6287 10009
rect 6313 9983 6319 10009
rect 9137 9983 9143 10009
rect 9169 9983 9175 10009
rect 9305 9983 9311 10009
rect 9337 9983 9343 10009
rect 10145 9983 10151 10009
rect 10177 9983 10183 10009
rect 7911 9977 7937 9983
rect 11271 9977 11297 9983
rect 11607 10009 11633 10015
rect 11607 9977 11633 9983
rect 12223 10009 12249 10015
rect 12223 9977 12249 9983
rect 12727 10009 12753 10015
rect 12727 9977 12753 9983
rect 12951 10009 12977 10015
rect 13449 9983 13455 10009
rect 13481 9983 13487 10009
rect 18825 9983 18831 10009
rect 18857 9983 18863 10009
rect 12951 9977 12977 9983
rect 8751 9953 8777 9959
rect 11327 9953 11353 9959
rect 4825 9927 4831 9953
rect 4857 9927 4863 9953
rect 5889 9927 5895 9953
rect 5921 9927 5927 9953
rect 9081 9927 9087 9953
rect 9113 9927 9119 9953
rect 9361 9927 9367 9953
rect 9393 9927 9399 9953
rect 8751 9921 8777 9927
rect 11327 9921 11353 9927
rect 12839 9953 12865 9959
rect 13001 9927 13007 9953
rect 13033 9927 13039 9953
rect 13841 9927 13847 9953
rect 13873 9927 13879 9953
rect 14905 9927 14911 9953
rect 14937 9927 14943 9953
rect 12839 9921 12865 9927
rect 6511 9897 6537 9903
rect 6511 9865 6537 9871
rect 8807 9897 8833 9903
rect 8807 9865 8833 9871
rect 8975 9897 9001 9903
rect 8975 9865 9001 9871
rect 12615 9897 12641 9903
rect 12615 9865 12641 9871
rect 20007 9897 20033 9903
rect 20007 9865 20033 9871
rect 672 9813 20328 9830
rect 672 9787 2239 9813
rect 2265 9787 2291 9813
rect 2317 9787 2343 9813
rect 2369 9787 17599 9813
rect 17625 9787 17651 9813
rect 17677 9787 17703 9813
rect 17729 9787 20328 9813
rect 672 9770 20328 9787
rect 13175 9729 13201 9735
rect 13175 9697 13201 9703
rect 8359 9673 8385 9679
rect 12615 9673 12641 9679
rect 7177 9647 7183 9673
rect 7209 9647 7215 9673
rect 10817 9647 10823 9673
rect 10849 9647 10855 9673
rect 8359 9641 8385 9647
rect 12615 9641 12641 9647
rect 13287 9673 13313 9679
rect 13287 9641 13313 9647
rect 8807 9617 8833 9623
rect 10599 9617 10625 9623
rect 7345 9591 7351 9617
rect 7377 9591 7383 9617
rect 9361 9591 9367 9617
rect 9393 9591 9399 9617
rect 9753 9591 9759 9617
rect 9785 9591 9791 9617
rect 9977 9591 9983 9617
rect 10009 9591 10015 9617
rect 8807 9585 8833 9591
rect 10599 9585 10625 9591
rect 11271 9617 11297 9623
rect 11775 9617 11801 9623
rect 11545 9591 11551 9617
rect 11577 9591 11583 9617
rect 11271 9585 11297 9591
rect 11775 9585 11801 9591
rect 13399 9617 13425 9623
rect 13399 9585 13425 9591
rect 9479 9561 9505 9567
rect 7289 9535 7295 9561
rect 7321 9535 7327 9561
rect 8633 9535 8639 9561
rect 8665 9535 8671 9561
rect 9137 9535 9143 9561
rect 9169 9535 9175 9561
rect 9479 9529 9505 9535
rect 10879 9561 10905 9567
rect 10879 9529 10905 9535
rect 11327 9561 11353 9567
rect 11327 9529 11353 9535
rect 11999 9561 12025 9567
rect 11999 9529 12025 9535
rect 14295 9561 14321 9567
rect 14295 9529 14321 9535
rect 7015 9505 7041 9511
rect 7015 9473 7041 9479
rect 7463 9505 7489 9511
rect 7463 9473 7489 9479
rect 7575 9505 7601 9511
rect 8135 9505 8161 9511
rect 7961 9479 7967 9505
rect 7993 9479 7999 9505
rect 7575 9473 7601 9479
rect 8135 9473 8161 9479
rect 8975 9505 9001 9511
rect 8975 9473 9001 9479
rect 10039 9505 10065 9511
rect 10039 9473 10065 9479
rect 10767 9505 10793 9511
rect 10767 9473 10793 9479
rect 11383 9505 11409 9511
rect 11383 9473 11409 9479
rect 12447 9505 12473 9511
rect 12447 9473 12473 9479
rect 13511 9505 13537 9511
rect 13511 9473 13537 9479
rect 13567 9505 13593 9511
rect 13567 9473 13593 9479
rect 13623 9505 13649 9511
rect 13623 9473 13649 9479
rect 14239 9505 14265 9511
rect 14239 9473 14265 9479
rect 672 9421 20328 9438
rect 672 9395 9919 9421
rect 9945 9395 9971 9421
rect 9997 9395 10023 9421
rect 10049 9395 20328 9421
rect 672 9378 20328 9395
rect 7575 9337 7601 9343
rect 7575 9305 7601 9311
rect 7687 9337 7713 9343
rect 7687 9305 7713 9311
rect 7799 9337 7825 9343
rect 7799 9305 7825 9311
rect 11103 9337 11129 9343
rect 11103 9305 11129 9311
rect 11383 9337 11409 9343
rect 11383 9305 11409 9311
rect 12111 9337 12137 9343
rect 12111 9305 12137 9311
rect 13007 9337 13033 9343
rect 13007 9305 13033 9311
rect 8863 9281 8889 9287
rect 8863 9249 8889 9255
rect 10207 9281 10233 9287
rect 10207 9249 10233 9255
rect 11047 9281 11073 9287
rect 11047 9249 11073 9255
rect 11439 9281 11465 9287
rect 12783 9281 12809 9287
rect 11937 9255 11943 9281
rect 11969 9255 11975 9281
rect 11439 9249 11465 9255
rect 12783 9249 12809 9255
rect 12951 9281 12977 9287
rect 13729 9255 13735 9281
rect 13761 9255 13767 9281
rect 12951 9249 12977 9255
rect 7239 9225 7265 9231
rect 2137 9199 2143 9225
rect 2169 9199 2175 9225
rect 6505 9199 6511 9225
rect 6537 9199 6543 9225
rect 6897 9199 6903 9225
rect 6929 9199 6935 9225
rect 7239 9193 7265 9199
rect 8695 9225 8721 9231
rect 8695 9193 8721 9199
rect 9143 9225 9169 9231
rect 9143 9193 9169 9199
rect 9423 9225 9449 9231
rect 9423 9193 9449 9199
rect 9927 9225 9953 9231
rect 9927 9193 9953 9199
rect 11215 9225 11241 9231
rect 11215 9193 11241 9199
rect 11271 9225 11297 9231
rect 12609 9199 12615 9225
rect 12641 9199 12647 9225
rect 13393 9199 13399 9225
rect 13425 9199 13431 9225
rect 11271 9193 11297 9199
rect 7351 9169 7377 9175
rect 5441 9143 5447 9169
rect 5473 9143 5479 9169
rect 7351 9137 7377 9143
rect 7631 9169 7657 9175
rect 7631 9137 7657 9143
rect 8359 9169 8385 9175
rect 8359 9137 8385 9143
rect 12335 9169 12361 9175
rect 14793 9143 14799 9169
rect 14825 9143 14831 9169
rect 12335 9137 12361 9143
rect 967 9113 993 9119
rect 8415 9113 8441 9119
rect 7065 9087 7071 9113
rect 7097 9087 7103 9113
rect 967 9081 993 9087
rect 8415 9081 8441 9087
rect 12615 9113 12641 9119
rect 12615 9081 12641 9087
rect 13007 9113 13033 9119
rect 13007 9081 13033 9087
rect 672 9029 20328 9046
rect 672 9003 2239 9029
rect 2265 9003 2291 9029
rect 2317 9003 2343 9029
rect 2369 9003 17599 9029
rect 17625 9003 17651 9029
rect 17677 9003 17703 9029
rect 17729 9003 20328 9029
rect 672 8986 20328 9003
rect 7239 8945 7265 8951
rect 7239 8913 7265 8919
rect 11047 8945 11073 8951
rect 11047 8913 11073 8919
rect 11159 8945 11185 8951
rect 11159 8913 11185 8919
rect 12167 8945 12193 8951
rect 12167 8913 12193 8919
rect 12223 8945 12249 8951
rect 12223 8913 12249 8919
rect 967 8889 993 8895
rect 967 8857 993 8863
rect 7519 8889 7545 8895
rect 7519 8857 7545 8863
rect 10935 8889 10961 8895
rect 20007 8889 20033 8895
rect 12665 8863 12671 8889
rect 12697 8863 12703 8889
rect 13225 8863 13231 8889
rect 13257 8863 13263 8889
rect 14289 8863 14295 8889
rect 14321 8863 14327 8889
rect 10935 8857 10961 8863
rect 20007 8857 20033 8863
rect 6343 8833 6369 8839
rect 2137 8807 2143 8833
rect 2169 8807 2175 8833
rect 6343 8801 6369 8807
rect 7015 8833 7041 8839
rect 7015 8801 7041 8807
rect 7295 8833 7321 8839
rect 7295 8801 7321 8807
rect 10823 8833 10849 8839
rect 10823 8801 10849 8807
rect 11719 8833 11745 8839
rect 11719 8801 11745 8807
rect 12055 8833 12081 8839
rect 14631 8833 14657 8839
rect 12497 8807 12503 8833
rect 12529 8807 12535 8833
rect 12833 8807 12839 8833
rect 12865 8807 12871 8833
rect 18825 8807 18831 8833
rect 18857 8807 18863 8833
rect 12055 8801 12081 8807
rect 14631 8801 14657 8807
rect 6175 8777 6201 8783
rect 7239 8777 7265 8783
rect 6841 8751 6847 8777
rect 6873 8751 6879 8777
rect 6175 8745 6201 8751
rect 7239 8745 7265 8751
rect 12615 8777 12641 8783
rect 12615 8745 12641 8751
rect 7463 8721 7489 8727
rect 7463 8689 7489 8695
rect 10711 8721 10737 8727
rect 10711 8689 10737 8695
rect 10767 8721 10793 8727
rect 10767 8689 10793 8695
rect 11775 8721 11801 8727
rect 11775 8689 11801 8695
rect 11831 8721 11857 8727
rect 11831 8689 11857 8695
rect 12391 8721 12417 8727
rect 12391 8689 12417 8695
rect 672 8637 20328 8654
rect 672 8611 9919 8637
rect 9945 8611 9971 8637
rect 9997 8611 10023 8637
rect 10049 8611 20328 8637
rect 672 8594 20328 8611
rect 8751 8553 8777 8559
rect 8751 8521 8777 8527
rect 9815 8553 9841 8559
rect 9815 8521 9841 8527
rect 11999 8553 12025 8559
rect 11999 8521 12025 8527
rect 13903 8553 13929 8559
rect 13903 8521 13929 8527
rect 9647 8497 9673 8503
rect 10599 8497 10625 8503
rect 12727 8497 12753 8503
rect 7345 8471 7351 8497
rect 7377 8471 7383 8497
rect 9977 8471 9983 8497
rect 10009 8471 10015 8497
rect 11825 8471 11831 8497
rect 11857 8471 11863 8497
rect 9647 8465 9673 8471
rect 10599 8465 10625 8471
rect 12727 8465 12753 8471
rect 13959 8497 13985 8503
rect 13959 8465 13985 8471
rect 9479 8441 9505 8447
rect 6953 8415 6959 8441
rect 6985 8415 6991 8441
rect 9249 8415 9255 8441
rect 9281 8415 9287 8441
rect 9479 8409 9505 8415
rect 12615 8441 12641 8447
rect 12833 8415 12839 8441
rect 12865 8415 12871 8441
rect 12945 8415 12951 8441
rect 12977 8415 12983 8441
rect 18825 8415 18831 8441
rect 18857 8415 18863 8441
rect 12615 8409 12641 8415
rect 9591 8385 9617 8391
rect 8409 8359 8415 8385
rect 8441 8359 8447 8385
rect 9591 8353 9617 8359
rect 10487 8385 10513 8391
rect 12671 8385 12697 8391
rect 10649 8359 10655 8385
rect 10681 8359 10687 8385
rect 10487 8353 10513 8359
rect 12671 8353 12697 8359
rect 9423 8329 9449 8335
rect 9423 8297 9449 8303
rect 20007 8329 20033 8335
rect 20007 8297 20033 8303
rect 672 8245 20328 8262
rect 672 8219 2239 8245
rect 2265 8219 2291 8245
rect 2317 8219 2343 8245
rect 2369 8219 17599 8245
rect 17625 8219 17651 8245
rect 17677 8219 17703 8245
rect 17729 8219 20328 8245
rect 672 8202 20328 8219
rect 9535 8161 9561 8167
rect 9535 8129 9561 8135
rect 9703 8161 9729 8167
rect 9703 8129 9729 8135
rect 13623 8105 13649 8111
rect 12329 8079 12335 8105
rect 12361 8079 12367 8105
rect 13393 8079 13399 8105
rect 13425 8079 13431 8105
rect 13623 8073 13649 8079
rect 11937 8023 11943 8049
rect 11969 8023 11975 8049
rect 9591 7937 9617 7943
rect 9591 7905 9617 7911
rect 672 7853 20328 7870
rect 672 7827 9919 7853
rect 9945 7827 9971 7853
rect 9997 7827 10023 7853
rect 10049 7827 20328 7853
rect 672 7810 20328 7827
rect 12615 7769 12641 7775
rect 12615 7737 12641 7743
rect 12839 7769 12865 7775
rect 12839 7737 12865 7743
rect 13063 7769 13089 7775
rect 13063 7737 13089 7743
rect 11327 7713 11353 7719
rect 10761 7687 10767 7713
rect 10793 7687 10799 7713
rect 11327 7681 11353 7687
rect 11439 7713 11465 7719
rect 11439 7681 11465 7687
rect 12727 7657 12753 7663
rect 11153 7631 11159 7657
rect 11185 7631 11191 7657
rect 12727 7625 12753 7631
rect 11383 7601 11409 7607
rect 9697 7575 9703 7601
rect 9729 7575 9735 7601
rect 11383 7569 11409 7575
rect 11719 7601 11745 7607
rect 11719 7569 11745 7575
rect 12671 7601 12697 7607
rect 12671 7569 12697 7575
rect 13119 7601 13145 7607
rect 13119 7569 13145 7575
rect 672 7461 20328 7478
rect 672 7435 2239 7461
rect 2265 7435 2291 7461
rect 2317 7435 2343 7461
rect 2369 7435 17599 7461
rect 17625 7435 17651 7461
rect 17677 7435 17703 7461
rect 17729 7435 20328 7461
rect 672 7418 20328 7435
rect 10879 7377 10905 7383
rect 10879 7345 10905 7351
rect 13511 7321 13537 7327
rect 8689 7295 8695 7321
rect 8721 7295 8727 7321
rect 9753 7295 9759 7321
rect 9785 7295 9791 7321
rect 10705 7295 10711 7321
rect 10737 7295 10743 7321
rect 12217 7295 12223 7321
rect 12249 7295 12255 7321
rect 13281 7295 13287 7321
rect 13313 7295 13319 7321
rect 13511 7289 13537 7295
rect 9983 7265 10009 7271
rect 8353 7239 8359 7265
rect 8385 7239 8391 7265
rect 11825 7239 11831 7265
rect 11857 7239 11863 7265
rect 9983 7233 10009 7239
rect 10767 7209 10793 7215
rect 10767 7177 10793 7183
rect 672 7069 20328 7086
rect 672 7043 9919 7069
rect 9945 7043 9971 7069
rect 9997 7043 10023 7069
rect 10049 7043 20328 7069
rect 672 7026 20328 7043
rect 12839 6985 12865 6991
rect 12839 6953 12865 6959
rect 10201 6903 10207 6929
rect 10233 6903 10239 6929
rect 11495 6873 11521 6879
rect 9865 6847 9871 6873
rect 9897 6847 9903 6873
rect 11495 6841 11521 6847
rect 12895 6817 12921 6823
rect 11265 6791 11271 6817
rect 11297 6791 11303 6817
rect 12895 6785 12921 6791
rect 672 6677 20328 6694
rect 672 6651 2239 6677
rect 2265 6651 2291 6677
rect 2317 6651 2343 6677
rect 2369 6651 17599 6677
rect 17625 6651 17651 6677
rect 17677 6651 17703 6677
rect 17729 6651 20328 6677
rect 672 6634 20328 6651
rect 672 6285 20328 6302
rect 672 6259 9919 6285
rect 9945 6259 9971 6285
rect 9997 6259 10023 6285
rect 10049 6259 20328 6285
rect 672 6242 20328 6259
rect 672 5893 20328 5910
rect 672 5867 2239 5893
rect 2265 5867 2291 5893
rect 2317 5867 2343 5893
rect 2369 5867 17599 5893
rect 17625 5867 17651 5893
rect 17677 5867 17703 5893
rect 17729 5867 20328 5893
rect 672 5850 20328 5867
rect 672 5501 20328 5518
rect 672 5475 9919 5501
rect 9945 5475 9971 5501
rect 9997 5475 10023 5501
rect 10049 5475 20328 5501
rect 672 5458 20328 5475
rect 672 5109 20328 5126
rect 672 5083 2239 5109
rect 2265 5083 2291 5109
rect 2317 5083 2343 5109
rect 2369 5083 17599 5109
rect 17625 5083 17651 5109
rect 17677 5083 17703 5109
rect 17729 5083 20328 5109
rect 672 5066 20328 5083
rect 672 4717 20328 4734
rect 672 4691 9919 4717
rect 9945 4691 9971 4717
rect 9997 4691 10023 4717
rect 10049 4691 20328 4717
rect 672 4674 20328 4691
rect 672 4325 20328 4342
rect 672 4299 2239 4325
rect 2265 4299 2291 4325
rect 2317 4299 2343 4325
rect 2369 4299 17599 4325
rect 17625 4299 17651 4325
rect 17677 4299 17703 4325
rect 17729 4299 20328 4325
rect 672 4282 20328 4299
rect 672 3933 20328 3950
rect 672 3907 9919 3933
rect 9945 3907 9971 3933
rect 9997 3907 10023 3933
rect 10049 3907 20328 3933
rect 672 3890 20328 3907
rect 672 3541 20328 3558
rect 672 3515 2239 3541
rect 2265 3515 2291 3541
rect 2317 3515 2343 3541
rect 2369 3515 17599 3541
rect 17625 3515 17651 3541
rect 17677 3515 17703 3541
rect 17729 3515 20328 3541
rect 672 3498 20328 3515
rect 672 3149 20328 3166
rect 672 3123 9919 3149
rect 9945 3123 9971 3149
rect 9997 3123 10023 3149
rect 10049 3123 20328 3149
rect 672 3106 20328 3123
rect 672 2757 20328 2774
rect 672 2731 2239 2757
rect 2265 2731 2291 2757
rect 2317 2731 2343 2757
rect 2369 2731 17599 2757
rect 17625 2731 17651 2757
rect 17677 2731 17703 2757
rect 17729 2731 20328 2757
rect 672 2714 20328 2731
rect 672 2365 20328 2382
rect 672 2339 9919 2365
rect 9945 2339 9971 2365
rect 9997 2339 10023 2365
rect 10049 2339 20328 2365
rect 672 2322 20328 2339
rect 9417 2143 9423 2169
rect 9449 2143 9455 2169
rect 10929 2143 10935 2169
rect 10961 2143 10967 2169
rect 13225 2143 13231 2169
rect 13257 2143 13263 2169
rect 9927 2057 9953 2063
rect 9927 2025 9953 2031
rect 11383 2057 11409 2063
rect 11383 2025 11409 2031
rect 13735 2057 13761 2063
rect 13735 2025 13761 2031
rect 672 1973 20328 1990
rect 672 1947 2239 1973
rect 2265 1947 2291 1973
rect 2317 1947 2343 1973
rect 2369 1947 17599 1973
rect 17625 1947 17651 1973
rect 17677 1947 17703 1973
rect 17729 1947 20328 1973
rect 672 1930 20328 1947
rect 11937 1751 11943 1777
rect 11969 1751 11975 1777
rect 11097 1695 11103 1721
rect 11129 1695 11135 1721
rect 9199 1665 9225 1671
rect 9199 1633 9225 1639
rect 672 1581 20328 1598
rect 672 1555 9919 1581
rect 9945 1555 9971 1581
rect 9997 1555 10023 1581
rect 10049 1555 20328 1581
rect 672 1538 20328 1555
<< via1 >>
rect 2239 19195 2265 19221
rect 2291 19195 2317 19221
rect 2343 19195 2369 19221
rect 17599 19195 17625 19221
rect 17651 19195 17677 19221
rect 17703 19195 17729 19221
rect 9031 19111 9057 19137
rect 10879 19111 10905 19137
rect 12783 19111 12809 19137
rect 14687 19111 14713 19137
rect 8527 18999 8553 19025
rect 10375 18999 10401 19025
rect 12279 18999 12305 19025
rect 14295 18999 14321 19025
rect 9919 18803 9945 18829
rect 9971 18803 9997 18829
rect 10023 18803 10049 18829
rect 10039 18719 10065 18745
rect 12615 18719 12641 18745
rect 13399 18719 13425 18745
rect 9535 18607 9561 18633
rect 12895 18607 12921 18633
rect 2239 18411 2265 18437
rect 2291 18411 2317 18437
rect 2343 18411 2369 18437
rect 17599 18411 17625 18437
rect 17651 18411 17677 18437
rect 17703 18411 17729 18437
rect 9919 18019 9945 18045
rect 9971 18019 9997 18045
rect 10023 18019 10049 18045
rect 2239 17627 2265 17653
rect 2291 17627 2317 17653
rect 2343 17627 2369 17653
rect 17599 17627 17625 17653
rect 17651 17627 17677 17653
rect 17703 17627 17729 17653
rect 9919 17235 9945 17261
rect 9971 17235 9997 17261
rect 10023 17235 10049 17261
rect 2239 16843 2265 16869
rect 2291 16843 2317 16869
rect 2343 16843 2369 16869
rect 17599 16843 17625 16869
rect 17651 16843 17677 16869
rect 17703 16843 17729 16869
rect 9919 16451 9945 16477
rect 9971 16451 9997 16477
rect 10023 16451 10049 16477
rect 2239 16059 2265 16085
rect 2291 16059 2317 16085
rect 2343 16059 2369 16085
rect 17599 16059 17625 16085
rect 17651 16059 17677 16085
rect 17703 16059 17729 16085
rect 9919 15667 9945 15693
rect 9971 15667 9997 15693
rect 10023 15667 10049 15693
rect 2239 15275 2265 15301
rect 2291 15275 2317 15301
rect 2343 15275 2369 15301
rect 17599 15275 17625 15301
rect 17651 15275 17677 15301
rect 17703 15275 17729 15301
rect 9919 14883 9945 14909
rect 9971 14883 9997 14909
rect 10023 14883 10049 14909
rect 2239 14491 2265 14517
rect 2291 14491 2317 14517
rect 2343 14491 2369 14517
rect 17599 14491 17625 14517
rect 17651 14491 17677 14517
rect 17703 14491 17729 14517
rect 9535 14351 9561 14377
rect 12111 14351 12137 14377
rect 8135 14295 8161 14321
rect 9759 14295 9785 14321
rect 10711 14295 10737 14321
rect 11047 14295 11073 14321
rect 12335 14295 12361 14321
rect 8471 14239 8497 14265
rect 9919 14099 9945 14125
rect 9971 14099 9997 14125
rect 10023 14099 10049 14125
rect 8415 14015 8441 14041
rect 10879 14015 10905 14041
rect 11271 14015 11297 14041
rect 10767 13959 10793 13985
rect 11159 13959 11185 13985
rect 8919 13903 8945 13929
rect 10711 13903 10737 13929
rect 11327 13903 11353 13929
rect 9255 13847 9281 13873
rect 10319 13847 10345 13873
rect 2239 13707 2265 13733
rect 2291 13707 2317 13733
rect 2343 13707 2369 13733
rect 17599 13707 17625 13733
rect 17651 13707 17677 13733
rect 17703 13707 17729 13733
rect 9647 13623 9673 13649
rect 8471 13567 8497 13593
rect 8695 13567 8721 13593
rect 13231 13567 13257 13593
rect 7071 13511 7097 13537
rect 9031 13511 9057 13537
rect 9311 13511 9337 13537
rect 9479 13511 9505 13537
rect 11831 13511 11857 13537
rect 7407 13455 7433 13481
rect 9143 13455 9169 13481
rect 9199 13455 9225 13481
rect 9423 13455 9449 13481
rect 9703 13455 9729 13481
rect 12167 13455 12193 13481
rect 13455 13455 13481 13481
rect 9919 13315 9945 13341
rect 9971 13315 9997 13341
rect 10023 13315 10049 13341
rect 7463 13231 7489 13257
rect 7911 13231 7937 13257
rect 8807 13231 8833 13257
rect 9367 13231 9393 13257
rect 9927 13231 9953 13257
rect 9983 13231 10009 13257
rect 12167 13231 12193 13257
rect 7183 13175 7209 13201
rect 8695 13175 8721 13201
rect 12839 13175 12865 13201
rect 2143 13119 2169 13145
rect 6959 13119 6985 13145
rect 7127 13119 7153 13145
rect 8919 13119 8945 13145
rect 9031 13119 9057 13145
rect 9535 13119 9561 13145
rect 9759 13119 9785 13145
rect 9871 13119 9897 13145
rect 10095 13119 10121 13145
rect 11383 13119 11409 13145
rect 11439 13119 11465 13145
rect 11663 13119 11689 13145
rect 11775 13119 11801 13145
rect 11887 13119 11913 13145
rect 12111 13119 12137 13145
rect 12223 13119 12249 13145
rect 12783 13119 12809 13145
rect 18831 13119 18857 13145
rect 5503 13063 5529 13089
rect 6567 13063 6593 13089
rect 7967 13063 7993 13089
rect 8863 13063 8889 13089
rect 11551 13063 11577 13089
rect 11999 13063 12025 13089
rect 19951 13063 19977 13089
rect 967 13007 993 13033
rect 7183 13007 7209 13033
rect 2239 12923 2265 12949
rect 2291 12923 2317 12949
rect 2343 12923 2369 12949
rect 17599 12923 17625 12949
rect 17651 12923 17677 12949
rect 17703 12923 17729 12949
rect 10935 12839 10961 12865
rect 11719 12783 11745 12809
rect 12783 12783 12809 12809
rect 20007 12783 20033 12809
rect 6903 12727 6929 12753
rect 9759 12727 9785 12753
rect 10655 12727 10681 12753
rect 10767 12727 10793 12753
rect 11383 12727 11409 12753
rect 14631 12727 14657 12753
rect 18831 12727 18857 12753
rect 6735 12671 6761 12697
rect 6791 12671 6817 12697
rect 9871 12671 9897 12697
rect 13903 12671 13929 12697
rect 14743 12671 14769 12697
rect 7127 12615 7153 12641
rect 13007 12615 13033 12641
rect 13231 12615 13257 12641
rect 13847 12615 13873 12641
rect 9919 12531 9945 12557
rect 9971 12531 9997 12557
rect 10023 12531 10049 12557
rect 6511 12447 6537 12473
rect 11999 12447 12025 12473
rect 13063 12447 13089 12473
rect 13119 12447 13145 12473
rect 9479 12391 9505 12417
rect 9703 12391 9729 12417
rect 10039 12391 10065 12417
rect 11663 12391 11689 12417
rect 12111 12391 12137 12417
rect 13791 12391 13817 12417
rect 9311 12335 9337 12361
rect 11551 12335 11577 12361
rect 11943 12335 11969 12361
rect 12223 12335 12249 12361
rect 12951 12335 12977 12361
rect 13007 12335 13033 12361
rect 13231 12335 13257 12361
rect 13399 12335 13425 12361
rect 9983 12279 10009 12305
rect 14855 12279 14881 12305
rect 9647 12223 9673 12249
rect 9815 12223 9841 12249
rect 10151 12223 10177 12249
rect 2239 12139 2265 12165
rect 2291 12139 2317 12165
rect 2343 12139 2369 12165
rect 17599 12139 17625 12165
rect 17651 12139 17677 12165
rect 17703 12139 17729 12165
rect 10431 12055 10457 12081
rect 967 11999 993 12025
rect 4943 11999 4969 12025
rect 7071 11999 7097 12025
rect 8695 11999 8721 12025
rect 8919 11999 8945 12025
rect 11607 11999 11633 12025
rect 20007 11999 20033 12025
rect 2143 11943 2169 11969
rect 6399 11943 6425 11969
rect 6847 11943 6873 11969
rect 7239 11943 7265 11969
rect 9423 11943 9449 11969
rect 10095 11943 10121 11969
rect 10711 11943 10737 11969
rect 13007 11943 13033 11969
rect 13847 11943 13873 11969
rect 18831 11943 18857 11969
rect 6007 11887 6033 11913
rect 6791 11887 6817 11913
rect 7631 11887 7657 11913
rect 9255 11887 9281 11913
rect 9535 11887 9561 11913
rect 9815 11887 9841 11913
rect 12671 11887 12697 11913
rect 13903 11887 13929 11913
rect 6679 11831 6705 11857
rect 9087 11831 9113 11857
rect 9647 11831 9673 11857
rect 10263 11831 10289 11857
rect 10375 11831 10401 11857
rect 10823 11831 10849 11857
rect 13287 11831 13313 11857
rect 14015 11831 14041 11857
rect 9919 11747 9945 11773
rect 9971 11747 9997 11773
rect 10023 11747 10049 11773
rect 6175 11663 6201 11689
rect 9479 11663 9505 11689
rect 12671 11663 12697 11689
rect 13063 11663 13089 11689
rect 6287 11607 6313 11633
rect 6343 11607 6369 11633
rect 7743 11607 7769 11633
rect 8023 11607 8049 11633
rect 9255 11607 9281 11633
rect 9311 11607 9337 11633
rect 11887 11607 11913 11633
rect 8135 11551 8161 11577
rect 9031 11551 9057 11577
rect 9143 11551 9169 11577
rect 10039 11551 10065 11577
rect 10655 11551 10681 11577
rect 11047 11551 11073 11577
rect 11663 11551 11689 11577
rect 12839 11551 12865 11577
rect 12951 11551 12977 11577
rect 13287 11551 13313 11577
rect 7687 11495 7713 11521
rect 7855 11495 7881 11521
rect 9759 11495 9785 11521
rect 9927 11495 9953 11521
rect 10879 11495 10905 11521
rect 11327 11495 11353 11521
rect 11719 11495 11745 11521
rect 12895 11495 12921 11521
rect 13679 11495 13705 11521
rect 14743 11495 14769 11521
rect 8975 11439 9001 11465
rect 10207 11439 10233 11465
rect 11831 11439 11857 11465
rect 2239 11355 2265 11381
rect 2291 11355 2317 11381
rect 2343 11355 2369 11381
rect 17599 11355 17625 11381
rect 17651 11355 17677 11381
rect 17703 11355 17729 11381
rect 12727 11271 12753 11297
rect 967 11215 993 11241
rect 8919 11215 8945 11241
rect 11159 11215 11185 11241
rect 2143 11159 2169 11185
rect 7015 11159 7041 11185
rect 7127 11159 7153 11185
rect 9703 11159 9729 11185
rect 10935 11159 10961 11185
rect 12223 11159 12249 11185
rect 12447 11159 12473 11185
rect 12559 11159 12585 11185
rect 12951 11159 12977 11185
rect 7351 11103 7377 11129
rect 10991 11103 11017 11129
rect 11439 11103 11465 11129
rect 6959 11047 6985 11073
rect 7239 11047 7265 11073
rect 13063 11047 13089 11073
rect 9919 10963 9945 10989
rect 9971 10963 9997 10989
rect 10023 10963 10049 10989
rect 7743 10879 7769 10905
rect 12671 10879 12697 10905
rect 6735 10823 6761 10849
rect 7687 10823 7713 10849
rect 8975 10823 9001 10849
rect 2143 10767 2169 10793
rect 7127 10767 7153 10793
rect 7519 10767 7545 10793
rect 7799 10767 7825 10793
rect 7911 10767 7937 10793
rect 8135 10767 8161 10793
rect 8247 10767 8273 10793
rect 8863 10767 8889 10793
rect 9255 10767 9281 10793
rect 9591 10767 9617 10793
rect 18831 10767 18857 10793
rect 5671 10711 5697 10737
rect 7351 10711 7377 10737
rect 8191 10711 8217 10737
rect 9143 10711 9169 10737
rect 11327 10711 11353 10737
rect 13287 10711 13313 10737
rect 14575 10711 14601 10737
rect 967 10655 993 10681
rect 9423 10655 9449 10681
rect 14519 10655 14545 10681
rect 20007 10655 20033 10681
rect 2239 10571 2265 10597
rect 2291 10571 2317 10597
rect 2343 10571 2369 10597
rect 17599 10571 17625 10597
rect 17651 10571 17677 10597
rect 17703 10571 17729 10597
rect 6063 10487 6089 10513
rect 9199 10487 9225 10513
rect 7127 10431 7153 10457
rect 8191 10431 8217 10457
rect 10711 10431 10737 10457
rect 11103 10431 11129 10457
rect 6119 10375 6145 10401
rect 6343 10375 6369 10401
rect 6791 10375 6817 10401
rect 8359 10375 8385 10401
rect 8751 10375 8777 10401
rect 9479 10375 9505 10401
rect 9647 10375 9673 10401
rect 10095 10375 10121 10401
rect 10319 10375 10345 10401
rect 10823 10375 10849 10401
rect 11047 10375 11073 10401
rect 11327 10375 11353 10401
rect 8863 10319 8889 10345
rect 9031 10319 9057 10345
rect 10263 10319 10289 10345
rect 13343 10319 13369 10345
rect 6063 10263 6089 10289
rect 8527 10263 8553 10289
rect 9143 10263 9169 10289
rect 9367 10263 9393 10289
rect 11159 10263 11185 10289
rect 20119 10263 20145 10289
rect 9919 10179 9945 10205
rect 9971 10179 9997 10205
rect 10023 10179 10049 10205
rect 7855 10095 7881 10121
rect 8303 10095 8329 10121
rect 11383 10095 11409 10121
rect 6455 10039 6481 10065
rect 6511 10039 6537 10065
rect 6791 10039 6817 10065
rect 7463 10039 7489 10065
rect 7743 10039 7769 10065
rect 8247 10039 8273 10065
rect 9591 10039 9617 10065
rect 10095 10039 10121 10065
rect 11719 10039 11745 10065
rect 11887 10039 11913 10065
rect 12279 10039 12305 10065
rect 12391 10039 12417 10065
rect 13063 10039 13089 10065
rect 6287 9983 6313 10009
rect 7911 9983 7937 10009
rect 9143 9983 9169 10009
rect 9311 9983 9337 10009
rect 10151 9983 10177 10009
rect 11271 9983 11297 10009
rect 11607 9983 11633 10009
rect 12223 9983 12249 10009
rect 12727 9983 12753 10009
rect 12951 9983 12977 10009
rect 13455 9983 13481 10009
rect 18831 9983 18857 10009
rect 4831 9927 4857 9953
rect 5895 9927 5921 9953
rect 8751 9927 8777 9953
rect 9087 9927 9113 9953
rect 9367 9927 9393 9953
rect 11327 9927 11353 9953
rect 12839 9927 12865 9953
rect 13007 9927 13033 9953
rect 13847 9927 13873 9953
rect 14911 9927 14937 9953
rect 6511 9871 6537 9897
rect 8807 9871 8833 9897
rect 8975 9871 9001 9897
rect 12615 9871 12641 9897
rect 20007 9871 20033 9897
rect 2239 9787 2265 9813
rect 2291 9787 2317 9813
rect 2343 9787 2369 9813
rect 17599 9787 17625 9813
rect 17651 9787 17677 9813
rect 17703 9787 17729 9813
rect 13175 9703 13201 9729
rect 7183 9647 7209 9673
rect 8359 9647 8385 9673
rect 10823 9647 10849 9673
rect 12615 9647 12641 9673
rect 13287 9647 13313 9673
rect 7351 9591 7377 9617
rect 8807 9591 8833 9617
rect 9367 9591 9393 9617
rect 9759 9591 9785 9617
rect 9983 9591 10009 9617
rect 10599 9591 10625 9617
rect 11271 9591 11297 9617
rect 11551 9591 11577 9617
rect 11775 9591 11801 9617
rect 13399 9591 13425 9617
rect 7295 9535 7321 9561
rect 8639 9535 8665 9561
rect 9143 9535 9169 9561
rect 9479 9535 9505 9561
rect 10879 9535 10905 9561
rect 11327 9535 11353 9561
rect 11999 9535 12025 9561
rect 14295 9535 14321 9561
rect 7015 9479 7041 9505
rect 7463 9479 7489 9505
rect 7575 9479 7601 9505
rect 7967 9479 7993 9505
rect 8135 9479 8161 9505
rect 8975 9479 9001 9505
rect 10039 9479 10065 9505
rect 10767 9479 10793 9505
rect 11383 9479 11409 9505
rect 12447 9479 12473 9505
rect 13511 9479 13537 9505
rect 13567 9479 13593 9505
rect 13623 9479 13649 9505
rect 14239 9479 14265 9505
rect 9919 9395 9945 9421
rect 9971 9395 9997 9421
rect 10023 9395 10049 9421
rect 7575 9311 7601 9337
rect 7687 9311 7713 9337
rect 7799 9311 7825 9337
rect 11103 9311 11129 9337
rect 11383 9311 11409 9337
rect 12111 9311 12137 9337
rect 13007 9311 13033 9337
rect 8863 9255 8889 9281
rect 10207 9255 10233 9281
rect 11047 9255 11073 9281
rect 11439 9255 11465 9281
rect 11943 9255 11969 9281
rect 12783 9255 12809 9281
rect 12951 9255 12977 9281
rect 13735 9255 13761 9281
rect 2143 9199 2169 9225
rect 6511 9199 6537 9225
rect 6903 9199 6929 9225
rect 7239 9199 7265 9225
rect 8695 9199 8721 9225
rect 9143 9199 9169 9225
rect 9423 9199 9449 9225
rect 9927 9199 9953 9225
rect 11215 9199 11241 9225
rect 11271 9199 11297 9225
rect 12615 9199 12641 9225
rect 13399 9199 13425 9225
rect 5447 9143 5473 9169
rect 7351 9143 7377 9169
rect 7631 9143 7657 9169
rect 8359 9143 8385 9169
rect 12335 9143 12361 9169
rect 14799 9143 14825 9169
rect 967 9087 993 9113
rect 7071 9087 7097 9113
rect 8415 9087 8441 9113
rect 12615 9087 12641 9113
rect 13007 9087 13033 9113
rect 2239 9003 2265 9029
rect 2291 9003 2317 9029
rect 2343 9003 2369 9029
rect 17599 9003 17625 9029
rect 17651 9003 17677 9029
rect 17703 9003 17729 9029
rect 7239 8919 7265 8945
rect 11047 8919 11073 8945
rect 11159 8919 11185 8945
rect 12167 8919 12193 8945
rect 12223 8919 12249 8945
rect 967 8863 993 8889
rect 7519 8863 7545 8889
rect 10935 8863 10961 8889
rect 12671 8863 12697 8889
rect 13231 8863 13257 8889
rect 14295 8863 14321 8889
rect 20007 8863 20033 8889
rect 2143 8807 2169 8833
rect 6343 8807 6369 8833
rect 7015 8807 7041 8833
rect 7295 8807 7321 8833
rect 10823 8807 10849 8833
rect 11719 8807 11745 8833
rect 12055 8807 12081 8833
rect 12503 8807 12529 8833
rect 12839 8807 12865 8833
rect 14631 8807 14657 8833
rect 18831 8807 18857 8833
rect 6175 8751 6201 8777
rect 6847 8751 6873 8777
rect 7239 8751 7265 8777
rect 12615 8751 12641 8777
rect 7463 8695 7489 8721
rect 10711 8695 10737 8721
rect 10767 8695 10793 8721
rect 11775 8695 11801 8721
rect 11831 8695 11857 8721
rect 12391 8695 12417 8721
rect 9919 8611 9945 8637
rect 9971 8611 9997 8637
rect 10023 8611 10049 8637
rect 8751 8527 8777 8553
rect 9815 8527 9841 8553
rect 11999 8527 12025 8553
rect 13903 8527 13929 8553
rect 7351 8471 7377 8497
rect 9647 8471 9673 8497
rect 9983 8471 10009 8497
rect 10599 8471 10625 8497
rect 11831 8471 11857 8497
rect 12727 8471 12753 8497
rect 13959 8471 13985 8497
rect 6959 8415 6985 8441
rect 9255 8415 9281 8441
rect 9479 8415 9505 8441
rect 12615 8415 12641 8441
rect 12839 8415 12865 8441
rect 12951 8415 12977 8441
rect 18831 8415 18857 8441
rect 8415 8359 8441 8385
rect 9591 8359 9617 8385
rect 10487 8359 10513 8385
rect 10655 8359 10681 8385
rect 12671 8359 12697 8385
rect 9423 8303 9449 8329
rect 20007 8303 20033 8329
rect 2239 8219 2265 8245
rect 2291 8219 2317 8245
rect 2343 8219 2369 8245
rect 17599 8219 17625 8245
rect 17651 8219 17677 8245
rect 17703 8219 17729 8245
rect 9535 8135 9561 8161
rect 9703 8135 9729 8161
rect 12335 8079 12361 8105
rect 13399 8079 13425 8105
rect 13623 8079 13649 8105
rect 11943 8023 11969 8049
rect 9591 7911 9617 7937
rect 9919 7827 9945 7853
rect 9971 7827 9997 7853
rect 10023 7827 10049 7853
rect 12615 7743 12641 7769
rect 12839 7743 12865 7769
rect 13063 7743 13089 7769
rect 10767 7687 10793 7713
rect 11327 7687 11353 7713
rect 11439 7687 11465 7713
rect 11159 7631 11185 7657
rect 12727 7631 12753 7657
rect 9703 7575 9729 7601
rect 11383 7575 11409 7601
rect 11719 7575 11745 7601
rect 12671 7575 12697 7601
rect 13119 7575 13145 7601
rect 2239 7435 2265 7461
rect 2291 7435 2317 7461
rect 2343 7435 2369 7461
rect 17599 7435 17625 7461
rect 17651 7435 17677 7461
rect 17703 7435 17729 7461
rect 10879 7351 10905 7377
rect 8695 7295 8721 7321
rect 9759 7295 9785 7321
rect 10711 7295 10737 7321
rect 12223 7295 12249 7321
rect 13287 7295 13313 7321
rect 13511 7295 13537 7321
rect 8359 7239 8385 7265
rect 9983 7239 10009 7265
rect 11831 7239 11857 7265
rect 10767 7183 10793 7209
rect 9919 7043 9945 7069
rect 9971 7043 9997 7069
rect 10023 7043 10049 7069
rect 12839 6959 12865 6985
rect 10207 6903 10233 6929
rect 9871 6847 9897 6873
rect 11495 6847 11521 6873
rect 11271 6791 11297 6817
rect 12895 6791 12921 6817
rect 2239 6651 2265 6677
rect 2291 6651 2317 6677
rect 2343 6651 2369 6677
rect 17599 6651 17625 6677
rect 17651 6651 17677 6677
rect 17703 6651 17729 6677
rect 9919 6259 9945 6285
rect 9971 6259 9997 6285
rect 10023 6259 10049 6285
rect 2239 5867 2265 5893
rect 2291 5867 2317 5893
rect 2343 5867 2369 5893
rect 17599 5867 17625 5893
rect 17651 5867 17677 5893
rect 17703 5867 17729 5893
rect 9919 5475 9945 5501
rect 9971 5475 9997 5501
rect 10023 5475 10049 5501
rect 2239 5083 2265 5109
rect 2291 5083 2317 5109
rect 2343 5083 2369 5109
rect 17599 5083 17625 5109
rect 17651 5083 17677 5109
rect 17703 5083 17729 5109
rect 9919 4691 9945 4717
rect 9971 4691 9997 4717
rect 10023 4691 10049 4717
rect 2239 4299 2265 4325
rect 2291 4299 2317 4325
rect 2343 4299 2369 4325
rect 17599 4299 17625 4325
rect 17651 4299 17677 4325
rect 17703 4299 17729 4325
rect 9919 3907 9945 3933
rect 9971 3907 9997 3933
rect 10023 3907 10049 3933
rect 2239 3515 2265 3541
rect 2291 3515 2317 3541
rect 2343 3515 2369 3541
rect 17599 3515 17625 3541
rect 17651 3515 17677 3541
rect 17703 3515 17729 3541
rect 9919 3123 9945 3149
rect 9971 3123 9997 3149
rect 10023 3123 10049 3149
rect 2239 2731 2265 2757
rect 2291 2731 2317 2757
rect 2343 2731 2369 2757
rect 17599 2731 17625 2757
rect 17651 2731 17677 2757
rect 17703 2731 17729 2757
rect 9919 2339 9945 2365
rect 9971 2339 9997 2365
rect 10023 2339 10049 2365
rect 9423 2143 9449 2169
rect 10935 2143 10961 2169
rect 13231 2143 13257 2169
rect 9927 2031 9953 2057
rect 11383 2031 11409 2057
rect 13735 2031 13761 2057
rect 2239 1947 2265 1973
rect 2291 1947 2317 1973
rect 2343 1947 2369 1973
rect 17599 1947 17625 1973
rect 17651 1947 17677 1973
rect 17703 1947 17729 1973
rect 11943 1751 11969 1777
rect 11103 1695 11129 1721
rect 9199 1639 9225 1665
rect 9919 1555 9945 1581
rect 9971 1555 9997 1581
rect 10023 1555 10049 1581
<< metal2 >>
rect 8400 20600 8456 21000
rect 9408 20600 9464 21000
rect 10080 20600 10136 21000
rect 11424 20600 11480 21000
rect 12432 20600 12488 21000
rect 12768 20600 12824 21000
rect 13104 20600 13160 21000
rect 2238 19222 2370 19227
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2238 19189 2370 19194
rect 8414 19138 8442 20600
rect 8414 19105 8442 19110
rect 9030 19138 9058 19143
rect 9030 19091 9058 19110
rect 8526 19025 8554 19031
rect 8526 18999 8527 19025
rect 8553 18999 8554 19025
rect 2238 18438 2370 18443
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2238 18405 2370 18410
rect 2238 17654 2370 17659
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2238 17621 2370 17626
rect 2238 16870 2370 16875
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2238 16837 2370 16842
rect 2238 16086 2370 16091
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2238 16053 2370 16058
rect 2238 15302 2370 15307
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2238 15269 2370 15274
rect 2238 14518 2370 14523
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2238 14485 2370 14490
rect 7630 14322 7658 14327
rect 7574 14294 7630 14322
rect 7574 14266 7602 14294
rect 7630 14289 7658 14294
rect 8134 14322 8162 14327
rect 8134 14275 8162 14294
rect 8414 14322 8442 14327
rect 7462 14238 7602 14266
rect 2086 14154 2114 14159
rect 966 13033 994 13039
rect 966 13007 967 13033
rect 993 13007 994 13033
rect 966 12810 994 13007
rect 966 12777 994 12782
rect 966 12025 994 12031
rect 966 11999 967 12025
rect 993 11999 994 12025
rect 966 11802 994 11999
rect 966 11769 994 11774
rect 966 11242 994 11247
rect 966 11195 994 11214
rect 2086 10794 2114 14126
rect 2238 13734 2370 13739
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2238 13701 2370 13706
rect 7462 13594 7490 14238
rect 8414 14041 8442 14294
rect 8470 14266 8498 14271
rect 8470 14219 8498 14238
rect 8414 14015 8415 14041
rect 8441 14015 8442 14041
rect 8414 14009 8442 14015
rect 7070 13566 7490 13594
rect 7070 13538 7098 13566
rect 7014 13537 7098 13538
rect 7014 13511 7071 13537
rect 7097 13511 7098 13537
rect 7014 13510 7098 13511
rect 2142 13146 2170 13151
rect 2142 13099 2170 13118
rect 5502 13146 5530 13151
rect 5502 13089 5530 13118
rect 6790 13146 6818 13151
rect 5502 13063 5503 13089
rect 5529 13063 5530 13089
rect 5502 13057 5530 13063
rect 6566 13089 6594 13095
rect 6566 13063 6567 13089
rect 6593 13063 6594 13089
rect 6566 13034 6594 13063
rect 6566 13001 6594 13006
rect 2238 12950 2370 12955
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2238 12917 2370 12922
rect 6734 12697 6762 12703
rect 6734 12671 6735 12697
rect 6761 12671 6762 12697
rect 6510 12474 6538 12479
rect 6398 12446 6510 12474
rect 2238 12166 2370 12171
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2238 12133 2370 12138
rect 4942 12025 4970 12031
rect 4942 11999 4943 12025
rect 4969 11999 4970 12025
rect 2142 11970 2170 11975
rect 2142 11923 2170 11942
rect 4942 11914 4970 11999
rect 6398 11969 6426 12446
rect 6510 12427 6538 12446
rect 6734 12418 6762 12671
rect 6790 12697 6818 13118
rect 6958 13145 6986 13151
rect 6958 13119 6959 13145
rect 6985 13119 6986 13145
rect 6958 13090 6986 13119
rect 7014 13090 7042 13510
rect 7070 13505 7098 13510
rect 7406 13481 7434 13487
rect 7406 13455 7407 13481
rect 7433 13455 7434 13481
rect 7406 13258 7434 13455
rect 7406 13225 7434 13230
rect 7462 13257 7490 13566
rect 8470 13594 8498 13599
rect 8526 13594 8554 18999
rect 9422 18746 9450 20600
rect 10094 19138 10122 20600
rect 10094 19105 10122 19110
rect 10878 19138 10906 19143
rect 10878 19091 10906 19110
rect 11438 19138 11466 20600
rect 12446 19306 12474 20600
rect 12782 19306 12810 20600
rect 12446 19278 12642 19306
rect 11438 19105 11466 19110
rect 10374 19025 10402 19031
rect 10374 18999 10375 19025
rect 10401 18999 10402 19025
rect 9918 18830 10050 18835
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 9918 18797 10050 18802
rect 9422 18713 9450 18718
rect 10038 18746 10066 18751
rect 10038 18699 10066 18718
rect 9534 18633 9562 18639
rect 9534 18607 9535 18633
rect 9561 18607 9562 18633
rect 9534 14377 9562 18607
rect 9918 18046 10050 18051
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 9918 18013 10050 18018
rect 9918 17262 10050 17267
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 9918 17229 10050 17234
rect 9918 16478 10050 16483
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 9918 16445 10050 16450
rect 10374 15974 10402 18999
rect 12278 19025 12306 19031
rect 12278 18999 12279 19025
rect 12305 18999 12306 19025
rect 12278 15974 12306 18999
rect 12614 18745 12642 19278
rect 12782 19273 12810 19278
rect 12782 19138 12810 19143
rect 12782 19091 12810 19110
rect 13118 19138 13146 20600
rect 13118 19105 13146 19110
rect 13398 19306 13426 19311
rect 12614 18719 12615 18745
rect 12641 18719 12642 18745
rect 12614 18713 12642 18719
rect 13398 18745 13426 19278
rect 17598 19222 17730 19227
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17598 19189 17730 19194
rect 14686 19138 14714 19143
rect 14686 19091 14714 19110
rect 13398 18719 13399 18745
rect 13425 18719 13426 18745
rect 13398 18713 13426 18719
rect 14294 19025 14322 19031
rect 14294 18999 14295 19025
rect 14321 18999 14322 19025
rect 12894 18633 12922 18639
rect 12894 18607 12895 18633
rect 12921 18607 12922 18633
rect 12894 15974 12922 18607
rect 10318 15946 10402 15974
rect 12110 15946 12306 15974
rect 12726 15946 12922 15974
rect 9918 15694 10050 15699
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 9918 15661 10050 15666
rect 9918 14910 10050 14915
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 9918 14877 10050 14882
rect 9534 14351 9535 14377
rect 9561 14351 9562 14377
rect 8918 14322 8946 14327
rect 8918 13930 8946 14294
rect 8974 14266 9002 14271
rect 9002 14238 9058 14266
rect 8974 14233 9002 14238
rect 8694 13929 8946 13930
rect 8694 13903 8919 13929
rect 8945 13903 8946 13929
rect 8694 13902 8946 13903
rect 8694 13594 8722 13902
rect 8918 13897 8946 13902
rect 8470 13593 8666 13594
rect 8470 13567 8471 13593
rect 8497 13567 8666 13593
rect 8470 13566 8666 13567
rect 8470 13561 8498 13566
rect 8638 13454 8666 13566
rect 8694 13593 8778 13594
rect 8694 13567 8695 13593
rect 8721 13567 8778 13593
rect 8694 13566 8778 13567
rect 8694 13561 8722 13566
rect 8638 13426 8722 13454
rect 7462 13231 7463 13257
rect 7489 13231 7490 13257
rect 7462 13225 7490 13231
rect 7910 13258 7938 13263
rect 7910 13211 7938 13230
rect 7182 13202 7210 13207
rect 7182 13201 7266 13202
rect 7182 13175 7183 13201
rect 7209 13175 7266 13201
rect 7182 13174 7266 13175
rect 7182 13169 7210 13174
rect 7126 13146 7154 13151
rect 6790 12671 6791 12697
rect 6817 12671 6818 12697
rect 6790 12665 6818 12671
rect 6846 13062 7042 13090
rect 7070 13145 7154 13146
rect 7070 13119 7127 13145
rect 7153 13119 7154 13145
rect 7070 13118 7154 13119
rect 6846 12474 6874 13062
rect 7070 12922 7098 13118
rect 7126 13113 7154 13118
rect 7182 13034 7210 13039
rect 7182 12987 7210 13006
rect 6902 12894 7098 12922
rect 6902 12753 6930 12894
rect 7238 12754 7266 13174
rect 8694 13201 8722 13426
rect 8694 13175 8695 13201
rect 8721 13175 8722 13201
rect 8694 13169 8722 13175
rect 7966 13090 7994 13095
rect 7966 13043 7994 13062
rect 7294 12754 7322 12759
rect 6902 12727 6903 12753
rect 6929 12727 6930 12753
rect 6902 12721 6930 12727
rect 7182 12726 7294 12754
rect 6846 12441 6874 12446
rect 7126 12641 7154 12647
rect 7126 12615 7127 12641
rect 7153 12615 7154 12641
rect 7126 12418 7154 12615
rect 6734 12385 6762 12390
rect 7070 12390 7126 12418
rect 7070 12026 7098 12390
rect 7126 12385 7154 12390
rect 6398 11943 6399 11969
rect 6425 11943 6426 11969
rect 6398 11937 6426 11943
rect 6846 12025 7098 12026
rect 6846 11999 7071 12025
rect 7097 11999 7098 12025
rect 6846 11998 7098 11999
rect 6846 11969 6874 11998
rect 7070 11993 7098 11998
rect 6846 11943 6847 11969
rect 6873 11943 6874 11969
rect 4942 11881 4970 11886
rect 6006 11914 6034 11919
rect 6790 11914 6818 11919
rect 6006 11913 6202 11914
rect 6006 11887 6007 11913
rect 6033 11887 6202 11913
rect 6006 11886 6202 11887
rect 6006 11881 6034 11886
rect 6006 11802 6034 11807
rect 2238 11382 2370 11387
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2238 11349 2370 11354
rect 2142 11186 2170 11191
rect 2142 11139 2170 11158
rect 5670 11186 5698 11191
rect 5670 10850 5698 11158
rect 2086 10761 2114 10766
rect 2142 10793 2170 10799
rect 2142 10767 2143 10793
rect 2169 10767 2170 10793
rect 966 10681 994 10687
rect 966 10655 967 10681
rect 993 10655 994 10681
rect 966 10458 994 10655
rect 966 10425 994 10430
rect 2142 10346 2170 10767
rect 5670 10737 5698 10822
rect 5670 10711 5671 10737
rect 5697 10711 5698 10737
rect 5670 10705 5698 10711
rect 2238 10598 2370 10603
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2238 10565 2370 10570
rect 6006 10402 6034 11774
rect 6174 11689 6202 11886
rect 6790 11867 6818 11886
rect 6678 11858 6706 11863
rect 6174 11663 6175 11689
rect 6201 11663 6202 11689
rect 6174 11657 6202 11663
rect 6342 11857 6706 11858
rect 6342 11831 6679 11857
rect 6705 11831 6706 11857
rect 6342 11830 6706 11831
rect 6286 11634 6314 11639
rect 6286 11587 6314 11606
rect 6342 11633 6370 11830
rect 6678 11825 6706 11830
rect 6846 11802 6874 11943
rect 6846 11769 6874 11774
rect 6342 11607 6343 11633
rect 6369 11607 6370 11633
rect 6342 11601 6370 11607
rect 7014 11634 7042 11639
rect 7014 11186 7042 11606
rect 7014 11139 7042 11158
rect 7126 11186 7154 11191
rect 7182 11186 7210 12726
rect 7294 12721 7322 12726
rect 7238 12474 7266 12479
rect 7238 11969 7266 12446
rect 7238 11943 7239 11969
rect 7265 11943 7266 11969
rect 7238 11937 7266 11943
rect 8078 12250 8106 12255
rect 7630 11914 7658 11919
rect 7630 11913 7714 11914
rect 7630 11887 7631 11913
rect 7657 11887 7714 11913
rect 7630 11886 7714 11887
rect 7630 11881 7658 11886
rect 7686 11521 7714 11886
rect 7686 11495 7687 11521
rect 7713 11495 7714 11521
rect 7686 11489 7714 11495
rect 7742 11634 7770 11639
rect 8022 11634 8050 11639
rect 7742 11633 8050 11634
rect 7742 11607 7743 11633
rect 7769 11607 8023 11633
rect 8049 11607 8050 11633
rect 7742 11606 8050 11607
rect 7742 11410 7770 11606
rect 8022 11601 8050 11606
rect 7854 11522 7882 11527
rect 8078 11522 8106 12222
rect 8750 12082 8778 13566
rect 9030 13537 9058 14238
rect 9254 13874 9282 13879
rect 9254 13827 9282 13846
rect 9534 13650 9562 14351
rect 9758 14322 9786 14327
rect 9758 14275 9786 14294
rect 9918 14126 10050 14131
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 9918 14093 10050 14098
rect 9590 13874 9618 13879
rect 9618 13846 9674 13874
rect 9590 13841 9618 13846
rect 9422 13622 9562 13650
rect 9646 13649 9674 13846
rect 9646 13623 9647 13649
rect 9673 13623 9674 13649
rect 9030 13511 9031 13537
rect 9057 13511 9058 13537
rect 9030 13505 9058 13511
rect 9142 13566 9282 13594
rect 9142 13481 9170 13566
rect 9254 13538 9282 13566
rect 9310 13538 9338 13543
rect 9254 13537 9338 13538
rect 9254 13511 9311 13537
rect 9337 13511 9338 13537
rect 9254 13510 9338 13511
rect 9310 13505 9338 13510
rect 9142 13455 9143 13481
rect 9169 13455 9170 13481
rect 9142 13449 9170 13455
rect 9198 13481 9226 13487
rect 9198 13455 9199 13481
rect 9225 13455 9226 13481
rect 8806 13258 8834 13263
rect 8806 13211 8834 13230
rect 8918 13145 8946 13151
rect 8918 13119 8919 13145
rect 8945 13119 8946 13145
rect 8862 13090 8890 13095
rect 8862 13043 8890 13062
rect 8918 12250 8946 13119
rect 9030 13146 9058 13151
rect 9030 13099 9058 13118
rect 9198 12642 9226 13455
rect 9422 13481 9450 13622
rect 9646 13617 9674 13623
rect 10318 13873 10346 15946
rect 12110 14377 12138 15946
rect 12110 14351 12111 14377
rect 12137 14351 12138 14377
rect 10710 14322 10738 14327
rect 11046 14322 11074 14327
rect 10710 14275 10738 14294
rect 10878 14321 11074 14322
rect 10878 14295 11047 14321
rect 11073 14295 11074 14321
rect 10878 14294 11074 14295
rect 10878 14041 10906 14294
rect 11046 14289 11074 14294
rect 11830 14322 11858 14327
rect 10878 14015 10879 14041
rect 10905 14015 10906 14041
rect 10878 14009 10906 14015
rect 11270 14042 11298 14047
rect 11270 13995 11298 14014
rect 10766 13986 10794 13991
rect 10766 13939 10794 13958
rect 11158 13986 11186 13991
rect 11158 13939 11186 13958
rect 10318 13847 10319 13873
rect 10345 13847 10346 13873
rect 9422 13455 9423 13481
rect 9449 13455 9450 13481
rect 9422 13449 9450 13455
rect 9478 13538 9506 13543
rect 9366 13258 9394 13263
rect 9478 13258 9506 13510
rect 9702 13482 9730 13487
rect 9702 13481 9842 13482
rect 9702 13455 9703 13481
rect 9729 13455 9842 13481
rect 9702 13454 9842 13455
rect 9702 13449 9730 13454
rect 9394 13230 9506 13258
rect 9814 13258 9842 13454
rect 9918 13342 10050 13347
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 9918 13309 10050 13314
rect 9926 13258 9954 13263
rect 9814 13257 9954 13258
rect 9814 13231 9927 13257
rect 9953 13231 9954 13257
rect 9814 13230 9954 13231
rect 9366 13211 9394 13230
rect 9926 13225 9954 13230
rect 9982 13258 10010 13263
rect 9982 13211 10010 13230
rect 10318 13258 10346 13847
rect 10710 13929 10738 13935
rect 10710 13903 10711 13929
rect 10737 13903 10738 13929
rect 10710 13454 10738 13903
rect 11326 13930 11354 13935
rect 11326 13538 11354 13902
rect 11326 13505 11354 13510
rect 11830 13537 11858 14294
rect 12110 14042 12138 14351
rect 12334 14322 12362 14327
rect 12334 14275 12362 14294
rect 12110 14009 12138 14014
rect 11830 13511 11831 13537
rect 11857 13511 11858 13537
rect 11830 13454 11858 13511
rect 10710 13426 10794 13454
rect 10318 13225 10346 13230
rect 9198 12609 9226 12614
rect 9422 13146 9450 13151
rect 9422 12474 9450 13118
rect 9534 13145 9562 13151
rect 9534 13119 9535 13145
rect 9561 13119 9562 13145
rect 9534 12754 9562 13119
rect 9758 13146 9786 13151
rect 9870 13146 9898 13151
rect 9758 13099 9786 13118
rect 9814 13145 9898 13146
rect 9814 13119 9871 13145
rect 9897 13119 9898 13145
rect 9814 13118 9898 13119
rect 9758 12754 9786 12759
rect 9534 12753 9786 12754
rect 9534 12727 9759 12753
rect 9785 12727 9786 12753
rect 9534 12726 9786 12727
rect 8918 12217 8946 12222
rect 9254 12446 9450 12474
rect 8750 12054 8946 12082
rect 8694 12026 8722 12031
rect 8694 11979 8722 11998
rect 8918 12025 8946 12054
rect 8918 11999 8919 12025
rect 8945 11999 8946 12025
rect 7854 11521 8106 11522
rect 7854 11495 7855 11521
rect 7881 11495 8106 11521
rect 7854 11494 8106 11495
rect 8134 11577 8162 11583
rect 8134 11551 8135 11577
rect 8161 11551 8162 11577
rect 7854 11489 7882 11494
rect 7126 11185 7210 11186
rect 7126 11159 7127 11185
rect 7153 11159 7210 11185
rect 7126 11158 7210 11159
rect 7630 11382 7770 11410
rect 7126 11153 7154 11158
rect 7350 11129 7378 11135
rect 7350 11103 7351 11129
rect 7377 11103 7378 11129
rect 6958 11074 6986 11079
rect 6734 11073 6986 11074
rect 6734 11047 6959 11073
rect 6985 11047 6986 11073
rect 6734 11046 6986 11047
rect 6734 10849 6762 11046
rect 6958 11041 6986 11046
rect 7238 11073 7266 11079
rect 7238 11047 7239 11073
rect 7265 11047 7266 11073
rect 7238 10962 7266 11047
rect 7238 10929 7266 10934
rect 7350 10906 7378 11103
rect 7350 10873 7378 10878
rect 6734 10823 6735 10849
rect 6761 10823 6762 10849
rect 6734 10817 6762 10823
rect 7126 10793 7154 10799
rect 7126 10767 7127 10793
rect 7153 10767 7154 10793
rect 7126 10738 7154 10767
rect 7518 10793 7546 10799
rect 7518 10767 7519 10793
rect 7545 10767 7546 10793
rect 7350 10738 7378 10743
rect 7126 10737 7378 10738
rect 7126 10711 7351 10737
rect 7377 10711 7378 10737
rect 7126 10710 7378 10711
rect 7126 10570 7154 10575
rect 6062 10514 6090 10519
rect 6062 10513 6482 10514
rect 6062 10487 6063 10513
rect 6089 10487 6482 10513
rect 6062 10486 6482 10487
rect 6062 10481 6090 10486
rect 6118 10402 6146 10407
rect 6342 10402 6370 10407
rect 6006 10401 6370 10402
rect 6006 10375 6119 10401
rect 6145 10375 6343 10401
rect 6369 10375 6370 10401
rect 6006 10374 6370 10375
rect 6118 10369 6146 10374
rect 6342 10369 6370 10374
rect 2142 10313 2170 10318
rect 4830 10290 4858 10295
rect 4830 9953 4858 10262
rect 6062 10290 6090 10295
rect 6062 10243 6090 10262
rect 6286 10066 6314 10071
rect 6286 10009 6314 10038
rect 6454 10065 6482 10486
rect 7126 10457 7154 10542
rect 7126 10431 7127 10457
rect 7153 10431 7154 10457
rect 7126 10425 7154 10431
rect 6790 10401 6818 10407
rect 6790 10375 6791 10401
rect 6817 10375 6818 10401
rect 6454 10039 6455 10065
rect 6481 10039 6482 10065
rect 6454 10033 6482 10039
rect 6510 10066 6538 10071
rect 6790 10066 6818 10375
rect 6510 10065 6594 10066
rect 6510 10039 6511 10065
rect 6537 10039 6594 10065
rect 6510 10038 6594 10039
rect 6510 10033 6538 10038
rect 6286 9983 6287 10009
rect 6313 9983 6314 10009
rect 6286 9977 6314 9983
rect 4830 9927 4831 9953
rect 4857 9927 4858 9953
rect 4830 9921 4858 9927
rect 5894 9953 5922 9959
rect 5894 9927 5895 9953
rect 5921 9927 5922 9953
rect 5894 9898 5922 9927
rect 6566 9954 6594 10038
rect 6790 10019 6818 10038
rect 7014 10066 7042 10071
rect 6566 9921 6594 9926
rect 6510 9898 6538 9903
rect 5894 9897 6538 9898
rect 5894 9871 6511 9897
rect 6537 9871 6538 9897
rect 5894 9870 6538 9871
rect 6510 9865 6538 9870
rect 2238 9814 2370 9819
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2238 9781 2370 9786
rect 7014 9506 7042 10038
rect 7350 10066 7378 10710
rect 7350 10033 7378 10038
rect 7462 10065 7490 10071
rect 7462 10039 7463 10065
rect 7489 10039 7490 10065
rect 6958 9505 7042 9506
rect 6958 9479 7015 9505
rect 7041 9479 7042 9505
rect 6958 9478 7042 9479
rect 2142 9226 2170 9231
rect 2142 9179 2170 9198
rect 5446 9226 5474 9231
rect 6510 9226 6538 9231
rect 5446 9169 5474 9198
rect 5446 9143 5447 9169
rect 5473 9143 5474 9169
rect 5446 9137 5474 9143
rect 6174 9225 6538 9226
rect 6174 9199 6511 9225
rect 6537 9199 6538 9225
rect 6174 9198 6538 9199
rect 966 9114 994 9119
rect 966 9067 994 9086
rect 2238 9030 2370 9035
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2238 8997 2370 9002
rect 966 8890 994 8895
rect 966 8843 994 8862
rect 2142 8834 2170 8839
rect 2142 8787 2170 8806
rect 6174 8777 6202 9198
rect 6510 9193 6538 9198
rect 6902 9226 6930 9231
rect 6958 9226 6986 9478
rect 7014 9473 7042 9478
rect 7182 9673 7210 9679
rect 7182 9647 7183 9673
rect 7209 9647 7210 9673
rect 6902 9225 6986 9226
rect 6902 9199 6903 9225
rect 6929 9199 6986 9225
rect 6902 9198 6986 9199
rect 6902 9193 6930 9198
rect 6342 9114 6370 9119
rect 6342 8833 6370 9086
rect 6342 8807 6343 8833
rect 6369 8807 6370 8833
rect 6342 8801 6370 8807
rect 6846 8834 6874 8839
rect 6174 8751 6175 8777
rect 6201 8751 6202 8777
rect 6174 8745 6202 8751
rect 6846 8777 6874 8806
rect 6846 8751 6847 8777
rect 6873 8751 6874 8777
rect 6846 8745 6874 8751
rect 6958 8441 6986 9198
rect 7014 9226 7042 9231
rect 7182 9226 7210 9647
rect 7350 9617 7378 9623
rect 7350 9591 7351 9617
rect 7377 9591 7378 9617
rect 7294 9562 7322 9567
rect 7294 9515 7322 9534
rect 7350 9282 7378 9591
rect 7462 9505 7490 10039
rect 7518 9562 7546 10767
rect 7518 9529 7546 9534
rect 7574 10626 7602 10631
rect 7630 10626 7658 11382
rect 7910 11186 7938 11191
rect 7742 10906 7770 10911
rect 7742 10859 7770 10878
rect 7686 10850 7714 10855
rect 7686 10803 7714 10822
rect 7602 10598 7658 10626
rect 7798 10793 7826 10799
rect 7798 10767 7799 10793
rect 7825 10767 7826 10793
rect 7462 9479 7463 9505
rect 7489 9479 7490 9505
rect 7294 9254 7378 9282
rect 7406 9282 7434 9287
rect 7462 9282 7490 9479
rect 7574 9505 7602 10598
rect 7742 10122 7770 10127
rect 7742 10065 7770 10094
rect 7742 10039 7743 10065
rect 7769 10039 7770 10065
rect 7742 10033 7770 10039
rect 7798 9618 7826 10767
rect 7910 10793 7938 11158
rect 8134 10906 8162 11551
rect 8918 11242 8946 11999
rect 9086 11970 9114 11975
rect 9086 11857 9114 11942
rect 9086 11831 9087 11857
rect 9113 11831 9114 11857
rect 9030 11578 9058 11583
rect 7910 10767 7911 10793
rect 7937 10767 7938 10793
rect 7854 10122 7882 10127
rect 7910 10122 7938 10767
rect 7854 10121 7938 10122
rect 7854 10095 7855 10121
rect 7881 10095 7938 10121
rect 7854 10094 7938 10095
rect 7966 10878 8162 10906
rect 8470 11241 8946 11242
rect 8470 11215 8919 11241
rect 8945 11215 8946 11241
rect 8470 11214 8946 11215
rect 7966 10234 7994 10878
rect 7854 10089 7882 10094
rect 7910 10010 7938 10015
rect 7966 10010 7994 10206
rect 8134 10793 8162 10799
rect 8134 10767 8135 10793
rect 8161 10767 8162 10793
rect 8134 10122 8162 10767
rect 8246 10793 8274 10799
rect 8246 10767 8247 10793
rect 8273 10767 8274 10793
rect 8190 10737 8218 10743
rect 8190 10711 8191 10737
rect 8217 10711 8218 10737
rect 8190 10570 8218 10711
rect 8246 10626 8274 10767
rect 8246 10593 8274 10598
rect 8190 10537 8218 10542
rect 8190 10458 8218 10463
rect 8190 10457 8386 10458
rect 8190 10431 8191 10457
rect 8217 10431 8386 10457
rect 8190 10430 8386 10431
rect 8190 10425 8218 10430
rect 8162 10094 8218 10122
rect 8134 10089 8162 10094
rect 7910 10009 7994 10010
rect 7910 9983 7911 10009
rect 7937 9983 7994 10009
rect 7910 9982 7994 9983
rect 7910 9977 7938 9982
rect 7798 9585 7826 9590
rect 7966 9506 7994 9511
rect 7574 9479 7575 9505
rect 7601 9479 7602 9505
rect 7574 9337 7602 9479
rect 7574 9311 7575 9337
rect 7601 9311 7602 9337
rect 7574 9305 7602 9311
rect 7686 9505 7994 9506
rect 7686 9479 7967 9505
rect 7993 9479 7994 9505
rect 7686 9478 7994 9479
rect 7686 9338 7714 9478
rect 7966 9473 7994 9478
rect 8134 9506 8162 9511
rect 8134 9459 8162 9478
rect 7686 9291 7714 9310
rect 7798 9338 7826 9343
rect 7798 9291 7826 9310
rect 7434 9254 7490 9282
rect 7238 9226 7266 9231
rect 7182 9225 7266 9226
rect 7182 9199 7239 9225
rect 7265 9199 7266 9225
rect 7182 9198 7266 9199
rect 7014 8834 7042 9198
rect 7238 9193 7266 9198
rect 7070 9114 7098 9119
rect 7070 9067 7098 9086
rect 7238 8946 7266 8951
rect 7294 8946 7322 9254
rect 7350 9170 7378 9175
rect 7350 9123 7378 9142
rect 7238 8945 7322 8946
rect 7238 8919 7239 8945
rect 7265 8919 7322 8945
rect 7238 8918 7322 8919
rect 7238 8913 7266 8918
rect 7294 8834 7322 8839
rect 7406 8834 7434 9254
rect 7630 9169 7658 9175
rect 7630 9143 7631 9169
rect 7657 9143 7658 9169
rect 7518 8890 7546 8895
rect 7630 8890 7658 9143
rect 7518 8889 7658 8890
rect 7518 8863 7519 8889
rect 7545 8863 7658 8889
rect 7518 8862 7658 8863
rect 7518 8857 7546 8862
rect 7014 8833 7266 8834
rect 7014 8807 7015 8833
rect 7041 8807 7266 8833
rect 7014 8806 7266 8807
rect 7014 8801 7042 8806
rect 7238 8777 7266 8806
rect 7294 8833 7434 8834
rect 7294 8807 7295 8833
rect 7321 8807 7434 8833
rect 7294 8806 7434 8807
rect 7294 8801 7322 8806
rect 7238 8751 7239 8777
rect 7265 8751 7266 8777
rect 7238 8745 7266 8751
rect 7462 8722 7490 8727
rect 7350 8721 7490 8722
rect 7350 8695 7463 8721
rect 7489 8695 7490 8721
rect 7350 8694 7490 8695
rect 7350 8497 7378 8694
rect 7462 8689 7490 8694
rect 7350 8471 7351 8497
rect 7377 8471 7378 8497
rect 7350 8465 7378 8471
rect 6958 8415 6959 8441
rect 6985 8415 6986 8441
rect 6958 8409 6986 8415
rect 8190 8442 8218 10094
rect 8246 10065 8274 10430
rect 8358 10401 8386 10430
rect 8358 10375 8359 10401
rect 8385 10375 8386 10401
rect 8358 10369 8386 10375
rect 8302 10290 8330 10295
rect 8302 10121 8330 10262
rect 8302 10095 8303 10121
rect 8329 10095 8330 10121
rect 8302 10089 8330 10095
rect 8246 10039 8247 10065
rect 8273 10039 8274 10065
rect 8246 10033 8274 10039
rect 8470 10066 8498 11214
rect 8918 11209 8946 11214
rect 8974 11465 9002 11471
rect 8974 11439 8975 11465
rect 9001 11439 9002 11465
rect 8750 10962 8778 10967
rect 8974 10962 9002 11439
rect 9030 11018 9058 11550
rect 9030 10985 9058 10990
rect 8694 10934 8750 10962
rect 8526 10289 8554 10295
rect 8526 10263 8527 10289
rect 8553 10263 8554 10289
rect 8526 10066 8554 10263
rect 8638 10066 8666 10071
rect 8526 10038 8638 10066
rect 8358 9674 8386 9679
rect 8470 9674 8498 10038
rect 8638 9730 8666 10038
rect 8694 9954 8722 10934
rect 8750 10929 8778 10934
rect 8918 10934 9002 10962
rect 8862 10794 8890 10799
rect 8918 10794 8946 10934
rect 9086 10906 9114 11831
rect 9254 11913 9282 12446
rect 9254 11887 9255 11913
rect 9281 11887 9282 11913
rect 9254 11802 9282 11887
rect 9310 12361 9338 12367
rect 9310 12335 9311 12361
rect 9337 12335 9338 12361
rect 9310 12026 9338 12335
rect 9310 11858 9338 11998
rect 9422 11969 9450 12446
rect 9590 12642 9618 12647
rect 9422 11943 9423 11969
rect 9449 11943 9450 11969
rect 9422 11937 9450 11943
rect 9478 12417 9506 12423
rect 9478 12391 9479 12417
rect 9505 12391 9506 12417
rect 9478 11914 9506 12391
rect 9310 11830 9394 11858
rect 9254 11774 9338 11802
rect 9198 11746 9226 11751
rect 9142 11577 9170 11583
rect 9142 11551 9143 11577
rect 9169 11551 9170 11577
rect 9142 10962 9170 11551
rect 9142 10929 9170 10934
rect 9030 10878 9114 10906
rect 8974 10850 9002 10855
rect 8974 10803 9002 10822
rect 8862 10793 8946 10794
rect 8862 10767 8863 10793
rect 8889 10767 8946 10793
rect 8862 10766 8946 10767
rect 8862 10761 8890 10766
rect 8750 10401 8778 10407
rect 8750 10375 8751 10401
rect 8777 10375 8778 10401
rect 8750 10066 8778 10375
rect 8862 10346 8890 10351
rect 8862 10299 8890 10318
rect 8750 10033 8778 10038
rect 8918 10010 8946 10766
rect 9030 10738 9058 10878
rect 9142 10738 9170 10757
rect 9030 10710 9114 10738
rect 9030 10345 9058 10351
rect 9030 10319 9031 10345
rect 9057 10319 9058 10345
rect 8974 10010 9002 10015
rect 8918 9982 8974 10010
rect 8974 9977 9002 9982
rect 8750 9954 8778 9959
rect 8694 9953 8778 9954
rect 8694 9927 8751 9953
rect 8777 9927 8778 9953
rect 8694 9926 8778 9927
rect 8750 9921 8778 9926
rect 8806 9898 8834 9903
rect 8806 9851 8834 9870
rect 8974 9897 9002 9903
rect 8974 9871 8975 9897
rect 9001 9871 9002 9897
rect 8918 9842 8946 9847
rect 8638 9702 8834 9730
rect 8358 9673 8778 9674
rect 8358 9647 8359 9673
rect 8385 9647 8778 9673
rect 8358 9646 8778 9647
rect 8358 9641 8386 9646
rect 8638 9562 8666 9567
rect 8638 9515 8666 9534
rect 8694 9225 8722 9231
rect 8694 9199 8695 9225
rect 8721 9199 8722 9225
rect 8358 9170 8386 9175
rect 8358 8946 8386 9142
rect 8694 9170 8722 9199
rect 8694 9137 8722 9142
rect 8414 9114 8442 9119
rect 8414 9067 8442 9086
rect 8358 8918 8442 8946
rect 8190 8409 8218 8414
rect 8414 8385 8442 8918
rect 8750 8553 8778 9646
rect 8806 9617 8834 9702
rect 8806 9591 8807 9617
rect 8833 9591 8834 9617
rect 8806 9585 8834 9591
rect 8918 9562 8946 9814
rect 8918 9529 8946 9534
rect 8974 9506 9002 9871
rect 8862 9281 8890 9287
rect 8862 9255 8863 9281
rect 8889 9255 8890 9281
rect 8862 9226 8890 9255
rect 8974 9226 9002 9478
rect 8862 9198 8974 9226
rect 8974 9193 9002 9198
rect 9030 9226 9058 10319
rect 9086 9953 9114 10710
rect 9142 10705 9170 10710
rect 9142 10626 9170 10631
rect 9142 10290 9170 10598
rect 9198 10513 9226 11718
rect 9254 11633 9282 11639
rect 9254 11607 9255 11633
rect 9281 11607 9282 11633
rect 9254 10906 9282 11607
rect 9310 11633 9338 11774
rect 9310 11607 9311 11633
rect 9337 11607 9338 11633
rect 9310 11601 9338 11607
rect 9254 10873 9282 10878
rect 9254 10794 9282 10799
rect 9366 10794 9394 11830
rect 9478 11689 9506 11886
rect 9478 11663 9479 11689
rect 9505 11663 9506 11689
rect 9478 11657 9506 11663
rect 9534 12026 9562 12031
rect 9534 11913 9562 11998
rect 9534 11887 9535 11913
rect 9561 11887 9562 11913
rect 9534 10850 9562 11887
rect 9590 11858 9618 12614
rect 9702 12417 9730 12423
rect 9702 12391 9703 12417
rect 9729 12391 9730 12417
rect 9646 12250 9674 12255
rect 9646 12203 9674 12222
rect 9646 11858 9674 11863
rect 9590 11857 9674 11858
rect 9590 11831 9647 11857
rect 9673 11831 9674 11857
rect 9590 11830 9674 11831
rect 9534 10817 9562 10822
rect 9254 10793 9394 10794
rect 9254 10767 9255 10793
rect 9281 10767 9394 10793
rect 9254 10766 9394 10767
rect 9590 10794 9618 10799
rect 9254 10761 9282 10766
rect 9590 10747 9618 10766
rect 9422 10682 9450 10687
rect 9422 10681 9506 10682
rect 9422 10655 9423 10681
rect 9449 10655 9506 10681
rect 9422 10654 9506 10655
rect 9422 10649 9450 10654
rect 9198 10487 9199 10513
rect 9225 10487 9226 10513
rect 9198 10481 9226 10487
rect 9142 10243 9170 10262
rect 9198 10402 9226 10407
rect 9142 10066 9170 10071
rect 9142 10009 9170 10038
rect 9142 9983 9143 10009
rect 9169 9983 9170 10009
rect 9142 9977 9170 9983
rect 9086 9927 9087 9953
rect 9113 9927 9114 9953
rect 9086 9921 9114 9927
rect 9142 9562 9170 9567
rect 9198 9562 9226 10374
rect 9478 10402 9506 10654
rect 9646 10626 9674 11830
rect 9702 11522 9730 12391
rect 9758 11746 9786 12726
rect 9814 12474 9842 13118
rect 9870 13113 9898 13118
rect 10094 13145 10122 13151
rect 10094 13119 10095 13145
rect 10121 13119 10122 13145
rect 9870 12698 9898 12703
rect 9870 12651 9898 12670
rect 10094 12698 10122 13119
rect 10654 12754 10682 12759
rect 10654 12707 10682 12726
rect 10766 12753 10794 13426
rect 11494 13426 11858 13454
rect 12110 13930 12138 13935
rect 11438 13258 11466 13263
rect 11382 13145 11410 13151
rect 11382 13119 11383 13145
rect 11409 13119 11410 13145
rect 11382 13090 11410 13119
rect 11382 13057 11410 13062
rect 11438 13145 11466 13230
rect 11438 13119 11439 13145
rect 11465 13119 11466 13145
rect 10934 12866 10962 12871
rect 10934 12819 10962 12838
rect 11438 12866 11466 13119
rect 11438 12833 11466 12838
rect 10766 12727 10767 12753
rect 10793 12727 10794 12753
rect 10094 12665 10122 12670
rect 9918 12558 10050 12563
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 9918 12525 10050 12530
rect 9814 12446 10010 12474
rect 9982 12305 10010 12446
rect 9982 12279 9983 12305
rect 10009 12279 10010 12305
rect 9982 12273 10010 12279
rect 10038 12417 10066 12423
rect 10038 12391 10039 12417
rect 10065 12391 10066 12417
rect 9814 12250 9842 12255
rect 9814 12203 9842 12222
rect 10038 12082 10066 12391
rect 10150 12250 10178 12255
rect 10178 12222 10234 12250
rect 10150 12203 10178 12222
rect 9982 12054 10066 12082
rect 9982 12026 10010 12054
rect 9982 11993 10010 11998
rect 10094 11970 10122 11975
rect 10094 11923 10122 11942
rect 9758 11713 9786 11718
rect 9814 11913 9842 11919
rect 9814 11887 9815 11913
rect 9841 11887 9842 11913
rect 9814 11858 9842 11887
rect 10038 11914 10066 11919
rect 10038 11858 10066 11886
rect 10206 11914 10234 12222
rect 10430 12082 10458 12087
rect 10766 12082 10794 12727
rect 10430 12081 10794 12082
rect 10430 12055 10431 12081
rect 10457 12055 10794 12081
rect 10430 12054 10794 12055
rect 11158 12754 11186 12759
rect 10430 12049 10458 12054
rect 10206 11881 10234 11886
rect 10710 11969 10738 11975
rect 10710 11943 10711 11969
rect 10737 11943 10738 11969
rect 10262 11858 10290 11863
rect 10038 11830 10122 11858
rect 9702 11489 9730 11494
rect 9758 11522 9786 11527
rect 9814 11522 9842 11830
rect 10094 11802 10122 11830
rect 10262 11811 10290 11830
rect 10374 11857 10402 11863
rect 10374 11831 10375 11857
rect 10401 11831 10402 11857
rect 9918 11774 10050 11779
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 9918 11741 10050 11746
rect 10094 11690 10122 11774
rect 10038 11662 10122 11690
rect 10038 11577 10066 11662
rect 10038 11551 10039 11577
rect 10065 11551 10066 11577
rect 10038 11545 10066 11551
rect 9758 11521 9842 11522
rect 9758 11495 9759 11521
rect 9785 11495 9842 11521
rect 9758 11494 9842 11495
rect 9926 11522 9954 11527
rect 9702 11185 9730 11191
rect 9702 11159 9703 11185
rect 9729 11159 9730 11185
rect 9702 10738 9730 11159
rect 9758 10906 9786 11494
rect 9926 11475 9954 11494
rect 10374 11522 10402 11831
rect 10710 11802 10738 11943
rect 11102 11914 11130 11919
rect 10822 11858 10850 11863
rect 10822 11811 10850 11830
rect 10710 11769 10738 11774
rect 10654 11578 10682 11583
rect 11046 11578 11074 11583
rect 10654 11531 10682 11550
rect 10934 11577 11074 11578
rect 10934 11551 11047 11577
rect 11073 11551 11074 11577
rect 10934 11550 11074 11551
rect 10374 11489 10402 11494
rect 10878 11522 10906 11527
rect 10206 11466 10234 11471
rect 10206 11419 10234 11438
rect 10878 11130 10906 11494
rect 10878 11097 10906 11102
rect 10934 11185 10962 11550
rect 11046 11545 11074 11550
rect 10934 11159 10935 11185
rect 10961 11159 10962 11185
rect 9918 10990 10050 10995
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 9918 10957 10050 10962
rect 9758 10873 9786 10878
rect 10150 10906 10178 10911
rect 9702 10705 9730 10710
rect 9646 10598 9730 10626
rect 9646 10402 9674 10407
rect 9478 10401 9674 10402
rect 9478 10375 9479 10401
rect 9505 10375 9647 10401
rect 9673 10375 9674 10401
rect 9478 10374 9674 10375
rect 9478 10369 9506 10374
rect 9646 10369 9674 10374
rect 9366 10289 9394 10295
rect 9366 10263 9367 10289
rect 9393 10263 9394 10289
rect 9366 10234 9394 10263
rect 9366 10201 9394 10206
rect 9310 10066 9338 10071
rect 9590 10066 9618 10071
rect 9310 10009 9338 10038
rect 9310 9983 9311 10009
rect 9337 9983 9338 10009
rect 9310 9977 9338 9983
rect 9422 10065 9618 10066
rect 9422 10039 9591 10065
rect 9617 10039 9618 10065
rect 9422 10038 9618 10039
rect 9366 9954 9394 9959
rect 9366 9907 9394 9926
rect 9142 9561 9226 9562
rect 9142 9535 9143 9561
rect 9169 9535 9226 9561
rect 9142 9534 9226 9535
rect 9310 9730 9338 9735
rect 9310 9618 9338 9702
rect 9142 9529 9170 9534
rect 9142 9226 9170 9231
rect 9030 9225 9170 9226
rect 9030 9199 9143 9225
rect 9169 9199 9170 9225
rect 9030 9198 9170 9199
rect 9030 9114 9058 9198
rect 9142 9193 9170 9198
rect 9030 9081 9058 9086
rect 9310 9058 9338 9590
rect 9366 9674 9394 9679
rect 9366 9617 9394 9646
rect 9366 9591 9367 9617
rect 9393 9591 9394 9617
rect 9366 9338 9394 9591
rect 9366 9305 9394 9310
rect 9422 9450 9450 10038
rect 9590 10033 9618 10038
rect 9478 9562 9506 9567
rect 9702 9562 9730 10598
rect 10094 10401 10122 10407
rect 10094 10375 10095 10401
rect 10121 10375 10122 10401
rect 10094 10346 10122 10375
rect 10094 10313 10122 10318
rect 9918 10206 10050 10211
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 9918 10173 10050 10178
rect 10094 10065 10122 10071
rect 10094 10039 10095 10065
rect 10121 10039 10122 10065
rect 10094 10010 10122 10039
rect 10094 9977 10122 9982
rect 10150 10009 10178 10878
rect 10710 10794 10738 10799
rect 10318 10570 10346 10575
rect 10318 10402 10346 10542
rect 10710 10457 10738 10766
rect 10934 10626 10962 11159
rect 10934 10593 10962 10598
rect 10990 11129 11018 11135
rect 10990 11103 10991 11129
rect 11017 11103 11018 11129
rect 10878 10570 10906 10575
rect 10710 10431 10711 10457
rect 10737 10431 10738 10457
rect 10710 10425 10738 10431
rect 10822 10542 10878 10570
rect 10318 10355 10346 10374
rect 10822 10401 10850 10542
rect 10878 10537 10906 10542
rect 10822 10375 10823 10401
rect 10849 10375 10850 10401
rect 10822 10369 10850 10375
rect 10150 9983 10151 10009
rect 10177 9983 10178 10009
rect 10150 9977 10178 9983
rect 10262 10345 10290 10351
rect 10262 10319 10263 10345
rect 10289 10319 10290 10345
rect 9982 9954 10010 9959
rect 9478 9561 9730 9562
rect 9478 9535 9479 9561
rect 9505 9535 9730 9561
rect 9478 9534 9730 9535
rect 9758 9617 9786 9623
rect 9758 9591 9759 9617
rect 9785 9591 9786 9617
rect 9758 9562 9786 9591
rect 9982 9618 10010 9926
rect 10262 9674 10290 10319
rect 10934 9898 10962 9903
rect 10262 9641 10290 9646
rect 10822 9673 10850 9679
rect 10822 9647 10823 9673
rect 10849 9647 10850 9673
rect 9982 9571 10010 9590
rect 10598 9618 10626 9623
rect 10598 9571 10626 9590
rect 9478 9529 9506 9534
rect 9758 9529 9786 9534
rect 10766 9562 10794 9567
rect 10038 9506 10066 9511
rect 10206 9506 10234 9511
rect 10038 9505 10122 9506
rect 10038 9479 10039 9505
rect 10065 9479 10122 9505
rect 10038 9478 10122 9479
rect 10038 9473 10066 9478
rect 9422 9422 9842 9450
rect 9422 9225 9450 9422
rect 9422 9199 9423 9225
rect 9449 9199 9450 9225
rect 9422 9193 9450 9199
rect 9646 9338 9674 9343
rect 9310 9030 9506 9058
rect 8750 8527 8751 8553
rect 8777 8527 8778 8553
rect 8414 8359 8415 8385
rect 8441 8359 8442 8385
rect 8414 8353 8442 8359
rect 8694 8386 8722 8391
rect 2238 8246 2370 8251
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2238 8213 2370 8218
rect 2238 7462 2370 7467
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2238 7429 2370 7434
rect 8694 7321 8722 8358
rect 8694 7295 8695 7321
rect 8721 7295 8722 7321
rect 8694 7289 8722 7295
rect 8358 7266 8386 7271
rect 8358 7219 8386 7238
rect 8750 7266 8778 8527
rect 9478 8498 9506 9030
rect 9254 8442 9282 8447
rect 9254 8395 9282 8414
rect 9478 8441 9506 8470
rect 9646 8497 9674 9310
rect 9814 8554 9842 9422
rect 9918 9422 10050 9427
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 9918 9389 10050 9394
rect 10094 9338 10122 9478
rect 10038 9310 10122 9338
rect 9926 9226 9954 9231
rect 9926 9179 9954 9198
rect 10038 9170 10066 9310
rect 10206 9281 10234 9478
rect 10206 9255 10207 9281
rect 10233 9255 10234 9281
rect 10206 9249 10234 9255
rect 10766 9505 10794 9534
rect 10766 9479 10767 9505
rect 10793 9479 10794 9505
rect 10766 9282 10794 9479
rect 10766 9249 10794 9254
rect 10038 9137 10066 9142
rect 10822 8946 10850 9647
rect 10878 9674 10906 9679
rect 10878 9561 10906 9646
rect 10878 9535 10879 9561
rect 10905 9535 10906 9561
rect 10878 9529 10906 9535
rect 10934 9226 10962 9870
rect 10990 9506 11018 11103
rect 11102 10570 11130 11886
rect 11158 11241 11186 12726
rect 11382 12754 11410 12759
rect 11494 12754 11522 13426
rect 11886 13258 11914 13263
rect 11662 13145 11690 13151
rect 11662 13119 11663 13145
rect 11689 13119 11690 13145
rect 11550 13089 11578 13095
rect 11550 13063 11551 13089
rect 11577 13063 11578 13089
rect 11550 12922 11578 13063
rect 11662 12978 11690 13119
rect 11774 13145 11802 13151
rect 11774 13119 11775 13145
rect 11801 13119 11802 13145
rect 11774 13034 11802 13119
rect 11886 13145 11914 13230
rect 11886 13119 11887 13145
rect 11913 13119 11914 13145
rect 11886 13113 11914 13119
rect 12110 13145 12138 13902
rect 12166 13481 12194 13487
rect 12166 13455 12167 13481
rect 12193 13455 12194 13481
rect 12166 13257 12194 13455
rect 12166 13231 12167 13257
rect 12193 13231 12194 13257
rect 12166 13225 12194 13231
rect 12110 13119 12111 13145
rect 12137 13119 12138 13145
rect 12110 13113 12138 13119
rect 12222 13146 12250 13151
rect 12222 13099 12250 13118
rect 11998 13090 12026 13095
rect 11998 13043 12026 13062
rect 12390 13090 12418 13095
rect 11774 13006 11858 13034
rect 11662 12950 11802 12978
rect 11550 12894 11746 12922
rect 11718 12809 11746 12894
rect 11718 12783 11719 12809
rect 11745 12783 11746 12809
rect 11718 12777 11746 12783
rect 11382 12753 11522 12754
rect 11382 12727 11383 12753
rect 11409 12727 11522 12753
rect 11382 12726 11522 12727
rect 11382 12642 11410 12726
rect 11382 12609 11410 12614
rect 11550 12698 11578 12703
rect 11550 12361 11578 12670
rect 11774 12530 11802 12950
rect 11830 12698 11858 13006
rect 11830 12665 11858 12670
rect 11774 12502 12026 12530
rect 11998 12473 12026 12502
rect 11998 12447 11999 12473
rect 12025 12447 12026 12473
rect 11998 12441 12026 12447
rect 11550 12335 11551 12361
rect 11577 12335 11578 12361
rect 11550 12306 11578 12335
rect 11550 12273 11578 12278
rect 11662 12418 11690 12423
rect 11606 12025 11634 12031
rect 11606 11999 11607 12025
rect 11633 11999 11634 12025
rect 11270 11858 11298 11863
rect 11158 11215 11159 11241
rect 11185 11215 11186 11241
rect 11158 11209 11186 11215
rect 11214 11634 11242 11639
rect 11046 10542 11130 10570
rect 11214 10570 11242 11606
rect 11270 11298 11298 11830
rect 11438 11802 11466 11807
rect 11326 11522 11354 11527
rect 11326 11475 11354 11494
rect 11382 11298 11410 11303
rect 11270 11270 11382 11298
rect 11046 10401 11074 10542
rect 11214 10537 11242 10542
rect 11326 10738 11354 10743
rect 11102 10458 11130 10463
rect 11102 10411 11130 10430
rect 11046 10375 11047 10401
rect 11073 10375 11074 10401
rect 11046 9842 11074 10375
rect 11326 10401 11354 10710
rect 11326 10375 11327 10401
rect 11353 10375 11354 10401
rect 11326 10369 11354 10375
rect 11046 9809 11074 9814
rect 11102 10346 11130 10351
rect 10990 9473 11018 9478
rect 11046 9618 11074 9623
rect 11046 9338 11074 9590
rect 11046 9281 11074 9310
rect 11102 9338 11130 10318
rect 11158 10290 11186 10295
rect 11158 9618 11186 10262
rect 11382 10121 11410 11270
rect 11438 11242 11466 11774
rect 11606 11578 11634 11999
rect 11662 11858 11690 12390
rect 12110 12418 12138 12423
rect 12110 12371 12138 12390
rect 11662 11825 11690 11830
rect 11886 12362 11914 12367
rect 11606 11545 11634 11550
rect 11662 11634 11690 11639
rect 11662 11577 11690 11606
rect 11886 11633 11914 12334
rect 11942 12361 11970 12367
rect 11942 12335 11943 12361
rect 11969 12335 11970 12361
rect 11942 11914 11970 12335
rect 12222 12362 12250 12367
rect 12222 12315 12250 12334
rect 11942 11881 11970 11886
rect 11886 11607 11887 11633
rect 11913 11607 11914 11633
rect 11886 11601 11914 11607
rect 11662 11551 11663 11577
rect 11689 11551 11690 11577
rect 11662 11545 11690 11551
rect 11718 11522 11746 11527
rect 11438 11214 11690 11242
rect 11438 11130 11466 11135
rect 11438 11083 11466 11102
rect 11382 10095 11383 10121
rect 11409 10095 11410 10121
rect 11382 10089 11410 10095
rect 11438 10570 11466 10575
rect 11270 10009 11298 10015
rect 11270 9983 11271 10009
rect 11297 9983 11298 10009
rect 11270 9730 11298 9983
rect 11326 9954 11354 9959
rect 11326 9907 11354 9926
rect 11270 9697 11298 9702
rect 11270 9618 11298 9623
rect 11158 9617 11298 9618
rect 11158 9591 11271 9617
rect 11297 9591 11298 9617
rect 11158 9590 11298 9591
rect 11270 9585 11298 9590
rect 11326 9562 11354 9567
rect 11326 9515 11354 9534
rect 11382 9506 11410 9511
rect 11382 9459 11410 9478
rect 11158 9338 11186 9343
rect 11102 9337 11158 9338
rect 11102 9311 11103 9337
rect 11129 9311 11158 9337
rect 11102 9310 11158 9311
rect 11102 9305 11130 9310
rect 11158 9305 11186 9310
rect 11382 9338 11410 9343
rect 11382 9291 11410 9310
rect 11046 9255 11047 9281
rect 11073 9255 11074 9281
rect 11046 9249 11074 9255
rect 11438 9281 11466 10542
rect 11606 10178 11634 10183
rect 11606 10009 11634 10150
rect 11662 10066 11690 11214
rect 11718 10402 11746 11494
rect 11830 11465 11858 11471
rect 11830 11439 11831 11465
rect 11857 11439 11858 11465
rect 11774 11298 11802 11303
rect 11830 11298 11858 11439
rect 11802 11270 11858 11298
rect 11774 11265 11802 11270
rect 12222 11186 12250 11191
rect 11886 11185 12250 11186
rect 11886 11159 12223 11185
rect 12249 11159 12250 11185
rect 11886 11158 12250 11159
rect 11718 10374 11802 10402
rect 11774 10122 11802 10374
rect 11718 10066 11746 10071
rect 11662 10065 11746 10066
rect 11662 10039 11719 10065
rect 11745 10039 11746 10065
rect 11662 10038 11746 10039
rect 11718 10033 11746 10038
rect 11606 9983 11607 10009
rect 11633 9983 11634 10009
rect 11550 9617 11578 9623
rect 11550 9591 11551 9617
rect 11577 9591 11578 9617
rect 11494 9338 11522 9343
rect 11550 9338 11578 9591
rect 11522 9310 11578 9338
rect 11494 9305 11522 9310
rect 11438 9255 11439 9281
rect 11465 9255 11466 9281
rect 11438 9249 11466 9255
rect 11102 9226 11130 9231
rect 11214 9226 11242 9231
rect 10934 9198 11018 9226
rect 10822 8913 10850 8918
rect 10934 9114 10962 9119
rect 10934 8889 10962 9086
rect 10990 8946 11018 9198
rect 11130 9198 11186 9226
rect 11102 9193 11130 9198
rect 11158 9114 11186 9198
rect 11214 9179 11242 9198
rect 11270 9225 11298 9231
rect 11270 9199 11271 9225
rect 11297 9199 11298 9225
rect 11270 9114 11298 9199
rect 11606 9226 11634 9983
rect 11606 9193 11634 9198
rect 11662 9954 11690 9959
rect 11158 9086 11298 9114
rect 11046 8946 11074 8951
rect 10990 8945 11074 8946
rect 10990 8919 11047 8945
rect 11073 8919 11074 8945
rect 10990 8918 11074 8919
rect 11046 8913 11074 8918
rect 11158 8946 11186 8951
rect 11158 8899 11186 8918
rect 10934 8863 10935 8889
rect 10961 8863 10962 8889
rect 10934 8857 10962 8863
rect 10822 8834 10850 8839
rect 10654 8833 10850 8834
rect 10654 8807 10823 8833
rect 10849 8807 10850 8833
rect 10654 8806 10850 8807
rect 9918 8638 10050 8643
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 9918 8605 10050 8610
rect 9646 8471 9647 8497
rect 9673 8471 9674 8497
rect 9646 8465 9674 8471
rect 9702 8553 9842 8554
rect 9702 8527 9815 8553
rect 9841 8527 9842 8553
rect 9702 8526 9842 8527
rect 9478 8415 9479 8441
rect 9505 8415 9506 8441
rect 9478 8409 9506 8415
rect 9590 8386 9618 8391
rect 9590 8339 9618 8358
rect 9702 8386 9730 8526
rect 9814 8521 9842 8526
rect 9422 8330 9450 8335
rect 9422 8329 9562 8330
rect 9422 8303 9423 8329
rect 9449 8303 9562 8329
rect 9422 8302 9562 8303
rect 9422 8297 9450 8302
rect 9534 8161 9562 8302
rect 9534 8135 9535 8161
rect 9561 8135 9562 8161
rect 9534 8129 9562 8135
rect 9702 8161 9730 8358
rect 9982 8498 10010 8503
rect 9982 8330 10010 8470
rect 10598 8497 10626 8503
rect 10598 8471 10599 8497
rect 10625 8471 10626 8497
rect 10486 8386 10514 8391
rect 10486 8339 10514 8358
rect 9982 8297 10010 8302
rect 9702 8135 9703 8161
rect 9729 8135 9730 8161
rect 9702 8129 9730 8135
rect 9590 7937 9618 7943
rect 9590 7911 9591 7937
rect 9617 7911 9618 7937
rect 9590 7322 9618 7911
rect 9918 7854 10050 7859
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 9918 7821 10050 7826
rect 9702 7658 9730 7663
rect 9702 7601 9730 7630
rect 10598 7658 10626 8471
rect 10654 8385 10682 8806
rect 10822 8801 10850 8806
rect 10654 8359 10655 8385
rect 10681 8359 10682 8385
rect 10654 8353 10682 8359
rect 10710 8721 10738 8727
rect 10710 8695 10711 8721
rect 10737 8695 10738 8721
rect 10710 8386 10738 8695
rect 10598 7625 10626 7630
rect 9702 7575 9703 7601
rect 9729 7575 9730 7601
rect 9702 7569 9730 7575
rect 10710 7574 10738 8358
rect 10766 8721 10794 8727
rect 10766 8695 10767 8721
rect 10793 8695 10794 8721
rect 10766 7713 10794 8695
rect 11662 8498 11690 9926
rect 11774 9617 11802 10094
rect 11886 10065 11914 11158
rect 12222 11153 12250 11158
rect 12390 10346 12418 13062
rect 12726 12810 12754 15946
rect 13230 14210 13258 14215
rect 12838 13594 12866 13599
rect 12838 13201 12866 13566
rect 13230 13594 13258 14182
rect 14294 14210 14322 18999
rect 17598 18438 17730 18443
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17598 18405 17730 18410
rect 17598 17654 17730 17659
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17598 17621 17730 17626
rect 17598 16870 17730 16875
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17598 16837 17730 16842
rect 17598 16086 17730 16091
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17598 16053 17730 16058
rect 17598 15302 17730 15307
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17598 15269 17730 15274
rect 17598 14518 17730 14523
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17598 14485 17730 14490
rect 14294 14177 14322 14182
rect 17598 13734 17730 13739
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17598 13701 17730 13706
rect 13230 13547 13258 13566
rect 12838 13175 12839 13201
rect 12865 13175 12866 13201
rect 12838 13169 12866 13175
rect 13454 13481 13482 13487
rect 13454 13455 13455 13481
rect 13481 13455 13482 13481
rect 12782 13146 12810 13151
rect 12782 13099 12810 13118
rect 12782 12810 12810 12815
rect 13454 12810 13482 13455
rect 18830 13146 18858 13151
rect 18718 13145 18858 13146
rect 18718 13119 18831 13145
rect 18857 13119 18858 13145
rect 18718 13118 18858 13119
rect 17598 12950 17730 12955
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17598 12917 17730 12922
rect 12726 12809 12810 12810
rect 12726 12783 12783 12809
rect 12809 12783 12810 12809
rect 12726 12782 12810 12783
rect 12726 12698 12754 12703
rect 12614 12026 12642 12031
rect 12614 11914 12642 11998
rect 12670 11914 12698 11919
rect 12614 11913 12698 11914
rect 12614 11887 12671 11913
rect 12697 11887 12698 11913
rect 12614 11886 12698 11887
rect 12446 11185 12474 11191
rect 12446 11159 12447 11185
rect 12473 11159 12474 11185
rect 12446 10458 12474 11159
rect 12446 10425 12474 10430
rect 12558 11185 12586 11191
rect 12558 11159 12559 11185
rect 12585 11159 12586 11185
rect 12390 10318 12474 10346
rect 12054 10122 12082 10127
rect 12278 10122 12306 10127
rect 12082 10094 12138 10122
rect 12054 10089 12082 10094
rect 11886 10039 11887 10065
rect 11913 10039 11914 10065
rect 11886 9674 11914 10039
rect 11886 9641 11914 9646
rect 11774 9591 11775 9617
rect 11801 9591 11802 9617
rect 11774 9585 11802 9591
rect 11942 9562 11970 9567
rect 11718 9450 11746 9455
rect 11718 8833 11746 9422
rect 11942 9394 11970 9534
rect 11998 9561 12026 9567
rect 11998 9535 11999 9561
rect 12025 9535 12026 9561
rect 11998 9506 12026 9535
rect 11998 9473 12026 9478
rect 12054 9394 12082 9399
rect 11942 9366 12026 9394
rect 11998 9338 12026 9366
rect 11718 8807 11719 8833
rect 11745 8807 11746 8833
rect 11718 8801 11746 8807
rect 11942 9281 11970 9287
rect 11942 9255 11943 9281
rect 11969 9255 11970 9281
rect 11662 8465 11690 8470
rect 11774 8721 11802 8727
rect 11774 8695 11775 8721
rect 11801 8695 11802 8721
rect 10766 7687 10767 7713
rect 10793 7687 10794 7713
rect 10766 7681 10794 7687
rect 11326 8330 11354 8335
rect 11326 7713 11354 8302
rect 11774 7770 11802 8695
rect 11830 8722 11858 8727
rect 11942 8722 11970 9255
rect 11830 8721 11970 8722
rect 11830 8695 11831 8721
rect 11857 8695 11970 8721
rect 11830 8694 11970 8695
rect 11830 8689 11858 8694
rect 11830 8497 11858 8503
rect 11830 8471 11831 8497
rect 11857 8471 11858 8497
rect 11830 8386 11858 8471
rect 11886 8442 11914 8694
rect 11886 8409 11914 8414
rect 11942 8610 11970 8615
rect 11830 8353 11858 8358
rect 11774 7737 11802 7742
rect 11942 8049 11970 8582
rect 11998 8553 12026 9310
rect 12054 8833 12082 9366
rect 12110 9337 12138 10094
rect 12278 10065 12306 10094
rect 12278 10039 12279 10065
rect 12305 10039 12306 10065
rect 12278 10033 12306 10039
rect 12390 10066 12418 10071
rect 12390 10019 12418 10038
rect 12222 10009 12250 10015
rect 12222 9983 12223 10009
rect 12249 9983 12250 10009
rect 12222 9506 12250 9983
rect 12222 9473 12250 9478
rect 12446 9505 12474 10318
rect 12558 10178 12586 11159
rect 12558 10145 12586 10150
rect 12446 9479 12447 9505
rect 12473 9479 12474 9505
rect 12446 9450 12474 9479
rect 12446 9417 12474 9422
rect 12502 10010 12530 10015
rect 12614 10010 12642 11886
rect 12670 11881 12698 11886
rect 12670 11802 12698 11807
rect 12670 11689 12698 11774
rect 12670 11663 12671 11689
rect 12697 11663 12698 11689
rect 12670 11657 12698 11663
rect 12726 11297 12754 12670
rect 12782 12418 12810 12782
rect 13398 12782 13482 12810
rect 12950 12698 12978 12703
rect 12950 12530 12978 12670
rect 13006 12642 13034 12647
rect 13230 12642 13258 12647
rect 13398 12642 13426 12782
rect 14630 12753 14658 12759
rect 14630 12727 14631 12753
rect 14657 12727 14658 12753
rect 13902 12698 13930 12703
rect 13902 12651 13930 12670
rect 13846 12642 13874 12647
rect 13034 12641 13426 12642
rect 13034 12615 13231 12641
rect 13257 12615 13426 12641
rect 13034 12614 13426 12615
rect 13006 12595 13034 12614
rect 13230 12609 13258 12614
rect 13118 12530 13146 12535
rect 12950 12502 13090 12530
rect 13062 12473 13090 12502
rect 13062 12447 13063 12473
rect 13089 12447 13090 12473
rect 13062 12441 13090 12447
rect 13118 12473 13146 12502
rect 13118 12447 13119 12473
rect 13145 12447 13146 12473
rect 13118 12441 13146 12447
rect 12782 12385 12810 12390
rect 12950 12361 12978 12367
rect 12950 12335 12951 12361
rect 12977 12335 12978 12361
rect 12950 12082 12978 12335
rect 13006 12362 13034 12367
rect 13006 12315 13034 12334
rect 13230 12362 13258 12367
rect 13230 12315 13258 12334
rect 13398 12361 13426 12614
rect 13790 12641 13874 12642
rect 13790 12615 13847 12641
rect 13873 12615 13874 12641
rect 13790 12614 13874 12615
rect 13790 12417 13818 12614
rect 13846 12609 13874 12614
rect 14630 12642 14658 12727
rect 14742 12698 14770 12703
rect 14742 12651 14770 12670
rect 18718 12698 18746 13118
rect 18830 13113 18858 13118
rect 19950 13089 19978 13095
rect 19950 13063 19951 13089
rect 19977 13063 19978 13089
rect 19950 12810 19978 13063
rect 19950 12777 19978 12782
rect 20006 12809 20034 12815
rect 20006 12783 20007 12809
rect 20033 12783 20034 12809
rect 18830 12754 18858 12759
rect 18830 12707 18858 12726
rect 18718 12665 18746 12670
rect 14630 12609 14658 12614
rect 14854 12642 14882 12647
rect 13790 12391 13791 12417
rect 13817 12391 13818 12417
rect 13790 12385 13818 12391
rect 13398 12335 13399 12361
rect 13425 12335 13426 12361
rect 12950 12054 13146 12082
rect 13006 11969 13034 11975
rect 13006 11943 13007 11969
rect 13033 11943 13034 11969
rect 12726 11271 12727 11297
rect 12753 11271 12754 11297
rect 12726 11265 12754 11271
rect 12782 11858 12810 11863
rect 12670 10906 12698 10911
rect 12782 10906 12810 11830
rect 13006 11802 13034 11943
rect 13006 11769 13034 11774
rect 13062 11858 13090 11863
rect 13062 11689 13090 11830
rect 13062 11663 13063 11689
rect 13089 11663 13090 11689
rect 13062 11657 13090 11663
rect 12670 10905 12810 10906
rect 12670 10879 12671 10905
rect 12697 10879 12810 10905
rect 12670 10878 12810 10879
rect 12838 11577 12866 11583
rect 12838 11551 12839 11577
rect 12865 11551 12866 11577
rect 12670 10873 12698 10878
rect 12614 9982 12698 10010
rect 12110 9311 12111 9337
rect 12137 9311 12138 9337
rect 12110 9305 12138 9311
rect 12502 9338 12530 9982
rect 12670 9954 12698 9982
rect 12726 10009 12754 10878
rect 12838 10066 12866 11551
rect 12950 11577 12978 11583
rect 12950 11551 12951 11577
rect 12977 11551 12978 11577
rect 12894 11522 12922 11527
rect 12894 11475 12922 11494
rect 12950 11466 12978 11551
rect 12950 11298 12978 11438
rect 12726 9983 12727 10009
rect 12753 9983 12754 10009
rect 12726 9977 12754 9983
rect 12782 10038 12838 10066
rect 12670 9921 12698 9926
rect 12614 9898 12642 9903
rect 12614 9851 12642 9870
rect 12614 9674 12642 9679
rect 12614 9627 12642 9646
rect 12222 9170 12250 9175
rect 12166 9114 12194 9119
rect 12166 8945 12194 9086
rect 12166 8919 12167 8945
rect 12193 8919 12194 8945
rect 12166 8913 12194 8919
rect 12222 8945 12250 9142
rect 12222 8919 12223 8945
rect 12249 8919 12250 8945
rect 12222 8913 12250 8919
rect 12334 9169 12362 9175
rect 12334 9143 12335 9169
rect 12361 9143 12362 9169
rect 12054 8807 12055 8833
rect 12081 8807 12082 8833
rect 12054 8801 12082 8807
rect 12334 8610 12362 9143
rect 12502 8833 12530 9310
rect 12670 9618 12698 9623
rect 12614 9226 12642 9231
rect 12670 9226 12698 9590
rect 12782 9281 12810 10038
rect 12838 10033 12866 10038
rect 12894 11270 12978 11298
rect 13006 11578 13034 11583
rect 12838 9954 12866 9959
rect 12838 9907 12866 9926
rect 12782 9255 12783 9281
rect 12809 9255 12810 9281
rect 12782 9249 12810 9255
rect 12614 9225 12698 9226
rect 12614 9199 12615 9225
rect 12641 9199 12698 9225
rect 12614 9198 12698 9199
rect 12614 9193 12642 9198
rect 12670 9170 12698 9198
rect 12894 9170 12922 11270
rect 12950 11186 12978 11191
rect 13006 11186 13034 11550
rect 12950 11185 13034 11186
rect 12950 11159 12951 11185
rect 12977 11159 13034 11185
rect 12950 11158 13034 11159
rect 12950 11153 12978 11158
rect 13062 11074 13090 11079
rect 13118 11074 13146 12054
rect 13062 11073 13146 11074
rect 13062 11047 13063 11073
rect 13089 11047 13146 11073
rect 13062 11046 13146 11047
rect 13062 11041 13090 11046
rect 13062 10682 13090 10687
rect 13062 10065 13090 10654
rect 13062 10039 13063 10065
rect 13089 10039 13090 10065
rect 13062 10033 13090 10039
rect 12950 10010 12978 10015
rect 12950 9963 12978 9982
rect 13006 9954 13034 9959
rect 13006 9907 13034 9926
rect 12950 9450 12978 9455
rect 12950 9281 12978 9422
rect 13006 9394 13034 9399
rect 13118 9394 13146 11046
rect 13286 11858 13314 11863
rect 13398 11858 13426 12335
rect 13846 12362 13874 12367
rect 13846 11969 13874 12334
rect 14854 12305 14882 12614
rect 20006 12474 20034 12783
rect 20006 12441 20034 12446
rect 14854 12279 14855 12305
rect 14881 12279 14882 12305
rect 14854 12273 14882 12279
rect 17598 12166 17730 12171
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17598 12133 17730 12138
rect 20006 12025 20034 12031
rect 20006 11999 20007 12025
rect 20033 11999 20034 12025
rect 13846 11943 13847 11969
rect 13873 11943 13874 11969
rect 13846 11937 13874 11943
rect 13902 11970 13930 11975
rect 13902 11913 13930 11942
rect 13902 11887 13903 11913
rect 13929 11887 13930 11913
rect 13902 11881 13930 11887
rect 14742 11970 14770 11975
rect 13286 11857 13426 11858
rect 13286 11831 13287 11857
rect 13313 11831 13426 11857
rect 13286 11830 13426 11831
rect 14014 11858 14042 11863
rect 13286 11802 13314 11830
rect 14014 11811 14042 11830
rect 13286 11577 13314 11774
rect 13286 11551 13287 11577
rect 13313 11551 13314 11577
rect 13286 10737 13314 11551
rect 13678 11522 13706 11527
rect 13678 11475 13706 11494
rect 14742 11521 14770 11942
rect 18830 11970 18858 11975
rect 18830 11923 18858 11942
rect 20006 11802 20034 11999
rect 20006 11769 20034 11774
rect 14742 11495 14743 11521
rect 14769 11495 14770 11521
rect 14742 11489 14770 11495
rect 17598 11382 17730 11387
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17598 11349 17730 11354
rect 18830 10793 18858 10799
rect 18830 10767 18831 10793
rect 18857 10767 18858 10793
rect 13286 10711 13287 10737
rect 13313 10711 13314 10737
rect 13286 10346 13314 10711
rect 14574 10737 14602 10743
rect 14574 10711 14575 10737
rect 14601 10711 14602 10737
rect 14518 10682 14546 10687
rect 14518 10635 14546 10654
rect 13342 10346 13370 10351
rect 13286 10345 13370 10346
rect 13286 10319 13343 10345
rect 13369 10319 13370 10345
rect 13286 10318 13370 10319
rect 13174 10066 13202 10071
rect 13174 9729 13202 10038
rect 13174 9703 13175 9729
rect 13201 9703 13202 9729
rect 13174 9697 13202 9703
rect 13342 10010 13370 10318
rect 14574 10094 14602 10711
rect 17598 10598 17730 10603
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17598 10565 17730 10570
rect 14910 10122 14938 10127
rect 14574 10066 14938 10094
rect 18830 10122 18858 10767
rect 20006 10681 20034 10687
rect 20006 10655 20007 10681
rect 20033 10655 20034 10681
rect 20006 10458 20034 10655
rect 20006 10425 20034 10430
rect 18830 10089 18858 10094
rect 20118 10289 20146 10295
rect 20118 10263 20119 10289
rect 20145 10263 20146 10289
rect 20118 10122 20146 10263
rect 20118 10089 20146 10094
rect 13454 10010 13482 10015
rect 13342 10009 13482 10010
rect 13342 9983 13455 10009
rect 13481 9983 13482 10009
rect 13342 9982 13482 9983
rect 13286 9674 13314 9679
rect 13286 9627 13314 9646
rect 13034 9366 13146 9394
rect 13006 9337 13034 9366
rect 13006 9311 13007 9337
rect 13033 9311 13034 9337
rect 13006 9305 13034 9311
rect 12950 9255 12951 9281
rect 12977 9255 12978 9281
rect 12950 9249 12978 9255
rect 13342 9226 13370 9982
rect 13454 9977 13482 9982
rect 13846 9954 13874 9959
rect 13846 9907 13874 9926
rect 14910 9953 14938 10066
rect 14910 9927 14911 9953
rect 14937 9927 14938 9953
rect 14910 9921 14938 9927
rect 18830 10009 18858 10015
rect 18830 9983 18831 10009
rect 18857 9983 18858 10009
rect 17598 9814 17730 9819
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17598 9781 17730 9786
rect 13398 9617 13426 9623
rect 13398 9591 13399 9617
rect 13425 9591 13426 9617
rect 13398 9394 13426 9591
rect 14294 9562 14322 9567
rect 14294 9515 14322 9534
rect 14798 9562 14826 9567
rect 13398 9361 13426 9366
rect 13510 9505 13538 9511
rect 13510 9479 13511 9505
rect 13537 9479 13538 9505
rect 13510 9282 13538 9479
rect 13566 9505 13594 9511
rect 13566 9479 13567 9505
rect 13593 9479 13594 9505
rect 13566 9338 13594 9479
rect 13622 9506 13650 9511
rect 14238 9506 14266 9511
rect 13622 9505 14266 9506
rect 13622 9479 13623 9505
rect 13649 9479 14239 9505
rect 14265 9479 14266 9505
rect 13622 9478 14266 9479
rect 13622 9473 13650 9478
rect 14238 9473 14266 9478
rect 13566 9310 13762 9338
rect 13510 9249 13538 9254
rect 13734 9281 13762 9310
rect 13734 9255 13735 9281
rect 13761 9255 13762 9281
rect 13734 9249 13762 9255
rect 13398 9226 13426 9231
rect 13342 9225 13426 9226
rect 13342 9199 13399 9225
rect 13425 9199 13426 9225
rect 13342 9198 13426 9199
rect 12670 9142 12922 9170
rect 12614 9114 12642 9119
rect 13006 9114 13034 9119
rect 12614 9067 12642 9086
rect 12894 9113 13034 9114
rect 12894 9087 13007 9113
rect 13033 9087 13034 9113
rect 12894 9086 13034 9087
rect 12670 8890 12698 8895
rect 12670 8843 12698 8862
rect 12502 8807 12503 8833
rect 12529 8807 12530 8833
rect 12502 8801 12530 8807
rect 12838 8834 12866 8839
rect 12614 8778 12642 8783
rect 12614 8731 12642 8750
rect 12390 8722 12418 8727
rect 12390 8675 12418 8694
rect 12334 8577 12362 8582
rect 12838 8610 12866 8806
rect 12838 8577 12866 8582
rect 12894 8722 12922 9086
rect 13006 9081 13034 9086
rect 13230 8890 13258 8895
rect 13230 8843 13258 8862
rect 13398 8834 13426 9198
rect 14798 9169 14826 9534
rect 18830 9562 18858 9983
rect 20006 9897 20034 9903
rect 20006 9871 20007 9897
rect 20033 9871 20034 9897
rect 20006 9786 20034 9871
rect 20006 9753 20034 9758
rect 18830 9529 18858 9534
rect 14798 9143 14799 9169
rect 14825 9143 14826 9169
rect 14798 9137 14826 9143
rect 17598 9030 17730 9035
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17598 8997 17730 9002
rect 13958 8890 13986 8895
rect 13426 8806 13538 8834
rect 13398 8801 13426 8806
rect 11998 8527 11999 8553
rect 12025 8527 12026 8553
rect 11998 8521 12026 8527
rect 12726 8497 12754 8503
rect 12726 8471 12727 8497
rect 12753 8471 12754 8497
rect 12614 8441 12642 8447
rect 12614 8415 12615 8441
rect 12641 8415 12642 8441
rect 12334 8386 12362 8391
rect 12334 8105 12362 8358
rect 12334 8079 12335 8105
rect 12361 8079 12362 8105
rect 12334 8073 12362 8079
rect 12614 8330 12642 8415
rect 12670 8386 12698 8391
rect 12670 8339 12698 8358
rect 11942 8023 11943 8049
rect 11969 8023 11970 8049
rect 11326 7687 11327 7713
rect 11353 7687 11354 7713
rect 11326 7681 11354 7687
rect 11438 7713 11466 7719
rect 11438 7687 11439 7713
rect 11465 7687 11466 7713
rect 10934 7658 10962 7663
rect 10878 7602 10906 7607
rect 10710 7546 10794 7574
rect 9758 7322 9786 7327
rect 10710 7322 10738 7327
rect 9590 7321 9786 7322
rect 9590 7295 9759 7321
rect 9785 7295 9786 7321
rect 9590 7294 9786 7295
rect 8750 7233 8778 7238
rect 2238 6678 2370 6683
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2238 6645 2370 6650
rect 2238 5894 2370 5899
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2238 5861 2370 5866
rect 2238 5110 2370 5115
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2238 5077 2370 5082
rect 2238 4326 2370 4331
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2238 4293 2370 4298
rect 9758 4214 9786 7294
rect 10206 7321 10738 7322
rect 10206 7295 10711 7321
rect 10737 7295 10738 7321
rect 10206 7294 10738 7295
rect 9982 7266 10010 7271
rect 9982 7219 10010 7238
rect 9918 7070 10050 7075
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 9918 7037 10050 7042
rect 10206 6929 10234 7294
rect 10710 7289 10738 7294
rect 10766 7209 10794 7546
rect 10878 7377 10906 7574
rect 10878 7351 10879 7377
rect 10905 7351 10906 7377
rect 10878 7345 10906 7351
rect 10766 7183 10767 7209
rect 10793 7183 10794 7209
rect 10766 7177 10794 7183
rect 10206 6903 10207 6929
rect 10233 6903 10234 6929
rect 10206 6897 10234 6903
rect 9870 6874 9898 6879
rect 9870 6827 9898 6846
rect 9918 6286 10050 6291
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 9918 6253 10050 6258
rect 9918 5502 10050 5507
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 9918 5469 10050 5474
rect 9918 4718 10050 4723
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 9918 4685 10050 4690
rect 9422 4186 9786 4214
rect 2238 3542 2370 3547
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2238 3509 2370 3514
rect 2238 2758 2370 2763
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2238 2725 2370 2730
rect 9422 2169 9450 4186
rect 9918 3934 10050 3939
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 9918 3901 10050 3906
rect 9918 3150 10050 3155
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 9918 3117 10050 3122
rect 9918 2366 10050 2371
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 9918 2333 10050 2338
rect 9422 2143 9423 2169
rect 9449 2143 9450 2169
rect 9422 2137 9450 2143
rect 10934 2169 10962 7630
rect 11158 7657 11186 7663
rect 11158 7631 11159 7657
rect 11185 7631 11186 7657
rect 11158 6874 11186 7631
rect 11382 7602 11410 7621
rect 11382 7569 11410 7574
rect 11158 6841 11186 6846
rect 11270 6817 11298 6823
rect 11270 6791 11271 6817
rect 11297 6791 11298 6817
rect 11270 6762 11298 6791
rect 11438 6762 11466 7687
rect 11718 7601 11746 7607
rect 11718 7575 11719 7601
rect 11745 7575 11746 7601
rect 11718 7266 11746 7575
rect 11830 7266 11858 7271
rect 11942 7266 11970 8023
rect 12614 7769 12642 8302
rect 12726 8050 12754 8471
rect 12838 8442 12866 8447
rect 12894 8442 12922 8694
rect 12838 8441 12922 8442
rect 12838 8415 12839 8441
rect 12865 8415 12922 8441
rect 12838 8414 12922 8415
rect 12950 8498 12978 8503
rect 12950 8441 12978 8470
rect 12950 8415 12951 8441
rect 12977 8415 12978 8441
rect 12838 8409 12866 8414
rect 12950 8409 12978 8415
rect 13398 8105 13426 8111
rect 13398 8079 13399 8105
rect 13425 8079 13426 8105
rect 12726 8022 13090 8050
rect 12614 7743 12615 7769
rect 12641 7743 12642 7769
rect 12614 7737 12642 7743
rect 12838 7770 12866 7775
rect 12838 7723 12866 7742
rect 13062 7769 13090 8022
rect 13062 7743 13063 7769
rect 13089 7743 13090 7769
rect 13062 7737 13090 7743
rect 12726 7657 12754 7663
rect 12726 7631 12727 7657
rect 12753 7631 12754 7657
rect 12222 7602 12250 7607
rect 12222 7321 12250 7574
rect 12670 7602 12698 7621
rect 12670 7569 12698 7574
rect 12726 7574 12754 7631
rect 13118 7602 13146 7621
rect 12726 7546 12866 7574
rect 13118 7569 13146 7574
rect 13398 7602 13426 8079
rect 13398 7569 13426 7574
rect 13510 8106 13538 8806
rect 13902 8778 13930 8783
rect 13902 8553 13930 8750
rect 13902 8527 13903 8553
rect 13929 8527 13930 8553
rect 13902 8521 13930 8527
rect 13958 8497 13986 8862
rect 14294 8890 14322 8895
rect 14294 8843 14322 8862
rect 20006 8889 20034 8895
rect 20006 8863 20007 8889
rect 20033 8863 20034 8889
rect 14630 8834 14658 8839
rect 14630 8787 14658 8806
rect 18830 8834 18858 8839
rect 18830 8787 18858 8806
rect 20006 8778 20034 8863
rect 20006 8745 20034 8750
rect 13958 8471 13959 8497
rect 13985 8471 13986 8497
rect 13958 8465 13986 8471
rect 18830 8441 18858 8447
rect 18830 8415 18831 8441
rect 18857 8415 18858 8441
rect 17598 8246 17730 8251
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17598 8213 17730 8218
rect 13622 8106 13650 8111
rect 13510 8105 13650 8106
rect 13510 8079 13623 8105
rect 13649 8079 13650 8105
rect 13510 8078 13650 8079
rect 12222 7295 12223 7321
rect 12249 7295 12250 7321
rect 12222 7289 12250 7295
rect 11718 7265 11970 7266
rect 11718 7239 11831 7265
rect 11857 7239 11970 7265
rect 11718 7238 11970 7239
rect 11494 6874 11522 6879
rect 11494 6827 11522 6846
rect 11830 6874 11858 7238
rect 12838 6985 12866 7546
rect 12838 6959 12839 6985
rect 12865 6959 12866 6985
rect 12838 6953 12866 6959
rect 13286 7321 13314 7327
rect 13286 7295 13287 7321
rect 13313 7295 13314 7321
rect 11830 6841 11858 6846
rect 12894 6818 12922 6823
rect 13286 6818 13314 7295
rect 13510 7321 13538 8078
rect 13622 8073 13650 8078
rect 18830 7602 18858 8415
rect 20006 8329 20034 8335
rect 20006 8303 20007 8329
rect 20033 8303 20034 8329
rect 20006 8106 20034 8303
rect 20006 8073 20034 8078
rect 18830 7569 18858 7574
rect 17598 7462 17730 7467
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17598 7429 17730 7434
rect 13510 7295 13511 7321
rect 13537 7295 13538 7321
rect 13510 7289 13538 7295
rect 12894 6817 13314 6818
rect 12894 6791 12895 6817
rect 12921 6791 13314 6817
rect 12894 6790 13314 6791
rect 11494 6762 11522 6767
rect 11438 6734 11494 6762
rect 11270 6729 11298 6734
rect 11494 6729 11522 6734
rect 11942 6762 11970 6767
rect 10934 2143 10935 2169
rect 10961 2143 10962 2169
rect 10934 2137 10962 2143
rect 9926 2058 9954 2063
rect 9758 2057 9954 2058
rect 9758 2031 9927 2057
rect 9953 2031 9954 2057
rect 9758 2030 9954 2031
rect 2238 1974 2370 1979
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2238 1941 2370 1946
rect 9198 1666 9226 1671
rect 9086 1665 9226 1666
rect 9086 1639 9199 1665
rect 9225 1639 9226 1665
rect 9086 1638 9226 1639
rect 9086 400 9114 1638
rect 9198 1633 9226 1638
rect 9758 400 9786 2030
rect 9926 2025 9954 2030
rect 10766 2058 10794 2063
rect 9918 1582 10050 1587
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 9918 1549 10050 1554
rect 10766 400 10794 2030
rect 11382 2058 11410 2063
rect 11382 2011 11410 2030
rect 11942 1777 11970 6734
rect 12894 4214 12922 6790
rect 17598 6678 17730 6683
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17598 6645 17730 6650
rect 17598 5894 17730 5899
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17598 5861 17730 5866
rect 17598 5110 17730 5115
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17598 5077 17730 5082
rect 17598 4326 17730 4331
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17598 4293 17730 4298
rect 12894 4186 13258 4214
rect 13230 2169 13258 4186
rect 17598 3542 17730 3547
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17598 3509 17730 3514
rect 17598 2758 17730 2763
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17598 2725 17730 2730
rect 13230 2143 13231 2169
rect 13257 2143 13258 2169
rect 13230 2137 13258 2143
rect 11942 1751 11943 1777
rect 11969 1751 11970 1777
rect 11942 1745 11970 1751
rect 13118 2058 13146 2063
rect 11102 1721 11130 1727
rect 11102 1695 11103 1721
rect 11129 1695 11130 1721
rect 11102 400 11130 1695
rect 13118 400 13146 2030
rect 13734 2058 13762 2063
rect 13734 2011 13762 2030
rect 17598 1974 17730 1979
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17598 1941 17730 1946
rect 9072 0 9128 400
rect 9744 0 9800 400
rect 10752 0 10808 400
rect 11088 0 11144 400
rect 13104 0 13160 400
<< via2 >>
rect 2238 19221 2266 19222
rect 2238 19195 2239 19221
rect 2239 19195 2265 19221
rect 2265 19195 2266 19221
rect 2238 19194 2266 19195
rect 2290 19221 2318 19222
rect 2290 19195 2291 19221
rect 2291 19195 2317 19221
rect 2317 19195 2318 19221
rect 2290 19194 2318 19195
rect 2342 19221 2370 19222
rect 2342 19195 2343 19221
rect 2343 19195 2369 19221
rect 2369 19195 2370 19221
rect 2342 19194 2370 19195
rect 8414 19110 8442 19138
rect 9030 19137 9058 19138
rect 9030 19111 9031 19137
rect 9031 19111 9057 19137
rect 9057 19111 9058 19137
rect 9030 19110 9058 19111
rect 2238 18437 2266 18438
rect 2238 18411 2239 18437
rect 2239 18411 2265 18437
rect 2265 18411 2266 18437
rect 2238 18410 2266 18411
rect 2290 18437 2318 18438
rect 2290 18411 2291 18437
rect 2291 18411 2317 18437
rect 2317 18411 2318 18437
rect 2290 18410 2318 18411
rect 2342 18437 2370 18438
rect 2342 18411 2343 18437
rect 2343 18411 2369 18437
rect 2369 18411 2370 18437
rect 2342 18410 2370 18411
rect 2238 17653 2266 17654
rect 2238 17627 2239 17653
rect 2239 17627 2265 17653
rect 2265 17627 2266 17653
rect 2238 17626 2266 17627
rect 2290 17653 2318 17654
rect 2290 17627 2291 17653
rect 2291 17627 2317 17653
rect 2317 17627 2318 17653
rect 2290 17626 2318 17627
rect 2342 17653 2370 17654
rect 2342 17627 2343 17653
rect 2343 17627 2369 17653
rect 2369 17627 2370 17653
rect 2342 17626 2370 17627
rect 2238 16869 2266 16870
rect 2238 16843 2239 16869
rect 2239 16843 2265 16869
rect 2265 16843 2266 16869
rect 2238 16842 2266 16843
rect 2290 16869 2318 16870
rect 2290 16843 2291 16869
rect 2291 16843 2317 16869
rect 2317 16843 2318 16869
rect 2290 16842 2318 16843
rect 2342 16869 2370 16870
rect 2342 16843 2343 16869
rect 2343 16843 2369 16869
rect 2369 16843 2370 16869
rect 2342 16842 2370 16843
rect 2238 16085 2266 16086
rect 2238 16059 2239 16085
rect 2239 16059 2265 16085
rect 2265 16059 2266 16085
rect 2238 16058 2266 16059
rect 2290 16085 2318 16086
rect 2290 16059 2291 16085
rect 2291 16059 2317 16085
rect 2317 16059 2318 16085
rect 2290 16058 2318 16059
rect 2342 16085 2370 16086
rect 2342 16059 2343 16085
rect 2343 16059 2369 16085
rect 2369 16059 2370 16085
rect 2342 16058 2370 16059
rect 2238 15301 2266 15302
rect 2238 15275 2239 15301
rect 2239 15275 2265 15301
rect 2265 15275 2266 15301
rect 2238 15274 2266 15275
rect 2290 15301 2318 15302
rect 2290 15275 2291 15301
rect 2291 15275 2317 15301
rect 2317 15275 2318 15301
rect 2290 15274 2318 15275
rect 2342 15301 2370 15302
rect 2342 15275 2343 15301
rect 2343 15275 2369 15301
rect 2369 15275 2370 15301
rect 2342 15274 2370 15275
rect 2238 14517 2266 14518
rect 2238 14491 2239 14517
rect 2239 14491 2265 14517
rect 2265 14491 2266 14517
rect 2238 14490 2266 14491
rect 2290 14517 2318 14518
rect 2290 14491 2291 14517
rect 2291 14491 2317 14517
rect 2317 14491 2318 14517
rect 2290 14490 2318 14491
rect 2342 14517 2370 14518
rect 2342 14491 2343 14517
rect 2343 14491 2369 14517
rect 2369 14491 2370 14517
rect 2342 14490 2370 14491
rect 7630 14294 7658 14322
rect 8134 14321 8162 14322
rect 8134 14295 8135 14321
rect 8135 14295 8161 14321
rect 8161 14295 8162 14321
rect 8134 14294 8162 14295
rect 8414 14294 8442 14322
rect 2086 14126 2114 14154
rect 966 12782 994 12810
rect 966 11774 994 11802
rect 966 11241 994 11242
rect 966 11215 967 11241
rect 967 11215 993 11241
rect 993 11215 994 11241
rect 966 11214 994 11215
rect 2238 13733 2266 13734
rect 2238 13707 2239 13733
rect 2239 13707 2265 13733
rect 2265 13707 2266 13733
rect 2238 13706 2266 13707
rect 2290 13733 2318 13734
rect 2290 13707 2291 13733
rect 2291 13707 2317 13733
rect 2317 13707 2318 13733
rect 2290 13706 2318 13707
rect 2342 13733 2370 13734
rect 2342 13707 2343 13733
rect 2343 13707 2369 13733
rect 2369 13707 2370 13733
rect 2342 13706 2370 13707
rect 8470 14265 8498 14266
rect 8470 14239 8471 14265
rect 8471 14239 8497 14265
rect 8497 14239 8498 14265
rect 8470 14238 8498 14239
rect 2142 13145 2170 13146
rect 2142 13119 2143 13145
rect 2143 13119 2169 13145
rect 2169 13119 2170 13145
rect 2142 13118 2170 13119
rect 5502 13118 5530 13146
rect 6790 13118 6818 13146
rect 6566 13006 6594 13034
rect 2238 12949 2266 12950
rect 2238 12923 2239 12949
rect 2239 12923 2265 12949
rect 2265 12923 2266 12949
rect 2238 12922 2266 12923
rect 2290 12949 2318 12950
rect 2290 12923 2291 12949
rect 2291 12923 2317 12949
rect 2317 12923 2318 12949
rect 2290 12922 2318 12923
rect 2342 12949 2370 12950
rect 2342 12923 2343 12949
rect 2343 12923 2369 12949
rect 2369 12923 2370 12949
rect 2342 12922 2370 12923
rect 6510 12473 6538 12474
rect 6510 12447 6511 12473
rect 6511 12447 6537 12473
rect 6537 12447 6538 12473
rect 6510 12446 6538 12447
rect 2238 12165 2266 12166
rect 2238 12139 2239 12165
rect 2239 12139 2265 12165
rect 2265 12139 2266 12165
rect 2238 12138 2266 12139
rect 2290 12165 2318 12166
rect 2290 12139 2291 12165
rect 2291 12139 2317 12165
rect 2317 12139 2318 12165
rect 2290 12138 2318 12139
rect 2342 12165 2370 12166
rect 2342 12139 2343 12165
rect 2343 12139 2369 12165
rect 2369 12139 2370 12165
rect 2342 12138 2370 12139
rect 2142 11969 2170 11970
rect 2142 11943 2143 11969
rect 2143 11943 2169 11969
rect 2169 11943 2170 11969
rect 2142 11942 2170 11943
rect 7406 13230 7434 13258
rect 10094 19110 10122 19138
rect 10878 19137 10906 19138
rect 10878 19111 10879 19137
rect 10879 19111 10905 19137
rect 10905 19111 10906 19137
rect 10878 19110 10906 19111
rect 11438 19110 11466 19138
rect 9918 18829 9946 18830
rect 9918 18803 9919 18829
rect 9919 18803 9945 18829
rect 9945 18803 9946 18829
rect 9918 18802 9946 18803
rect 9970 18829 9998 18830
rect 9970 18803 9971 18829
rect 9971 18803 9997 18829
rect 9997 18803 9998 18829
rect 9970 18802 9998 18803
rect 10022 18829 10050 18830
rect 10022 18803 10023 18829
rect 10023 18803 10049 18829
rect 10049 18803 10050 18829
rect 10022 18802 10050 18803
rect 9422 18718 9450 18746
rect 10038 18745 10066 18746
rect 10038 18719 10039 18745
rect 10039 18719 10065 18745
rect 10065 18719 10066 18745
rect 10038 18718 10066 18719
rect 9918 18045 9946 18046
rect 9918 18019 9919 18045
rect 9919 18019 9945 18045
rect 9945 18019 9946 18045
rect 9918 18018 9946 18019
rect 9970 18045 9998 18046
rect 9970 18019 9971 18045
rect 9971 18019 9997 18045
rect 9997 18019 9998 18045
rect 9970 18018 9998 18019
rect 10022 18045 10050 18046
rect 10022 18019 10023 18045
rect 10023 18019 10049 18045
rect 10049 18019 10050 18045
rect 10022 18018 10050 18019
rect 9918 17261 9946 17262
rect 9918 17235 9919 17261
rect 9919 17235 9945 17261
rect 9945 17235 9946 17261
rect 9918 17234 9946 17235
rect 9970 17261 9998 17262
rect 9970 17235 9971 17261
rect 9971 17235 9997 17261
rect 9997 17235 9998 17261
rect 9970 17234 9998 17235
rect 10022 17261 10050 17262
rect 10022 17235 10023 17261
rect 10023 17235 10049 17261
rect 10049 17235 10050 17261
rect 10022 17234 10050 17235
rect 9918 16477 9946 16478
rect 9918 16451 9919 16477
rect 9919 16451 9945 16477
rect 9945 16451 9946 16477
rect 9918 16450 9946 16451
rect 9970 16477 9998 16478
rect 9970 16451 9971 16477
rect 9971 16451 9997 16477
rect 9997 16451 9998 16477
rect 9970 16450 9998 16451
rect 10022 16477 10050 16478
rect 10022 16451 10023 16477
rect 10023 16451 10049 16477
rect 10049 16451 10050 16477
rect 10022 16450 10050 16451
rect 12782 19278 12810 19306
rect 12782 19137 12810 19138
rect 12782 19111 12783 19137
rect 12783 19111 12809 19137
rect 12809 19111 12810 19137
rect 12782 19110 12810 19111
rect 13118 19110 13146 19138
rect 13398 19278 13426 19306
rect 17598 19221 17626 19222
rect 17598 19195 17599 19221
rect 17599 19195 17625 19221
rect 17625 19195 17626 19221
rect 17598 19194 17626 19195
rect 17650 19221 17678 19222
rect 17650 19195 17651 19221
rect 17651 19195 17677 19221
rect 17677 19195 17678 19221
rect 17650 19194 17678 19195
rect 17702 19221 17730 19222
rect 17702 19195 17703 19221
rect 17703 19195 17729 19221
rect 17729 19195 17730 19221
rect 17702 19194 17730 19195
rect 14686 19137 14714 19138
rect 14686 19111 14687 19137
rect 14687 19111 14713 19137
rect 14713 19111 14714 19137
rect 14686 19110 14714 19111
rect 9918 15693 9946 15694
rect 9918 15667 9919 15693
rect 9919 15667 9945 15693
rect 9945 15667 9946 15693
rect 9918 15666 9946 15667
rect 9970 15693 9998 15694
rect 9970 15667 9971 15693
rect 9971 15667 9997 15693
rect 9997 15667 9998 15693
rect 9970 15666 9998 15667
rect 10022 15693 10050 15694
rect 10022 15667 10023 15693
rect 10023 15667 10049 15693
rect 10049 15667 10050 15693
rect 10022 15666 10050 15667
rect 9918 14909 9946 14910
rect 9918 14883 9919 14909
rect 9919 14883 9945 14909
rect 9945 14883 9946 14909
rect 9918 14882 9946 14883
rect 9970 14909 9998 14910
rect 9970 14883 9971 14909
rect 9971 14883 9997 14909
rect 9997 14883 9998 14909
rect 9970 14882 9998 14883
rect 10022 14909 10050 14910
rect 10022 14883 10023 14909
rect 10023 14883 10049 14909
rect 10049 14883 10050 14909
rect 10022 14882 10050 14883
rect 8918 14294 8946 14322
rect 8974 14238 9002 14266
rect 7910 13257 7938 13258
rect 7910 13231 7911 13257
rect 7911 13231 7937 13257
rect 7937 13231 7938 13257
rect 7910 13230 7938 13231
rect 7182 13033 7210 13034
rect 7182 13007 7183 13033
rect 7183 13007 7209 13033
rect 7209 13007 7210 13033
rect 7182 13006 7210 13007
rect 7966 13089 7994 13090
rect 7966 13063 7967 13089
rect 7967 13063 7993 13089
rect 7993 13063 7994 13089
rect 7966 13062 7994 13063
rect 7294 12726 7322 12754
rect 6846 12446 6874 12474
rect 6734 12390 6762 12418
rect 7126 12390 7154 12418
rect 4942 11886 4970 11914
rect 6006 11774 6034 11802
rect 2238 11381 2266 11382
rect 2238 11355 2239 11381
rect 2239 11355 2265 11381
rect 2265 11355 2266 11381
rect 2238 11354 2266 11355
rect 2290 11381 2318 11382
rect 2290 11355 2291 11381
rect 2291 11355 2317 11381
rect 2317 11355 2318 11381
rect 2290 11354 2318 11355
rect 2342 11381 2370 11382
rect 2342 11355 2343 11381
rect 2343 11355 2369 11381
rect 2369 11355 2370 11381
rect 2342 11354 2370 11355
rect 2142 11185 2170 11186
rect 2142 11159 2143 11185
rect 2143 11159 2169 11185
rect 2169 11159 2170 11185
rect 2142 11158 2170 11159
rect 5670 11158 5698 11186
rect 5670 10822 5698 10850
rect 2086 10766 2114 10794
rect 966 10430 994 10458
rect 2238 10597 2266 10598
rect 2238 10571 2239 10597
rect 2239 10571 2265 10597
rect 2265 10571 2266 10597
rect 2238 10570 2266 10571
rect 2290 10597 2318 10598
rect 2290 10571 2291 10597
rect 2291 10571 2317 10597
rect 2317 10571 2318 10597
rect 2290 10570 2318 10571
rect 2342 10597 2370 10598
rect 2342 10571 2343 10597
rect 2343 10571 2369 10597
rect 2369 10571 2370 10597
rect 2342 10570 2370 10571
rect 6790 11913 6818 11914
rect 6790 11887 6791 11913
rect 6791 11887 6817 11913
rect 6817 11887 6818 11913
rect 6790 11886 6818 11887
rect 6286 11633 6314 11634
rect 6286 11607 6287 11633
rect 6287 11607 6313 11633
rect 6313 11607 6314 11633
rect 6286 11606 6314 11607
rect 6846 11774 6874 11802
rect 7014 11606 7042 11634
rect 7014 11185 7042 11186
rect 7014 11159 7015 11185
rect 7015 11159 7041 11185
rect 7041 11159 7042 11185
rect 7014 11158 7042 11159
rect 7238 12446 7266 12474
rect 8078 12222 8106 12250
rect 9254 13873 9282 13874
rect 9254 13847 9255 13873
rect 9255 13847 9281 13873
rect 9281 13847 9282 13873
rect 9254 13846 9282 13847
rect 9758 14321 9786 14322
rect 9758 14295 9759 14321
rect 9759 14295 9785 14321
rect 9785 14295 9786 14321
rect 9758 14294 9786 14295
rect 9918 14125 9946 14126
rect 9918 14099 9919 14125
rect 9919 14099 9945 14125
rect 9945 14099 9946 14125
rect 9918 14098 9946 14099
rect 9970 14125 9998 14126
rect 9970 14099 9971 14125
rect 9971 14099 9997 14125
rect 9997 14099 9998 14125
rect 9970 14098 9998 14099
rect 10022 14125 10050 14126
rect 10022 14099 10023 14125
rect 10023 14099 10049 14125
rect 10049 14099 10050 14125
rect 10022 14098 10050 14099
rect 9590 13846 9618 13874
rect 8806 13257 8834 13258
rect 8806 13231 8807 13257
rect 8807 13231 8833 13257
rect 8833 13231 8834 13257
rect 8806 13230 8834 13231
rect 8862 13089 8890 13090
rect 8862 13063 8863 13089
rect 8863 13063 8889 13089
rect 8889 13063 8890 13089
rect 8862 13062 8890 13063
rect 9030 13145 9058 13146
rect 9030 13119 9031 13145
rect 9031 13119 9057 13145
rect 9057 13119 9058 13145
rect 9030 13118 9058 13119
rect 10710 14321 10738 14322
rect 10710 14295 10711 14321
rect 10711 14295 10737 14321
rect 10737 14295 10738 14321
rect 10710 14294 10738 14295
rect 11830 14294 11858 14322
rect 11270 14041 11298 14042
rect 11270 14015 11271 14041
rect 11271 14015 11297 14041
rect 11297 14015 11298 14041
rect 11270 14014 11298 14015
rect 10766 13985 10794 13986
rect 10766 13959 10767 13985
rect 10767 13959 10793 13985
rect 10793 13959 10794 13985
rect 10766 13958 10794 13959
rect 11158 13985 11186 13986
rect 11158 13959 11159 13985
rect 11159 13959 11185 13985
rect 11185 13959 11186 13985
rect 11158 13958 11186 13959
rect 9478 13537 9506 13538
rect 9478 13511 9479 13537
rect 9479 13511 9505 13537
rect 9505 13511 9506 13537
rect 9478 13510 9506 13511
rect 9366 13257 9394 13258
rect 9366 13231 9367 13257
rect 9367 13231 9393 13257
rect 9393 13231 9394 13257
rect 9366 13230 9394 13231
rect 9918 13341 9946 13342
rect 9918 13315 9919 13341
rect 9919 13315 9945 13341
rect 9945 13315 9946 13341
rect 9918 13314 9946 13315
rect 9970 13341 9998 13342
rect 9970 13315 9971 13341
rect 9971 13315 9997 13341
rect 9997 13315 9998 13341
rect 9970 13314 9998 13315
rect 10022 13341 10050 13342
rect 10022 13315 10023 13341
rect 10023 13315 10049 13341
rect 10049 13315 10050 13341
rect 10022 13314 10050 13315
rect 9982 13257 10010 13258
rect 9982 13231 9983 13257
rect 9983 13231 10009 13257
rect 10009 13231 10010 13257
rect 9982 13230 10010 13231
rect 11326 13929 11354 13930
rect 11326 13903 11327 13929
rect 11327 13903 11353 13929
rect 11353 13903 11354 13929
rect 11326 13902 11354 13903
rect 11326 13510 11354 13538
rect 12334 14321 12362 14322
rect 12334 14295 12335 14321
rect 12335 14295 12361 14321
rect 12361 14295 12362 14321
rect 12334 14294 12362 14295
rect 12110 14014 12138 14042
rect 10318 13230 10346 13258
rect 9198 12614 9226 12642
rect 9422 13118 9450 13146
rect 9758 13145 9786 13146
rect 9758 13119 9759 13145
rect 9759 13119 9785 13145
rect 9785 13119 9786 13145
rect 9758 13118 9786 13119
rect 8918 12222 8946 12250
rect 8694 12025 8722 12026
rect 8694 11999 8695 12025
rect 8695 11999 8721 12025
rect 8721 11999 8722 12025
rect 8694 11998 8722 11999
rect 7238 10934 7266 10962
rect 7350 10878 7378 10906
rect 7126 10542 7154 10570
rect 2142 10318 2170 10346
rect 4830 10262 4858 10290
rect 6062 10289 6090 10290
rect 6062 10263 6063 10289
rect 6063 10263 6089 10289
rect 6089 10263 6090 10289
rect 6062 10262 6090 10263
rect 6286 10038 6314 10066
rect 6790 10065 6818 10066
rect 6790 10039 6791 10065
rect 6791 10039 6817 10065
rect 6817 10039 6818 10065
rect 6790 10038 6818 10039
rect 7014 10038 7042 10066
rect 6566 9926 6594 9954
rect 2238 9813 2266 9814
rect 2238 9787 2239 9813
rect 2239 9787 2265 9813
rect 2265 9787 2266 9813
rect 2238 9786 2266 9787
rect 2290 9813 2318 9814
rect 2290 9787 2291 9813
rect 2291 9787 2317 9813
rect 2317 9787 2318 9813
rect 2290 9786 2318 9787
rect 2342 9813 2370 9814
rect 2342 9787 2343 9813
rect 2343 9787 2369 9813
rect 2369 9787 2370 9813
rect 2342 9786 2370 9787
rect 7350 10038 7378 10066
rect 2142 9225 2170 9226
rect 2142 9199 2143 9225
rect 2143 9199 2169 9225
rect 2169 9199 2170 9225
rect 2142 9198 2170 9199
rect 5446 9198 5474 9226
rect 966 9113 994 9114
rect 966 9087 967 9113
rect 967 9087 993 9113
rect 993 9087 994 9113
rect 966 9086 994 9087
rect 2238 9029 2266 9030
rect 2238 9003 2239 9029
rect 2239 9003 2265 9029
rect 2265 9003 2266 9029
rect 2238 9002 2266 9003
rect 2290 9029 2318 9030
rect 2290 9003 2291 9029
rect 2291 9003 2317 9029
rect 2317 9003 2318 9029
rect 2290 9002 2318 9003
rect 2342 9029 2370 9030
rect 2342 9003 2343 9029
rect 2343 9003 2369 9029
rect 2369 9003 2370 9029
rect 2342 9002 2370 9003
rect 966 8889 994 8890
rect 966 8863 967 8889
rect 967 8863 993 8889
rect 993 8863 994 8889
rect 966 8862 994 8863
rect 2142 8833 2170 8834
rect 2142 8807 2143 8833
rect 2143 8807 2169 8833
rect 2169 8807 2170 8833
rect 2142 8806 2170 8807
rect 6342 9086 6370 9114
rect 6846 8806 6874 8834
rect 7014 9198 7042 9226
rect 7294 9561 7322 9562
rect 7294 9535 7295 9561
rect 7295 9535 7321 9561
rect 7321 9535 7322 9561
rect 7294 9534 7322 9535
rect 7518 9534 7546 9562
rect 7910 11158 7938 11186
rect 7742 10905 7770 10906
rect 7742 10879 7743 10905
rect 7743 10879 7769 10905
rect 7769 10879 7770 10905
rect 7742 10878 7770 10879
rect 7686 10849 7714 10850
rect 7686 10823 7687 10849
rect 7687 10823 7713 10849
rect 7713 10823 7714 10849
rect 7686 10822 7714 10823
rect 7574 10598 7602 10626
rect 7742 10094 7770 10122
rect 9086 11942 9114 11970
rect 9030 11577 9058 11578
rect 9030 11551 9031 11577
rect 9031 11551 9057 11577
rect 9057 11551 9058 11577
rect 9030 11550 9058 11551
rect 7966 10206 7994 10234
rect 8246 10598 8274 10626
rect 8190 10542 8218 10570
rect 8134 10094 8162 10122
rect 7798 9590 7826 9618
rect 8134 9505 8162 9506
rect 8134 9479 8135 9505
rect 8135 9479 8161 9505
rect 8161 9479 8162 9505
rect 8134 9478 8162 9479
rect 7686 9337 7714 9338
rect 7686 9311 7687 9337
rect 7687 9311 7713 9337
rect 7713 9311 7714 9337
rect 7686 9310 7714 9311
rect 7798 9337 7826 9338
rect 7798 9311 7799 9337
rect 7799 9311 7825 9337
rect 7825 9311 7826 9337
rect 7798 9310 7826 9311
rect 7406 9254 7434 9282
rect 7070 9113 7098 9114
rect 7070 9087 7071 9113
rect 7071 9087 7097 9113
rect 7097 9087 7098 9113
rect 7070 9086 7098 9087
rect 7350 9169 7378 9170
rect 7350 9143 7351 9169
rect 7351 9143 7377 9169
rect 7377 9143 7378 9169
rect 7350 9142 7378 9143
rect 8302 10262 8330 10290
rect 9030 10990 9058 11018
rect 8750 10934 8778 10962
rect 8470 10038 8498 10066
rect 8638 10038 8666 10066
rect 9310 11998 9338 12026
rect 9590 12614 9618 12642
rect 9478 11886 9506 11914
rect 9198 11718 9226 11746
rect 9142 10934 9170 10962
rect 8974 10849 9002 10850
rect 8974 10823 8975 10849
rect 8975 10823 9001 10849
rect 9001 10823 9002 10849
rect 8974 10822 9002 10823
rect 8862 10345 8890 10346
rect 8862 10319 8863 10345
rect 8863 10319 8889 10345
rect 8889 10319 8890 10345
rect 8862 10318 8890 10319
rect 8750 10038 8778 10066
rect 8974 9982 9002 10010
rect 8806 9897 8834 9898
rect 8806 9871 8807 9897
rect 8807 9871 8833 9897
rect 8833 9871 8834 9897
rect 8806 9870 8834 9871
rect 8918 9814 8946 9842
rect 8638 9561 8666 9562
rect 8638 9535 8639 9561
rect 8639 9535 8665 9561
rect 8665 9535 8666 9561
rect 8638 9534 8666 9535
rect 8358 9169 8386 9170
rect 8358 9143 8359 9169
rect 8359 9143 8385 9169
rect 8385 9143 8386 9169
rect 8358 9142 8386 9143
rect 8694 9142 8722 9170
rect 8414 9113 8442 9114
rect 8414 9087 8415 9113
rect 8415 9087 8441 9113
rect 8441 9087 8442 9113
rect 8414 9086 8442 9087
rect 8190 8414 8218 8442
rect 8918 9534 8946 9562
rect 8974 9505 9002 9506
rect 8974 9479 8975 9505
rect 8975 9479 9001 9505
rect 9001 9479 9002 9505
rect 8974 9478 9002 9479
rect 8974 9198 9002 9226
rect 9142 10737 9170 10738
rect 9142 10711 9143 10737
rect 9143 10711 9169 10737
rect 9169 10711 9170 10737
rect 9142 10710 9170 10711
rect 9142 10598 9170 10626
rect 9254 10878 9282 10906
rect 9534 11998 9562 12026
rect 9646 12249 9674 12250
rect 9646 12223 9647 12249
rect 9647 12223 9673 12249
rect 9673 12223 9674 12249
rect 9646 12222 9674 12223
rect 9534 10822 9562 10850
rect 9590 10793 9618 10794
rect 9590 10767 9591 10793
rect 9591 10767 9617 10793
rect 9617 10767 9618 10793
rect 9590 10766 9618 10767
rect 9142 10289 9170 10290
rect 9142 10263 9143 10289
rect 9143 10263 9169 10289
rect 9169 10263 9170 10289
rect 9142 10262 9170 10263
rect 9198 10374 9226 10402
rect 9142 10038 9170 10066
rect 9870 12697 9898 12698
rect 9870 12671 9871 12697
rect 9871 12671 9897 12697
rect 9897 12671 9898 12697
rect 9870 12670 9898 12671
rect 10654 12753 10682 12754
rect 10654 12727 10655 12753
rect 10655 12727 10681 12753
rect 10681 12727 10682 12753
rect 10654 12726 10682 12727
rect 12110 13902 12138 13930
rect 11438 13230 11466 13258
rect 11382 13062 11410 13090
rect 10934 12865 10962 12866
rect 10934 12839 10935 12865
rect 10935 12839 10961 12865
rect 10961 12839 10962 12865
rect 10934 12838 10962 12839
rect 11438 12838 11466 12866
rect 10094 12670 10122 12698
rect 9918 12557 9946 12558
rect 9918 12531 9919 12557
rect 9919 12531 9945 12557
rect 9945 12531 9946 12557
rect 9918 12530 9946 12531
rect 9970 12557 9998 12558
rect 9970 12531 9971 12557
rect 9971 12531 9997 12557
rect 9997 12531 9998 12557
rect 9970 12530 9998 12531
rect 10022 12557 10050 12558
rect 10022 12531 10023 12557
rect 10023 12531 10049 12557
rect 10049 12531 10050 12557
rect 10022 12530 10050 12531
rect 9814 12249 9842 12250
rect 9814 12223 9815 12249
rect 9815 12223 9841 12249
rect 9841 12223 9842 12249
rect 9814 12222 9842 12223
rect 10150 12249 10178 12250
rect 10150 12223 10151 12249
rect 10151 12223 10177 12249
rect 10177 12223 10178 12249
rect 10150 12222 10178 12223
rect 9982 11998 10010 12026
rect 10094 11969 10122 11970
rect 10094 11943 10095 11969
rect 10095 11943 10121 11969
rect 10121 11943 10122 11969
rect 10094 11942 10122 11943
rect 9758 11718 9786 11746
rect 9814 11830 9842 11858
rect 10038 11886 10066 11914
rect 11158 12726 11186 12754
rect 10206 11886 10234 11914
rect 9702 11494 9730 11522
rect 10262 11857 10290 11858
rect 10262 11831 10263 11857
rect 10263 11831 10289 11857
rect 10289 11831 10290 11857
rect 10262 11830 10290 11831
rect 9918 11773 9946 11774
rect 9918 11747 9919 11773
rect 9919 11747 9945 11773
rect 9945 11747 9946 11773
rect 9918 11746 9946 11747
rect 9970 11773 9998 11774
rect 9970 11747 9971 11773
rect 9971 11747 9997 11773
rect 9997 11747 9998 11773
rect 9970 11746 9998 11747
rect 10022 11773 10050 11774
rect 10022 11747 10023 11773
rect 10023 11747 10049 11773
rect 10049 11747 10050 11773
rect 10022 11746 10050 11747
rect 10094 11774 10122 11802
rect 9926 11521 9954 11522
rect 9926 11495 9927 11521
rect 9927 11495 9953 11521
rect 9953 11495 9954 11521
rect 9926 11494 9954 11495
rect 11102 11886 11130 11914
rect 10822 11857 10850 11858
rect 10822 11831 10823 11857
rect 10823 11831 10849 11857
rect 10849 11831 10850 11857
rect 10822 11830 10850 11831
rect 10710 11774 10738 11802
rect 10654 11577 10682 11578
rect 10654 11551 10655 11577
rect 10655 11551 10681 11577
rect 10681 11551 10682 11577
rect 10654 11550 10682 11551
rect 10374 11494 10402 11522
rect 10878 11521 10906 11522
rect 10878 11495 10879 11521
rect 10879 11495 10905 11521
rect 10905 11495 10906 11521
rect 10878 11494 10906 11495
rect 10206 11465 10234 11466
rect 10206 11439 10207 11465
rect 10207 11439 10233 11465
rect 10233 11439 10234 11465
rect 10206 11438 10234 11439
rect 10878 11102 10906 11130
rect 9918 10989 9946 10990
rect 9918 10963 9919 10989
rect 9919 10963 9945 10989
rect 9945 10963 9946 10989
rect 9918 10962 9946 10963
rect 9970 10989 9998 10990
rect 9970 10963 9971 10989
rect 9971 10963 9997 10989
rect 9997 10963 9998 10989
rect 9970 10962 9998 10963
rect 10022 10989 10050 10990
rect 10022 10963 10023 10989
rect 10023 10963 10049 10989
rect 10049 10963 10050 10989
rect 10022 10962 10050 10963
rect 9758 10878 9786 10906
rect 10150 10878 10178 10906
rect 9702 10710 9730 10738
rect 9366 10206 9394 10234
rect 9310 10038 9338 10066
rect 9366 9953 9394 9954
rect 9366 9927 9367 9953
rect 9367 9927 9393 9953
rect 9393 9927 9394 9953
rect 9366 9926 9394 9927
rect 9310 9702 9338 9730
rect 9310 9590 9338 9618
rect 9030 9086 9058 9114
rect 9366 9646 9394 9674
rect 9366 9310 9394 9338
rect 10094 10318 10122 10346
rect 9918 10205 9946 10206
rect 9918 10179 9919 10205
rect 9919 10179 9945 10205
rect 9945 10179 9946 10205
rect 9918 10178 9946 10179
rect 9970 10205 9998 10206
rect 9970 10179 9971 10205
rect 9971 10179 9997 10205
rect 9997 10179 9998 10205
rect 9970 10178 9998 10179
rect 10022 10205 10050 10206
rect 10022 10179 10023 10205
rect 10023 10179 10049 10205
rect 10049 10179 10050 10205
rect 10022 10178 10050 10179
rect 10094 9982 10122 10010
rect 10710 10766 10738 10794
rect 10318 10542 10346 10570
rect 10934 10598 10962 10626
rect 10878 10542 10906 10570
rect 10318 10401 10346 10402
rect 10318 10375 10319 10401
rect 10319 10375 10345 10401
rect 10345 10375 10346 10401
rect 10318 10374 10346 10375
rect 9982 9926 10010 9954
rect 10934 9870 10962 9898
rect 10262 9646 10290 9674
rect 9982 9617 10010 9618
rect 9982 9591 9983 9617
rect 9983 9591 10009 9617
rect 10009 9591 10010 9617
rect 9982 9590 10010 9591
rect 10598 9617 10626 9618
rect 10598 9591 10599 9617
rect 10599 9591 10625 9617
rect 10625 9591 10626 9617
rect 10598 9590 10626 9591
rect 9758 9534 9786 9562
rect 10766 9534 10794 9562
rect 9646 9310 9674 9338
rect 8694 8358 8722 8386
rect 2238 8245 2266 8246
rect 2238 8219 2239 8245
rect 2239 8219 2265 8245
rect 2265 8219 2266 8245
rect 2238 8218 2266 8219
rect 2290 8245 2318 8246
rect 2290 8219 2291 8245
rect 2291 8219 2317 8245
rect 2317 8219 2318 8245
rect 2290 8218 2318 8219
rect 2342 8245 2370 8246
rect 2342 8219 2343 8245
rect 2343 8219 2369 8245
rect 2369 8219 2370 8245
rect 2342 8218 2370 8219
rect 2238 7461 2266 7462
rect 2238 7435 2239 7461
rect 2239 7435 2265 7461
rect 2265 7435 2266 7461
rect 2238 7434 2266 7435
rect 2290 7461 2318 7462
rect 2290 7435 2291 7461
rect 2291 7435 2317 7461
rect 2317 7435 2318 7461
rect 2290 7434 2318 7435
rect 2342 7461 2370 7462
rect 2342 7435 2343 7461
rect 2343 7435 2369 7461
rect 2369 7435 2370 7461
rect 2342 7434 2370 7435
rect 8358 7265 8386 7266
rect 8358 7239 8359 7265
rect 8359 7239 8385 7265
rect 8385 7239 8386 7265
rect 8358 7238 8386 7239
rect 9478 8470 9506 8498
rect 9254 8441 9282 8442
rect 9254 8415 9255 8441
rect 9255 8415 9281 8441
rect 9281 8415 9282 8441
rect 9254 8414 9282 8415
rect 9918 9421 9946 9422
rect 9918 9395 9919 9421
rect 9919 9395 9945 9421
rect 9945 9395 9946 9421
rect 9918 9394 9946 9395
rect 9970 9421 9998 9422
rect 9970 9395 9971 9421
rect 9971 9395 9997 9421
rect 9997 9395 9998 9421
rect 9970 9394 9998 9395
rect 10022 9421 10050 9422
rect 10022 9395 10023 9421
rect 10023 9395 10049 9421
rect 10049 9395 10050 9421
rect 10022 9394 10050 9395
rect 10206 9478 10234 9506
rect 9926 9225 9954 9226
rect 9926 9199 9927 9225
rect 9927 9199 9953 9225
rect 9953 9199 9954 9225
rect 9926 9198 9954 9199
rect 10766 9254 10794 9282
rect 10038 9142 10066 9170
rect 10878 9646 10906 9674
rect 11886 13230 11914 13258
rect 12222 13145 12250 13146
rect 12222 13119 12223 13145
rect 12223 13119 12249 13145
rect 12249 13119 12250 13145
rect 12222 13118 12250 13119
rect 11998 13089 12026 13090
rect 11998 13063 11999 13089
rect 11999 13063 12025 13089
rect 12025 13063 12026 13089
rect 11998 13062 12026 13063
rect 12390 13062 12418 13090
rect 11382 12614 11410 12642
rect 11550 12670 11578 12698
rect 11830 12670 11858 12698
rect 11550 12278 11578 12306
rect 11662 12417 11690 12418
rect 11662 12391 11663 12417
rect 11663 12391 11689 12417
rect 11689 12391 11690 12417
rect 11662 12390 11690 12391
rect 11270 11830 11298 11858
rect 11214 11606 11242 11634
rect 11438 11774 11466 11802
rect 11326 11521 11354 11522
rect 11326 11495 11327 11521
rect 11327 11495 11353 11521
rect 11353 11495 11354 11521
rect 11326 11494 11354 11495
rect 11382 11270 11410 11298
rect 11214 10542 11242 10570
rect 11326 10737 11354 10738
rect 11326 10711 11327 10737
rect 11327 10711 11353 10737
rect 11353 10711 11354 10737
rect 11326 10710 11354 10711
rect 11102 10457 11130 10458
rect 11102 10431 11103 10457
rect 11103 10431 11129 10457
rect 11129 10431 11130 10457
rect 11102 10430 11130 10431
rect 11046 9814 11074 9842
rect 11102 10318 11130 10346
rect 10990 9478 11018 9506
rect 11046 9590 11074 9618
rect 11046 9310 11074 9338
rect 11158 10289 11186 10290
rect 11158 10263 11159 10289
rect 11159 10263 11185 10289
rect 11185 10263 11186 10289
rect 11158 10262 11186 10263
rect 12110 12417 12138 12418
rect 12110 12391 12111 12417
rect 12111 12391 12137 12417
rect 12137 12391 12138 12417
rect 12110 12390 12138 12391
rect 11662 11830 11690 11858
rect 11886 12334 11914 12362
rect 11606 11550 11634 11578
rect 11662 11606 11690 11634
rect 12222 12361 12250 12362
rect 12222 12335 12223 12361
rect 12223 12335 12249 12361
rect 12249 12335 12250 12361
rect 12222 12334 12250 12335
rect 11942 11886 11970 11914
rect 11718 11521 11746 11522
rect 11718 11495 11719 11521
rect 11719 11495 11745 11521
rect 11745 11495 11746 11521
rect 11718 11494 11746 11495
rect 11438 11129 11466 11130
rect 11438 11103 11439 11129
rect 11439 11103 11465 11129
rect 11465 11103 11466 11129
rect 11438 11102 11466 11103
rect 11438 10542 11466 10570
rect 11326 9953 11354 9954
rect 11326 9927 11327 9953
rect 11327 9927 11353 9953
rect 11353 9927 11354 9953
rect 11326 9926 11354 9927
rect 11270 9702 11298 9730
rect 11326 9561 11354 9562
rect 11326 9535 11327 9561
rect 11327 9535 11353 9561
rect 11353 9535 11354 9561
rect 11326 9534 11354 9535
rect 11382 9505 11410 9506
rect 11382 9479 11383 9505
rect 11383 9479 11409 9505
rect 11409 9479 11410 9505
rect 11382 9478 11410 9479
rect 11158 9310 11186 9338
rect 11382 9337 11410 9338
rect 11382 9311 11383 9337
rect 11383 9311 11409 9337
rect 11409 9311 11410 9337
rect 11382 9310 11410 9311
rect 11606 10150 11634 10178
rect 11774 11270 11802 11298
rect 11774 10094 11802 10122
rect 11494 9310 11522 9338
rect 10822 8918 10850 8946
rect 10934 9086 10962 9114
rect 11102 9198 11130 9226
rect 11214 9225 11242 9226
rect 11214 9199 11215 9225
rect 11215 9199 11241 9225
rect 11241 9199 11242 9225
rect 11214 9198 11242 9199
rect 11606 9198 11634 9226
rect 11662 9926 11690 9954
rect 11158 8945 11186 8946
rect 11158 8919 11159 8945
rect 11159 8919 11185 8945
rect 11185 8919 11186 8945
rect 11158 8918 11186 8919
rect 9918 8637 9946 8638
rect 9918 8611 9919 8637
rect 9919 8611 9945 8637
rect 9945 8611 9946 8637
rect 9918 8610 9946 8611
rect 9970 8637 9998 8638
rect 9970 8611 9971 8637
rect 9971 8611 9997 8637
rect 9997 8611 9998 8637
rect 9970 8610 9998 8611
rect 10022 8637 10050 8638
rect 10022 8611 10023 8637
rect 10023 8611 10049 8637
rect 10049 8611 10050 8637
rect 10022 8610 10050 8611
rect 9590 8385 9618 8386
rect 9590 8359 9591 8385
rect 9591 8359 9617 8385
rect 9617 8359 9618 8385
rect 9590 8358 9618 8359
rect 9702 8358 9730 8386
rect 9982 8497 10010 8498
rect 9982 8471 9983 8497
rect 9983 8471 10009 8497
rect 10009 8471 10010 8497
rect 9982 8470 10010 8471
rect 10486 8385 10514 8386
rect 10486 8359 10487 8385
rect 10487 8359 10513 8385
rect 10513 8359 10514 8385
rect 10486 8358 10514 8359
rect 9982 8302 10010 8330
rect 9918 7853 9946 7854
rect 9918 7827 9919 7853
rect 9919 7827 9945 7853
rect 9945 7827 9946 7853
rect 9918 7826 9946 7827
rect 9970 7853 9998 7854
rect 9970 7827 9971 7853
rect 9971 7827 9997 7853
rect 9997 7827 9998 7853
rect 9970 7826 9998 7827
rect 10022 7853 10050 7854
rect 10022 7827 10023 7853
rect 10023 7827 10049 7853
rect 10049 7827 10050 7853
rect 10022 7826 10050 7827
rect 9702 7630 9730 7658
rect 10710 8358 10738 8386
rect 10598 7630 10626 7658
rect 13230 14182 13258 14210
rect 12838 13566 12866 13594
rect 17598 18437 17626 18438
rect 17598 18411 17599 18437
rect 17599 18411 17625 18437
rect 17625 18411 17626 18437
rect 17598 18410 17626 18411
rect 17650 18437 17678 18438
rect 17650 18411 17651 18437
rect 17651 18411 17677 18437
rect 17677 18411 17678 18437
rect 17650 18410 17678 18411
rect 17702 18437 17730 18438
rect 17702 18411 17703 18437
rect 17703 18411 17729 18437
rect 17729 18411 17730 18437
rect 17702 18410 17730 18411
rect 17598 17653 17626 17654
rect 17598 17627 17599 17653
rect 17599 17627 17625 17653
rect 17625 17627 17626 17653
rect 17598 17626 17626 17627
rect 17650 17653 17678 17654
rect 17650 17627 17651 17653
rect 17651 17627 17677 17653
rect 17677 17627 17678 17653
rect 17650 17626 17678 17627
rect 17702 17653 17730 17654
rect 17702 17627 17703 17653
rect 17703 17627 17729 17653
rect 17729 17627 17730 17653
rect 17702 17626 17730 17627
rect 17598 16869 17626 16870
rect 17598 16843 17599 16869
rect 17599 16843 17625 16869
rect 17625 16843 17626 16869
rect 17598 16842 17626 16843
rect 17650 16869 17678 16870
rect 17650 16843 17651 16869
rect 17651 16843 17677 16869
rect 17677 16843 17678 16869
rect 17650 16842 17678 16843
rect 17702 16869 17730 16870
rect 17702 16843 17703 16869
rect 17703 16843 17729 16869
rect 17729 16843 17730 16869
rect 17702 16842 17730 16843
rect 17598 16085 17626 16086
rect 17598 16059 17599 16085
rect 17599 16059 17625 16085
rect 17625 16059 17626 16085
rect 17598 16058 17626 16059
rect 17650 16085 17678 16086
rect 17650 16059 17651 16085
rect 17651 16059 17677 16085
rect 17677 16059 17678 16085
rect 17650 16058 17678 16059
rect 17702 16085 17730 16086
rect 17702 16059 17703 16085
rect 17703 16059 17729 16085
rect 17729 16059 17730 16085
rect 17702 16058 17730 16059
rect 17598 15301 17626 15302
rect 17598 15275 17599 15301
rect 17599 15275 17625 15301
rect 17625 15275 17626 15301
rect 17598 15274 17626 15275
rect 17650 15301 17678 15302
rect 17650 15275 17651 15301
rect 17651 15275 17677 15301
rect 17677 15275 17678 15301
rect 17650 15274 17678 15275
rect 17702 15301 17730 15302
rect 17702 15275 17703 15301
rect 17703 15275 17729 15301
rect 17729 15275 17730 15301
rect 17702 15274 17730 15275
rect 17598 14517 17626 14518
rect 17598 14491 17599 14517
rect 17599 14491 17625 14517
rect 17625 14491 17626 14517
rect 17598 14490 17626 14491
rect 17650 14517 17678 14518
rect 17650 14491 17651 14517
rect 17651 14491 17677 14517
rect 17677 14491 17678 14517
rect 17650 14490 17678 14491
rect 17702 14517 17730 14518
rect 17702 14491 17703 14517
rect 17703 14491 17729 14517
rect 17729 14491 17730 14517
rect 17702 14490 17730 14491
rect 14294 14182 14322 14210
rect 17598 13733 17626 13734
rect 17598 13707 17599 13733
rect 17599 13707 17625 13733
rect 17625 13707 17626 13733
rect 17598 13706 17626 13707
rect 17650 13733 17678 13734
rect 17650 13707 17651 13733
rect 17651 13707 17677 13733
rect 17677 13707 17678 13733
rect 17650 13706 17678 13707
rect 17702 13733 17730 13734
rect 17702 13707 17703 13733
rect 17703 13707 17729 13733
rect 17729 13707 17730 13733
rect 17702 13706 17730 13707
rect 13230 13593 13258 13594
rect 13230 13567 13231 13593
rect 13231 13567 13257 13593
rect 13257 13567 13258 13593
rect 13230 13566 13258 13567
rect 12782 13145 12810 13146
rect 12782 13119 12783 13145
rect 12783 13119 12809 13145
rect 12809 13119 12810 13145
rect 12782 13118 12810 13119
rect 17598 12949 17626 12950
rect 17598 12923 17599 12949
rect 17599 12923 17625 12949
rect 17625 12923 17626 12949
rect 17598 12922 17626 12923
rect 17650 12949 17678 12950
rect 17650 12923 17651 12949
rect 17651 12923 17677 12949
rect 17677 12923 17678 12949
rect 17650 12922 17678 12923
rect 17702 12949 17730 12950
rect 17702 12923 17703 12949
rect 17703 12923 17729 12949
rect 17729 12923 17730 12949
rect 17702 12922 17730 12923
rect 12726 12670 12754 12698
rect 12614 11998 12642 12026
rect 12446 10430 12474 10458
rect 12054 10094 12082 10122
rect 11886 9646 11914 9674
rect 11942 9534 11970 9562
rect 11718 9422 11746 9450
rect 11998 9478 12026 9506
rect 11998 9310 12026 9338
rect 11662 8470 11690 8498
rect 11326 8302 11354 8330
rect 11886 8414 11914 8442
rect 11942 8582 11970 8610
rect 11830 8358 11858 8386
rect 11774 7742 11802 7770
rect 12054 9366 12082 9394
rect 12278 10094 12306 10122
rect 12390 10065 12418 10066
rect 12390 10039 12391 10065
rect 12391 10039 12417 10065
rect 12417 10039 12418 10065
rect 12390 10038 12418 10039
rect 12222 9478 12250 9506
rect 12558 10150 12586 10178
rect 12446 9422 12474 9450
rect 12502 9982 12530 10010
rect 12670 11774 12698 11802
rect 12950 12670 12978 12698
rect 13902 12697 13930 12698
rect 13902 12671 13903 12697
rect 13903 12671 13929 12697
rect 13929 12671 13930 12697
rect 13902 12670 13930 12671
rect 13006 12641 13034 12642
rect 13006 12615 13007 12641
rect 13007 12615 13033 12641
rect 13033 12615 13034 12641
rect 13006 12614 13034 12615
rect 13118 12502 13146 12530
rect 12782 12390 12810 12418
rect 13006 12361 13034 12362
rect 13006 12335 13007 12361
rect 13007 12335 13033 12361
rect 13033 12335 13034 12361
rect 13006 12334 13034 12335
rect 13230 12361 13258 12362
rect 13230 12335 13231 12361
rect 13231 12335 13257 12361
rect 13257 12335 13258 12361
rect 13230 12334 13258 12335
rect 14742 12697 14770 12698
rect 14742 12671 14743 12697
rect 14743 12671 14769 12697
rect 14769 12671 14770 12697
rect 14742 12670 14770 12671
rect 19950 12782 19978 12810
rect 18830 12753 18858 12754
rect 18830 12727 18831 12753
rect 18831 12727 18857 12753
rect 18857 12727 18858 12753
rect 18830 12726 18858 12727
rect 18718 12670 18746 12698
rect 14630 12614 14658 12642
rect 14854 12614 14882 12642
rect 12782 11830 12810 11858
rect 13006 11774 13034 11802
rect 13062 11830 13090 11858
rect 12894 11521 12922 11522
rect 12894 11495 12895 11521
rect 12895 11495 12921 11521
rect 12921 11495 12922 11521
rect 12894 11494 12922 11495
rect 12950 11438 12978 11466
rect 12838 10038 12866 10066
rect 12670 9926 12698 9954
rect 12614 9897 12642 9898
rect 12614 9871 12615 9897
rect 12615 9871 12641 9897
rect 12641 9871 12642 9897
rect 12614 9870 12642 9871
rect 12614 9673 12642 9674
rect 12614 9647 12615 9673
rect 12615 9647 12641 9673
rect 12641 9647 12642 9673
rect 12614 9646 12642 9647
rect 12502 9310 12530 9338
rect 12222 9142 12250 9170
rect 12166 9086 12194 9114
rect 12670 9590 12698 9618
rect 13006 11550 13034 11578
rect 12838 9953 12866 9954
rect 12838 9927 12839 9953
rect 12839 9927 12865 9953
rect 12865 9927 12866 9953
rect 12838 9926 12866 9927
rect 13062 10654 13090 10682
rect 12950 10009 12978 10010
rect 12950 9983 12951 10009
rect 12951 9983 12977 10009
rect 12977 9983 12978 10009
rect 12950 9982 12978 9983
rect 13006 9953 13034 9954
rect 13006 9927 13007 9953
rect 13007 9927 13033 9953
rect 13033 9927 13034 9953
rect 13006 9926 13034 9927
rect 12950 9422 12978 9450
rect 13846 12334 13874 12362
rect 20006 12446 20034 12474
rect 17598 12165 17626 12166
rect 17598 12139 17599 12165
rect 17599 12139 17625 12165
rect 17625 12139 17626 12165
rect 17598 12138 17626 12139
rect 17650 12165 17678 12166
rect 17650 12139 17651 12165
rect 17651 12139 17677 12165
rect 17677 12139 17678 12165
rect 17650 12138 17678 12139
rect 17702 12165 17730 12166
rect 17702 12139 17703 12165
rect 17703 12139 17729 12165
rect 17729 12139 17730 12165
rect 17702 12138 17730 12139
rect 13902 11942 13930 11970
rect 14742 11942 14770 11970
rect 14014 11857 14042 11858
rect 14014 11831 14015 11857
rect 14015 11831 14041 11857
rect 14041 11831 14042 11857
rect 14014 11830 14042 11831
rect 13286 11774 13314 11802
rect 13678 11521 13706 11522
rect 13678 11495 13679 11521
rect 13679 11495 13705 11521
rect 13705 11495 13706 11521
rect 13678 11494 13706 11495
rect 18830 11969 18858 11970
rect 18830 11943 18831 11969
rect 18831 11943 18857 11969
rect 18857 11943 18858 11969
rect 18830 11942 18858 11943
rect 20006 11774 20034 11802
rect 17598 11381 17626 11382
rect 17598 11355 17599 11381
rect 17599 11355 17625 11381
rect 17625 11355 17626 11381
rect 17598 11354 17626 11355
rect 17650 11381 17678 11382
rect 17650 11355 17651 11381
rect 17651 11355 17677 11381
rect 17677 11355 17678 11381
rect 17650 11354 17678 11355
rect 17702 11381 17730 11382
rect 17702 11355 17703 11381
rect 17703 11355 17729 11381
rect 17729 11355 17730 11381
rect 17702 11354 17730 11355
rect 14518 10681 14546 10682
rect 14518 10655 14519 10681
rect 14519 10655 14545 10681
rect 14545 10655 14546 10681
rect 14518 10654 14546 10655
rect 13174 10038 13202 10066
rect 17598 10597 17626 10598
rect 17598 10571 17599 10597
rect 17599 10571 17625 10597
rect 17625 10571 17626 10597
rect 17598 10570 17626 10571
rect 17650 10597 17678 10598
rect 17650 10571 17651 10597
rect 17651 10571 17677 10597
rect 17677 10571 17678 10597
rect 17650 10570 17678 10571
rect 17702 10597 17730 10598
rect 17702 10571 17703 10597
rect 17703 10571 17729 10597
rect 17729 10571 17730 10597
rect 17702 10570 17730 10571
rect 14910 10094 14938 10122
rect 20006 10430 20034 10458
rect 18830 10094 18858 10122
rect 20118 10094 20146 10122
rect 13286 9673 13314 9674
rect 13286 9647 13287 9673
rect 13287 9647 13313 9673
rect 13313 9647 13314 9673
rect 13286 9646 13314 9647
rect 13006 9366 13034 9394
rect 13846 9953 13874 9954
rect 13846 9927 13847 9953
rect 13847 9927 13873 9953
rect 13873 9927 13874 9953
rect 13846 9926 13874 9927
rect 17598 9813 17626 9814
rect 17598 9787 17599 9813
rect 17599 9787 17625 9813
rect 17625 9787 17626 9813
rect 17598 9786 17626 9787
rect 17650 9813 17678 9814
rect 17650 9787 17651 9813
rect 17651 9787 17677 9813
rect 17677 9787 17678 9813
rect 17650 9786 17678 9787
rect 17702 9813 17730 9814
rect 17702 9787 17703 9813
rect 17703 9787 17729 9813
rect 17729 9787 17730 9813
rect 17702 9786 17730 9787
rect 14294 9561 14322 9562
rect 14294 9535 14295 9561
rect 14295 9535 14321 9561
rect 14321 9535 14322 9561
rect 14294 9534 14322 9535
rect 14798 9534 14826 9562
rect 13398 9366 13426 9394
rect 13510 9254 13538 9282
rect 12614 9113 12642 9114
rect 12614 9087 12615 9113
rect 12615 9087 12641 9113
rect 12641 9087 12642 9113
rect 12614 9086 12642 9087
rect 12670 8889 12698 8890
rect 12670 8863 12671 8889
rect 12671 8863 12697 8889
rect 12697 8863 12698 8889
rect 12670 8862 12698 8863
rect 12838 8833 12866 8834
rect 12838 8807 12839 8833
rect 12839 8807 12865 8833
rect 12865 8807 12866 8833
rect 12838 8806 12866 8807
rect 12614 8777 12642 8778
rect 12614 8751 12615 8777
rect 12615 8751 12641 8777
rect 12641 8751 12642 8777
rect 12614 8750 12642 8751
rect 12390 8721 12418 8722
rect 12390 8695 12391 8721
rect 12391 8695 12417 8721
rect 12417 8695 12418 8721
rect 12390 8694 12418 8695
rect 12334 8582 12362 8610
rect 12838 8582 12866 8610
rect 13230 8889 13258 8890
rect 13230 8863 13231 8889
rect 13231 8863 13257 8889
rect 13257 8863 13258 8889
rect 13230 8862 13258 8863
rect 20006 9758 20034 9786
rect 18830 9534 18858 9562
rect 17598 9029 17626 9030
rect 17598 9003 17599 9029
rect 17599 9003 17625 9029
rect 17625 9003 17626 9029
rect 17598 9002 17626 9003
rect 17650 9029 17678 9030
rect 17650 9003 17651 9029
rect 17651 9003 17677 9029
rect 17677 9003 17678 9029
rect 17650 9002 17678 9003
rect 17702 9029 17730 9030
rect 17702 9003 17703 9029
rect 17703 9003 17729 9029
rect 17729 9003 17730 9029
rect 17702 9002 17730 9003
rect 13958 8862 13986 8890
rect 13398 8806 13426 8834
rect 12894 8694 12922 8722
rect 12334 8358 12362 8386
rect 12670 8385 12698 8386
rect 12670 8359 12671 8385
rect 12671 8359 12697 8385
rect 12697 8359 12698 8385
rect 12670 8358 12698 8359
rect 12614 8302 12642 8330
rect 10934 7630 10962 7658
rect 10878 7574 10906 7602
rect 8750 7238 8778 7266
rect 2238 6677 2266 6678
rect 2238 6651 2239 6677
rect 2239 6651 2265 6677
rect 2265 6651 2266 6677
rect 2238 6650 2266 6651
rect 2290 6677 2318 6678
rect 2290 6651 2291 6677
rect 2291 6651 2317 6677
rect 2317 6651 2318 6677
rect 2290 6650 2318 6651
rect 2342 6677 2370 6678
rect 2342 6651 2343 6677
rect 2343 6651 2369 6677
rect 2369 6651 2370 6677
rect 2342 6650 2370 6651
rect 2238 5893 2266 5894
rect 2238 5867 2239 5893
rect 2239 5867 2265 5893
rect 2265 5867 2266 5893
rect 2238 5866 2266 5867
rect 2290 5893 2318 5894
rect 2290 5867 2291 5893
rect 2291 5867 2317 5893
rect 2317 5867 2318 5893
rect 2290 5866 2318 5867
rect 2342 5893 2370 5894
rect 2342 5867 2343 5893
rect 2343 5867 2369 5893
rect 2369 5867 2370 5893
rect 2342 5866 2370 5867
rect 2238 5109 2266 5110
rect 2238 5083 2239 5109
rect 2239 5083 2265 5109
rect 2265 5083 2266 5109
rect 2238 5082 2266 5083
rect 2290 5109 2318 5110
rect 2290 5083 2291 5109
rect 2291 5083 2317 5109
rect 2317 5083 2318 5109
rect 2290 5082 2318 5083
rect 2342 5109 2370 5110
rect 2342 5083 2343 5109
rect 2343 5083 2369 5109
rect 2369 5083 2370 5109
rect 2342 5082 2370 5083
rect 2238 4325 2266 4326
rect 2238 4299 2239 4325
rect 2239 4299 2265 4325
rect 2265 4299 2266 4325
rect 2238 4298 2266 4299
rect 2290 4325 2318 4326
rect 2290 4299 2291 4325
rect 2291 4299 2317 4325
rect 2317 4299 2318 4325
rect 2290 4298 2318 4299
rect 2342 4325 2370 4326
rect 2342 4299 2343 4325
rect 2343 4299 2369 4325
rect 2369 4299 2370 4325
rect 2342 4298 2370 4299
rect 9982 7265 10010 7266
rect 9982 7239 9983 7265
rect 9983 7239 10009 7265
rect 10009 7239 10010 7265
rect 9982 7238 10010 7239
rect 9918 7069 9946 7070
rect 9918 7043 9919 7069
rect 9919 7043 9945 7069
rect 9945 7043 9946 7069
rect 9918 7042 9946 7043
rect 9970 7069 9998 7070
rect 9970 7043 9971 7069
rect 9971 7043 9997 7069
rect 9997 7043 9998 7069
rect 9970 7042 9998 7043
rect 10022 7069 10050 7070
rect 10022 7043 10023 7069
rect 10023 7043 10049 7069
rect 10049 7043 10050 7069
rect 10022 7042 10050 7043
rect 9870 6873 9898 6874
rect 9870 6847 9871 6873
rect 9871 6847 9897 6873
rect 9897 6847 9898 6873
rect 9870 6846 9898 6847
rect 9918 6285 9946 6286
rect 9918 6259 9919 6285
rect 9919 6259 9945 6285
rect 9945 6259 9946 6285
rect 9918 6258 9946 6259
rect 9970 6285 9998 6286
rect 9970 6259 9971 6285
rect 9971 6259 9997 6285
rect 9997 6259 9998 6285
rect 9970 6258 9998 6259
rect 10022 6285 10050 6286
rect 10022 6259 10023 6285
rect 10023 6259 10049 6285
rect 10049 6259 10050 6285
rect 10022 6258 10050 6259
rect 9918 5501 9946 5502
rect 9918 5475 9919 5501
rect 9919 5475 9945 5501
rect 9945 5475 9946 5501
rect 9918 5474 9946 5475
rect 9970 5501 9998 5502
rect 9970 5475 9971 5501
rect 9971 5475 9997 5501
rect 9997 5475 9998 5501
rect 9970 5474 9998 5475
rect 10022 5501 10050 5502
rect 10022 5475 10023 5501
rect 10023 5475 10049 5501
rect 10049 5475 10050 5501
rect 10022 5474 10050 5475
rect 9918 4717 9946 4718
rect 9918 4691 9919 4717
rect 9919 4691 9945 4717
rect 9945 4691 9946 4717
rect 9918 4690 9946 4691
rect 9970 4717 9998 4718
rect 9970 4691 9971 4717
rect 9971 4691 9997 4717
rect 9997 4691 9998 4717
rect 9970 4690 9998 4691
rect 10022 4717 10050 4718
rect 10022 4691 10023 4717
rect 10023 4691 10049 4717
rect 10049 4691 10050 4717
rect 10022 4690 10050 4691
rect 2238 3541 2266 3542
rect 2238 3515 2239 3541
rect 2239 3515 2265 3541
rect 2265 3515 2266 3541
rect 2238 3514 2266 3515
rect 2290 3541 2318 3542
rect 2290 3515 2291 3541
rect 2291 3515 2317 3541
rect 2317 3515 2318 3541
rect 2290 3514 2318 3515
rect 2342 3541 2370 3542
rect 2342 3515 2343 3541
rect 2343 3515 2369 3541
rect 2369 3515 2370 3541
rect 2342 3514 2370 3515
rect 2238 2757 2266 2758
rect 2238 2731 2239 2757
rect 2239 2731 2265 2757
rect 2265 2731 2266 2757
rect 2238 2730 2266 2731
rect 2290 2757 2318 2758
rect 2290 2731 2291 2757
rect 2291 2731 2317 2757
rect 2317 2731 2318 2757
rect 2290 2730 2318 2731
rect 2342 2757 2370 2758
rect 2342 2731 2343 2757
rect 2343 2731 2369 2757
rect 2369 2731 2370 2757
rect 2342 2730 2370 2731
rect 9918 3933 9946 3934
rect 9918 3907 9919 3933
rect 9919 3907 9945 3933
rect 9945 3907 9946 3933
rect 9918 3906 9946 3907
rect 9970 3933 9998 3934
rect 9970 3907 9971 3933
rect 9971 3907 9997 3933
rect 9997 3907 9998 3933
rect 9970 3906 9998 3907
rect 10022 3933 10050 3934
rect 10022 3907 10023 3933
rect 10023 3907 10049 3933
rect 10049 3907 10050 3933
rect 10022 3906 10050 3907
rect 9918 3149 9946 3150
rect 9918 3123 9919 3149
rect 9919 3123 9945 3149
rect 9945 3123 9946 3149
rect 9918 3122 9946 3123
rect 9970 3149 9998 3150
rect 9970 3123 9971 3149
rect 9971 3123 9997 3149
rect 9997 3123 9998 3149
rect 9970 3122 9998 3123
rect 10022 3149 10050 3150
rect 10022 3123 10023 3149
rect 10023 3123 10049 3149
rect 10049 3123 10050 3149
rect 10022 3122 10050 3123
rect 9918 2365 9946 2366
rect 9918 2339 9919 2365
rect 9919 2339 9945 2365
rect 9945 2339 9946 2365
rect 9918 2338 9946 2339
rect 9970 2365 9998 2366
rect 9970 2339 9971 2365
rect 9971 2339 9997 2365
rect 9997 2339 9998 2365
rect 9970 2338 9998 2339
rect 10022 2365 10050 2366
rect 10022 2339 10023 2365
rect 10023 2339 10049 2365
rect 10049 2339 10050 2365
rect 10022 2338 10050 2339
rect 11382 7601 11410 7602
rect 11382 7575 11383 7601
rect 11383 7575 11409 7601
rect 11409 7575 11410 7601
rect 11382 7574 11410 7575
rect 11158 6846 11186 6874
rect 11270 6734 11298 6762
rect 12950 8470 12978 8498
rect 12838 7769 12866 7770
rect 12838 7743 12839 7769
rect 12839 7743 12865 7769
rect 12865 7743 12866 7769
rect 12838 7742 12866 7743
rect 12222 7574 12250 7602
rect 12670 7601 12698 7602
rect 12670 7575 12671 7601
rect 12671 7575 12697 7601
rect 12697 7575 12698 7601
rect 12670 7574 12698 7575
rect 13118 7601 13146 7602
rect 13118 7575 13119 7601
rect 13119 7575 13145 7601
rect 13145 7575 13146 7601
rect 13118 7574 13146 7575
rect 13398 7574 13426 7602
rect 13902 8750 13930 8778
rect 14294 8889 14322 8890
rect 14294 8863 14295 8889
rect 14295 8863 14321 8889
rect 14321 8863 14322 8889
rect 14294 8862 14322 8863
rect 14630 8833 14658 8834
rect 14630 8807 14631 8833
rect 14631 8807 14657 8833
rect 14657 8807 14658 8833
rect 14630 8806 14658 8807
rect 18830 8833 18858 8834
rect 18830 8807 18831 8833
rect 18831 8807 18857 8833
rect 18857 8807 18858 8833
rect 18830 8806 18858 8807
rect 20006 8750 20034 8778
rect 17598 8245 17626 8246
rect 17598 8219 17599 8245
rect 17599 8219 17625 8245
rect 17625 8219 17626 8245
rect 17598 8218 17626 8219
rect 17650 8245 17678 8246
rect 17650 8219 17651 8245
rect 17651 8219 17677 8245
rect 17677 8219 17678 8245
rect 17650 8218 17678 8219
rect 17702 8245 17730 8246
rect 17702 8219 17703 8245
rect 17703 8219 17729 8245
rect 17729 8219 17730 8245
rect 17702 8218 17730 8219
rect 11494 6873 11522 6874
rect 11494 6847 11495 6873
rect 11495 6847 11521 6873
rect 11521 6847 11522 6873
rect 11494 6846 11522 6847
rect 11830 6846 11858 6874
rect 20006 8078 20034 8106
rect 18830 7574 18858 7602
rect 17598 7461 17626 7462
rect 17598 7435 17599 7461
rect 17599 7435 17625 7461
rect 17625 7435 17626 7461
rect 17598 7434 17626 7435
rect 17650 7461 17678 7462
rect 17650 7435 17651 7461
rect 17651 7435 17677 7461
rect 17677 7435 17678 7461
rect 17650 7434 17678 7435
rect 17702 7461 17730 7462
rect 17702 7435 17703 7461
rect 17703 7435 17729 7461
rect 17729 7435 17730 7461
rect 17702 7434 17730 7435
rect 11494 6734 11522 6762
rect 11942 6734 11970 6762
rect 2238 1973 2266 1974
rect 2238 1947 2239 1973
rect 2239 1947 2265 1973
rect 2265 1947 2266 1973
rect 2238 1946 2266 1947
rect 2290 1973 2318 1974
rect 2290 1947 2291 1973
rect 2291 1947 2317 1973
rect 2317 1947 2318 1973
rect 2290 1946 2318 1947
rect 2342 1973 2370 1974
rect 2342 1947 2343 1973
rect 2343 1947 2369 1973
rect 2369 1947 2370 1973
rect 2342 1946 2370 1947
rect 10766 2030 10794 2058
rect 9918 1581 9946 1582
rect 9918 1555 9919 1581
rect 9919 1555 9945 1581
rect 9945 1555 9946 1581
rect 9918 1554 9946 1555
rect 9970 1581 9998 1582
rect 9970 1555 9971 1581
rect 9971 1555 9997 1581
rect 9997 1555 9998 1581
rect 9970 1554 9998 1555
rect 10022 1581 10050 1582
rect 10022 1555 10023 1581
rect 10023 1555 10049 1581
rect 10049 1555 10050 1581
rect 10022 1554 10050 1555
rect 11382 2057 11410 2058
rect 11382 2031 11383 2057
rect 11383 2031 11409 2057
rect 11409 2031 11410 2057
rect 11382 2030 11410 2031
rect 17598 6677 17626 6678
rect 17598 6651 17599 6677
rect 17599 6651 17625 6677
rect 17625 6651 17626 6677
rect 17598 6650 17626 6651
rect 17650 6677 17678 6678
rect 17650 6651 17651 6677
rect 17651 6651 17677 6677
rect 17677 6651 17678 6677
rect 17650 6650 17678 6651
rect 17702 6677 17730 6678
rect 17702 6651 17703 6677
rect 17703 6651 17729 6677
rect 17729 6651 17730 6677
rect 17702 6650 17730 6651
rect 17598 5893 17626 5894
rect 17598 5867 17599 5893
rect 17599 5867 17625 5893
rect 17625 5867 17626 5893
rect 17598 5866 17626 5867
rect 17650 5893 17678 5894
rect 17650 5867 17651 5893
rect 17651 5867 17677 5893
rect 17677 5867 17678 5893
rect 17650 5866 17678 5867
rect 17702 5893 17730 5894
rect 17702 5867 17703 5893
rect 17703 5867 17729 5893
rect 17729 5867 17730 5893
rect 17702 5866 17730 5867
rect 17598 5109 17626 5110
rect 17598 5083 17599 5109
rect 17599 5083 17625 5109
rect 17625 5083 17626 5109
rect 17598 5082 17626 5083
rect 17650 5109 17678 5110
rect 17650 5083 17651 5109
rect 17651 5083 17677 5109
rect 17677 5083 17678 5109
rect 17650 5082 17678 5083
rect 17702 5109 17730 5110
rect 17702 5083 17703 5109
rect 17703 5083 17729 5109
rect 17729 5083 17730 5109
rect 17702 5082 17730 5083
rect 17598 4325 17626 4326
rect 17598 4299 17599 4325
rect 17599 4299 17625 4325
rect 17625 4299 17626 4325
rect 17598 4298 17626 4299
rect 17650 4325 17678 4326
rect 17650 4299 17651 4325
rect 17651 4299 17677 4325
rect 17677 4299 17678 4325
rect 17650 4298 17678 4299
rect 17702 4325 17730 4326
rect 17702 4299 17703 4325
rect 17703 4299 17729 4325
rect 17729 4299 17730 4325
rect 17702 4298 17730 4299
rect 17598 3541 17626 3542
rect 17598 3515 17599 3541
rect 17599 3515 17625 3541
rect 17625 3515 17626 3541
rect 17598 3514 17626 3515
rect 17650 3541 17678 3542
rect 17650 3515 17651 3541
rect 17651 3515 17677 3541
rect 17677 3515 17678 3541
rect 17650 3514 17678 3515
rect 17702 3541 17730 3542
rect 17702 3515 17703 3541
rect 17703 3515 17729 3541
rect 17729 3515 17730 3541
rect 17702 3514 17730 3515
rect 17598 2757 17626 2758
rect 17598 2731 17599 2757
rect 17599 2731 17625 2757
rect 17625 2731 17626 2757
rect 17598 2730 17626 2731
rect 17650 2757 17678 2758
rect 17650 2731 17651 2757
rect 17651 2731 17677 2757
rect 17677 2731 17678 2757
rect 17650 2730 17678 2731
rect 17702 2757 17730 2758
rect 17702 2731 17703 2757
rect 17703 2731 17729 2757
rect 17729 2731 17730 2757
rect 17702 2730 17730 2731
rect 13118 2030 13146 2058
rect 13734 2057 13762 2058
rect 13734 2031 13735 2057
rect 13735 2031 13761 2057
rect 13761 2031 13762 2057
rect 13734 2030 13762 2031
rect 17598 1973 17626 1974
rect 17598 1947 17599 1973
rect 17599 1947 17625 1973
rect 17625 1947 17626 1973
rect 17598 1946 17626 1947
rect 17650 1973 17678 1974
rect 17650 1947 17651 1973
rect 17651 1947 17677 1973
rect 17677 1947 17678 1973
rect 17650 1946 17678 1947
rect 17702 1973 17730 1974
rect 17702 1947 17703 1973
rect 17703 1947 17729 1973
rect 17729 1947 17730 1973
rect 17702 1946 17730 1947
<< metal3 >>
rect 12777 19278 12782 19306
rect 12810 19278 13398 19306
rect 13426 19278 13431 19306
rect 2233 19194 2238 19222
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2370 19194 2375 19222
rect 17593 19194 17598 19222
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17730 19194 17735 19222
rect 8409 19110 8414 19138
rect 8442 19110 9030 19138
rect 9058 19110 9063 19138
rect 10089 19110 10094 19138
rect 10122 19110 10878 19138
rect 10906 19110 10911 19138
rect 11433 19110 11438 19138
rect 11466 19110 12782 19138
rect 12810 19110 12815 19138
rect 13113 19110 13118 19138
rect 13146 19110 14686 19138
rect 14714 19110 14719 19138
rect 9913 18802 9918 18830
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 10050 18802 10055 18830
rect 9417 18718 9422 18746
rect 9450 18718 10038 18746
rect 10066 18718 10071 18746
rect 2233 18410 2238 18438
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2370 18410 2375 18438
rect 17593 18410 17598 18438
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17730 18410 17735 18438
rect 9913 18018 9918 18046
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 10050 18018 10055 18046
rect 2233 17626 2238 17654
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2370 17626 2375 17654
rect 17593 17626 17598 17654
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17730 17626 17735 17654
rect 9913 17234 9918 17262
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 10050 17234 10055 17262
rect 2233 16842 2238 16870
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2370 16842 2375 16870
rect 17593 16842 17598 16870
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17730 16842 17735 16870
rect 9913 16450 9918 16478
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 10050 16450 10055 16478
rect 2233 16058 2238 16086
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2370 16058 2375 16086
rect 17593 16058 17598 16086
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17730 16058 17735 16086
rect 9913 15666 9918 15694
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 10050 15666 10055 15694
rect 2233 15274 2238 15302
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2370 15274 2375 15302
rect 17593 15274 17598 15302
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17730 15274 17735 15302
rect 9913 14882 9918 14910
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 10050 14882 10055 14910
rect 2233 14490 2238 14518
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2370 14490 2375 14518
rect 17593 14490 17598 14518
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17730 14490 17735 14518
rect 7625 14294 7630 14322
rect 7658 14294 8134 14322
rect 8162 14294 8414 14322
rect 8442 14294 8918 14322
rect 8946 14294 9758 14322
rect 9786 14294 9791 14322
rect 10705 14294 10710 14322
rect 10738 14294 11830 14322
rect 11858 14294 12334 14322
rect 12362 14294 12367 14322
rect 8465 14238 8470 14266
rect 8498 14238 8974 14266
rect 9002 14238 9007 14266
rect 13225 14182 13230 14210
rect 13258 14182 14294 14210
rect 14322 14182 14327 14210
rect 0 14154 400 14168
rect 0 14126 2086 14154
rect 2114 14126 2119 14154
rect 0 14112 400 14126
rect 9913 14098 9918 14126
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 10050 14098 10055 14126
rect 11265 14014 11270 14042
rect 11298 14014 12110 14042
rect 12138 14014 12143 14042
rect 10761 13958 10766 13986
rect 10794 13958 11158 13986
rect 11186 13958 11191 13986
rect 11321 13902 11326 13930
rect 11354 13902 12110 13930
rect 12138 13902 12143 13930
rect 9249 13846 9254 13874
rect 9282 13846 9590 13874
rect 9618 13846 9623 13874
rect 2233 13706 2238 13734
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2370 13706 2375 13734
rect 17593 13706 17598 13734
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17730 13706 17735 13734
rect 12833 13566 12838 13594
rect 12866 13566 13230 13594
rect 13258 13566 13263 13594
rect 9473 13510 9478 13538
rect 9506 13510 11326 13538
rect 11354 13510 11359 13538
rect 9913 13314 9918 13342
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 10050 13314 10055 13342
rect 7401 13230 7406 13258
rect 7434 13230 7910 13258
rect 7938 13230 7943 13258
rect 8801 13230 8806 13258
rect 8834 13230 9366 13258
rect 9394 13230 9399 13258
rect 9977 13230 9982 13258
rect 10010 13230 10318 13258
rect 10346 13230 10351 13258
rect 11433 13230 11438 13258
rect 11466 13230 11886 13258
rect 11914 13230 11919 13258
rect 2137 13118 2142 13146
rect 2170 13118 5502 13146
rect 5530 13118 6790 13146
rect 6818 13118 6823 13146
rect 9025 13118 9030 13146
rect 9058 13118 9422 13146
rect 9450 13118 9758 13146
rect 9786 13118 9791 13146
rect 12217 13118 12222 13146
rect 12250 13118 12782 13146
rect 12810 13118 12815 13146
rect 7961 13062 7966 13090
rect 7994 13062 8862 13090
rect 8890 13062 8895 13090
rect 11377 13062 11382 13090
rect 11410 13062 11998 13090
rect 12026 13062 12390 13090
rect 12418 13062 12423 13090
rect 6561 13006 6566 13034
rect 6594 13006 7182 13034
rect 7210 13006 7215 13034
rect 2233 12922 2238 12950
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2370 12922 2375 12950
rect 17593 12922 17598 12950
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17730 12922 17735 12950
rect 10929 12838 10934 12866
rect 10962 12838 11438 12866
rect 11466 12838 11471 12866
rect 0 12810 400 12824
rect 20600 12810 21000 12824
rect 0 12782 966 12810
rect 994 12782 999 12810
rect 19945 12782 19950 12810
rect 19978 12782 21000 12810
rect 0 12768 400 12782
rect 20600 12768 21000 12782
rect 7289 12726 7294 12754
rect 7322 12726 10654 12754
rect 10682 12726 11158 12754
rect 11186 12726 11191 12754
rect 18825 12726 18830 12754
rect 18858 12726 18863 12754
rect 9865 12670 9870 12698
rect 9898 12670 10094 12698
rect 10122 12670 11550 12698
rect 11578 12670 11583 12698
rect 11825 12670 11830 12698
rect 11858 12670 12726 12698
rect 12754 12670 12759 12698
rect 12945 12670 12950 12698
rect 12978 12670 13902 12698
rect 13930 12670 13935 12698
rect 14737 12670 14742 12698
rect 14770 12670 18718 12698
rect 18746 12670 18751 12698
rect 18830 12642 18858 12726
rect 9193 12614 9198 12642
rect 9226 12614 9590 12642
rect 9618 12614 9623 12642
rect 11377 12614 11382 12642
rect 11410 12614 13006 12642
rect 13034 12614 13039 12642
rect 14625 12614 14630 12642
rect 14658 12614 14854 12642
rect 14882 12614 18858 12642
rect 14630 12586 14658 12614
rect 13118 12558 14658 12586
rect 9913 12530 9918 12558
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 10050 12530 10055 12558
rect 13118 12530 13146 12558
rect 13113 12502 13118 12530
rect 13146 12502 13151 12530
rect 20600 12474 21000 12488
rect 6505 12446 6510 12474
rect 6538 12446 6846 12474
rect 6874 12446 7238 12474
rect 7266 12446 7271 12474
rect 20001 12446 20006 12474
rect 20034 12446 21000 12474
rect 20600 12432 21000 12446
rect 6729 12390 6734 12418
rect 6762 12390 7126 12418
rect 7154 12390 11662 12418
rect 11690 12390 11695 12418
rect 12105 12390 12110 12418
rect 12138 12390 12782 12418
rect 12810 12390 12815 12418
rect 11881 12334 11886 12362
rect 11914 12334 12222 12362
rect 12250 12334 13006 12362
rect 13034 12334 13039 12362
rect 13225 12334 13230 12362
rect 13258 12334 13846 12362
rect 13874 12334 13879 12362
rect 13230 12306 13258 12334
rect 11545 12278 11550 12306
rect 11578 12278 13258 12306
rect 8073 12222 8078 12250
rect 8106 12222 8918 12250
rect 8946 12222 9646 12250
rect 9674 12222 9679 12250
rect 9809 12222 9814 12250
rect 9842 12222 10150 12250
rect 10178 12222 10183 12250
rect 2233 12138 2238 12166
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2370 12138 2375 12166
rect 17593 12138 17598 12166
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17730 12138 17735 12166
rect 8689 11998 8694 12026
rect 8722 11998 9310 12026
rect 9338 11998 9343 12026
rect 9529 11998 9534 12026
rect 9562 11998 9982 12026
rect 10010 11998 12614 12026
rect 12642 11998 12647 12026
rect 2137 11942 2142 11970
rect 2170 11942 4214 11970
rect 9081 11942 9086 11970
rect 9114 11942 10094 11970
rect 10122 11942 10127 11970
rect 13897 11942 13902 11970
rect 13930 11942 14742 11970
rect 14770 11942 18830 11970
rect 18858 11942 18863 11970
rect 4186 11914 4214 11942
rect 4186 11886 4942 11914
rect 4970 11886 6790 11914
rect 6818 11886 6823 11914
rect 9473 11886 9478 11914
rect 9506 11886 10038 11914
rect 10066 11886 10071 11914
rect 10201 11886 10206 11914
rect 10234 11886 10850 11914
rect 11097 11886 11102 11914
rect 11130 11886 11942 11914
rect 11970 11886 11975 11914
rect 10822 11858 10850 11886
rect 9809 11830 9814 11858
rect 9842 11830 10262 11858
rect 10290 11830 10295 11858
rect 10817 11830 10822 11858
rect 10850 11830 11270 11858
rect 11298 11830 11303 11858
rect 11657 11830 11662 11858
rect 11690 11830 12782 11858
rect 12810 11830 12815 11858
rect 13057 11830 13062 11858
rect 13090 11830 14014 11858
rect 14042 11830 14047 11858
rect 0 11802 400 11816
rect 20600 11802 21000 11816
rect 0 11774 966 11802
rect 994 11774 999 11802
rect 6001 11774 6006 11802
rect 6034 11774 6846 11802
rect 6874 11774 6879 11802
rect 10089 11774 10094 11802
rect 10122 11774 10710 11802
rect 10738 11774 11438 11802
rect 11466 11774 11471 11802
rect 12665 11774 12670 11802
rect 12698 11774 13006 11802
rect 13034 11774 13286 11802
rect 13314 11774 13319 11802
rect 20001 11774 20006 11802
rect 20034 11774 21000 11802
rect 0 11760 400 11774
rect 9913 11746 9918 11774
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 10050 11746 10055 11774
rect 20600 11760 21000 11774
rect 9193 11718 9198 11746
rect 9226 11718 9758 11746
rect 9786 11718 9791 11746
rect 6281 11606 6286 11634
rect 6314 11606 7014 11634
rect 7042 11606 7047 11634
rect 11209 11606 11214 11634
rect 11242 11606 11662 11634
rect 11690 11606 11695 11634
rect 9025 11550 9030 11578
rect 9058 11550 10654 11578
rect 10682 11550 11606 11578
rect 11634 11550 13006 11578
rect 13034 11550 13039 11578
rect 9697 11494 9702 11522
rect 9730 11494 9926 11522
rect 9954 11494 10374 11522
rect 10402 11494 10878 11522
rect 10906 11494 10911 11522
rect 11321 11494 11326 11522
rect 11354 11494 11718 11522
rect 11746 11494 11751 11522
rect 12889 11494 12894 11522
rect 12922 11494 13678 11522
rect 13706 11494 13711 11522
rect 10201 11438 10206 11466
rect 10234 11438 12950 11466
rect 12978 11438 12983 11466
rect 2233 11354 2238 11382
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2370 11354 2375 11382
rect 17593 11354 17598 11382
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17730 11354 17735 11382
rect 11377 11270 11382 11298
rect 11410 11270 11774 11298
rect 11802 11270 11807 11298
rect 961 11214 966 11242
rect 994 11214 999 11242
rect 0 11130 400 11144
rect 966 11130 994 11214
rect 2137 11158 2142 11186
rect 2170 11158 5670 11186
rect 5698 11158 5703 11186
rect 7009 11158 7014 11186
rect 7042 11158 7910 11186
rect 7938 11158 7943 11186
rect 0 11102 994 11130
rect 10873 11102 10878 11130
rect 10906 11102 11438 11130
rect 11466 11102 11471 11130
rect 0 11088 400 11102
rect 9025 10990 9030 11018
rect 9058 10990 9142 11018
rect 9170 10990 9175 11018
rect 9913 10962 9918 10990
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 10050 10962 10055 10990
rect 7233 10934 7238 10962
rect 7266 10934 8750 10962
rect 8778 10934 9142 10962
rect 9170 10934 9175 10962
rect 7345 10878 7350 10906
rect 7378 10878 7742 10906
rect 7770 10878 7775 10906
rect 9249 10878 9254 10906
rect 9282 10878 9758 10906
rect 9786 10878 10150 10906
rect 10178 10878 10183 10906
rect 5665 10822 5670 10850
rect 5698 10822 7686 10850
rect 7714 10822 7719 10850
rect 8969 10822 8974 10850
rect 9002 10822 9534 10850
rect 9562 10822 9567 10850
rect 2081 10766 2086 10794
rect 2114 10766 9590 10794
rect 9618 10766 10710 10794
rect 10738 10766 10743 10794
rect 9123 10710 9142 10738
rect 9170 10710 9175 10738
rect 9697 10710 9702 10738
rect 9730 10710 11326 10738
rect 11354 10710 11359 10738
rect 13057 10654 13062 10682
rect 13090 10654 14518 10682
rect 14546 10654 14551 10682
rect 7569 10598 7574 10626
rect 7602 10598 8246 10626
rect 8274 10598 8279 10626
rect 9137 10598 9142 10626
rect 9170 10598 10934 10626
rect 10962 10598 10967 10626
rect 2233 10570 2238 10598
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2370 10570 2375 10598
rect 17593 10570 17598 10598
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17730 10570 17735 10598
rect 7121 10542 7126 10570
rect 7154 10542 8190 10570
rect 8218 10542 8223 10570
rect 10313 10542 10318 10570
rect 10346 10542 10878 10570
rect 10906 10542 11214 10570
rect 11242 10542 11438 10570
rect 11466 10542 11471 10570
rect 0 10458 400 10472
rect 20600 10458 21000 10472
rect 0 10430 966 10458
rect 994 10430 999 10458
rect 11097 10430 11102 10458
rect 11130 10430 12446 10458
rect 12474 10430 12479 10458
rect 20001 10430 20006 10458
rect 20034 10430 21000 10458
rect 0 10416 400 10430
rect 20600 10416 21000 10430
rect 9193 10374 9198 10402
rect 9226 10374 10318 10402
rect 10346 10374 10351 10402
rect 2137 10318 2142 10346
rect 2170 10318 4214 10346
rect 8857 10318 8862 10346
rect 8890 10318 10094 10346
rect 10122 10318 11102 10346
rect 11130 10318 11135 10346
rect 4186 10290 4214 10318
rect 4186 10262 4830 10290
rect 4858 10262 6062 10290
rect 6090 10262 6095 10290
rect 8297 10262 8302 10290
rect 8330 10262 9142 10290
rect 9170 10262 9175 10290
rect 9366 10262 11158 10290
rect 11186 10262 11191 10290
rect 9366 10234 9394 10262
rect 7961 10206 7966 10234
rect 7994 10206 9366 10234
rect 9394 10206 9399 10234
rect 9913 10178 9918 10206
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 10050 10178 10055 10206
rect 11601 10150 11606 10178
rect 11634 10150 12558 10178
rect 12586 10150 12591 10178
rect 20600 10122 21000 10136
rect 7737 10094 7742 10122
rect 7770 10094 8134 10122
rect 8162 10094 8167 10122
rect 11769 10094 11774 10122
rect 11802 10094 12054 10122
rect 12082 10094 12278 10122
rect 12306 10094 12311 10122
rect 14905 10094 14910 10122
rect 14938 10094 18830 10122
rect 18858 10094 18863 10122
rect 20113 10094 20118 10122
rect 20146 10094 21000 10122
rect 20600 10080 21000 10094
rect 6281 10038 6286 10066
rect 6314 10038 6790 10066
rect 6818 10038 7014 10066
rect 7042 10038 7350 10066
rect 7378 10038 8470 10066
rect 8498 10038 8503 10066
rect 8633 10038 8638 10066
rect 8666 10038 8750 10066
rect 8778 10038 9142 10066
rect 9170 10038 9310 10066
rect 9338 10038 9343 10066
rect 12385 10038 12390 10066
rect 12418 10038 12838 10066
rect 12866 10038 13174 10066
rect 13202 10038 13207 10066
rect 8969 9982 8974 10010
rect 9002 9982 10094 10010
rect 10122 9982 10127 10010
rect 12497 9982 12502 10010
rect 12530 9982 12950 10010
rect 12978 9982 12983 10010
rect 6561 9926 6566 9954
rect 6594 9926 9366 9954
rect 9394 9926 9982 9954
rect 10010 9926 10015 9954
rect 11321 9926 11326 9954
rect 11354 9926 11662 9954
rect 11690 9926 11695 9954
rect 12665 9926 12670 9954
rect 12698 9926 12838 9954
rect 12866 9926 12871 9954
rect 13001 9926 13006 9954
rect 13034 9926 13846 9954
rect 13874 9926 13879 9954
rect 8801 9870 8806 9898
rect 8834 9870 10934 9898
rect 10962 9870 12614 9898
rect 12642 9870 12647 9898
rect 8913 9814 8918 9842
rect 8946 9814 11046 9842
rect 11074 9814 11079 9842
rect 2233 9786 2238 9814
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2370 9786 2375 9814
rect 17593 9786 17598 9814
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17730 9786 17735 9814
rect 20600 9786 21000 9800
rect 20001 9758 20006 9786
rect 20034 9758 21000 9786
rect 20600 9744 21000 9758
rect 9305 9702 9310 9730
rect 9338 9702 11270 9730
rect 11298 9702 11303 9730
rect 9361 9646 9366 9674
rect 9394 9646 10262 9674
rect 10290 9646 10878 9674
rect 10906 9646 10911 9674
rect 11881 9646 11886 9674
rect 11914 9646 12614 9674
rect 12642 9646 13286 9674
rect 13314 9646 13319 9674
rect 7793 9590 7798 9618
rect 7826 9590 9310 9618
rect 9338 9590 9343 9618
rect 9977 9590 9982 9618
rect 10010 9590 10598 9618
rect 10626 9590 10631 9618
rect 11041 9590 11046 9618
rect 11074 9590 12670 9618
rect 12698 9590 12703 9618
rect 7289 9534 7294 9562
rect 7322 9534 7518 9562
rect 7546 9534 8638 9562
rect 8666 9534 8918 9562
rect 8946 9534 8951 9562
rect 9753 9534 9758 9562
rect 9786 9534 10766 9562
rect 10794 9534 10799 9562
rect 11321 9534 11326 9562
rect 11354 9534 11942 9562
rect 11970 9534 11975 9562
rect 14289 9534 14294 9562
rect 14322 9534 14798 9562
rect 14826 9534 18830 9562
rect 18858 9534 18863 9562
rect 8129 9478 8134 9506
rect 8162 9478 8974 9506
rect 9002 9478 9007 9506
rect 10201 9478 10206 9506
rect 10234 9478 10990 9506
rect 11018 9478 11382 9506
rect 11410 9478 11998 9506
rect 12026 9478 12222 9506
rect 12250 9478 12255 9506
rect 11713 9422 11718 9450
rect 11746 9422 12446 9450
rect 12474 9422 12950 9450
rect 12978 9422 12983 9450
rect 9913 9394 9918 9422
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 10050 9394 10055 9422
rect 12049 9366 12054 9394
rect 12082 9366 13006 9394
rect 13034 9366 13398 9394
rect 13426 9366 13431 9394
rect 7546 9310 7686 9338
rect 7714 9310 7719 9338
rect 7793 9310 7798 9338
rect 7826 9310 9366 9338
rect 9394 9310 9399 9338
rect 9641 9310 9646 9338
rect 9674 9310 11046 9338
rect 11074 9310 11079 9338
rect 11153 9310 11158 9338
rect 11186 9310 11382 9338
rect 11410 9310 11494 9338
rect 11522 9310 11527 9338
rect 11993 9310 11998 9338
rect 12026 9310 12502 9338
rect 12530 9310 12535 9338
rect 7546 9282 7574 9310
rect 7401 9254 7406 9282
rect 7434 9254 7574 9282
rect 10761 9254 10766 9282
rect 10794 9254 13510 9282
rect 13538 9254 13543 9282
rect 11102 9226 11130 9254
rect 2137 9198 2142 9226
rect 2170 9198 5446 9226
rect 5474 9198 7014 9226
rect 7042 9198 7047 9226
rect 7350 9198 8834 9226
rect 8969 9198 8974 9226
rect 9002 9198 9926 9226
rect 9954 9198 9959 9226
rect 11097 9198 11102 9226
rect 11130 9198 11135 9226
rect 11209 9198 11214 9226
rect 11242 9198 11606 9226
rect 11634 9198 11639 9226
rect 7350 9170 7378 9198
rect 8806 9170 8834 9198
rect 7345 9142 7350 9170
rect 7378 9142 7383 9170
rect 8353 9142 8358 9170
rect 8386 9142 8694 9170
rect 8722 9142 8727 9170
rect 8806 9142 10038 9170
rect 10066 9142 12222 9170
rect 12250 9142 12255 9170
rect 0 9114 400 9128
rect 0 9086 966 9114
rect 994 9086 999 9114
rect 6337 9086 6342 9114
rect 6370 9086 7070 9114
rect 7098 9086 7103 9114
rect 8409 9086 8414 9114
rect 8442 9086 9030 9114
rect 9058 9086 9063 9114
rect 10929 9086 10934 9114
rect 10962 9086 12166 9114
rect 12194 9086 12614 9114
rect 12642 9086 12647 9114
rect 0 9072 400 9086
rect 2233 9002 2238 9030
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2370 9002 2375 9030
rect 17593 9002 17598 9030
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17730 9002 17735 9030
rect 10817 8918 10822 8946
rect 10850 8918 11158 8946
rect 11186 8918 11191 8946
rect 961 8862 966 8890
rect 994 8862 999 8890
rect 12665 8862 12670 8890
rect 12698 8862 13230 8890
rect 13258 8862 13263 8890
rect 13953 8862 13958 8890
rect 13986 8862 14294 8890
rect 14322 8862 15974 8890
rect 0 8778 400 8792
rect 966 8778 994 8862
rect 15946 8834 15974 8862
rect 2137 8806 2142 8834
rect 2170 8806 6846 8834
rect 6874 8806 6879 8834
rect 12833 8806 12838 8834
rect 12866 8806 13398 8834
rect 13426 8806 14630 8834
rect 14658 8806 14663 8834
rect 15946 8806 18830 8834
rect 18858 8806 18863 8834
rect 20600 8778 21000 8792
rect 0 8750 994 8778
rect 12609 8750 12614 8778
rect 12642 8750 13902 8778
rect 13930 8750 13935 8778
rect 20001 8750 20006 8778
rect 20034 8750 21000 8778
rect 0 8736 400 8750
rect 20600 8736 21000 8750
rect 12385 8694 12390 8722
rect 12418 8694 12894 8722
rect 12922 8694 12927 8722
rect 9913 8610 9918 8638
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 10050 8610 10055 8638
rect 11937 8582 11942 8610
rect 11970 8582 12334 8610
rect 12362 8582 12838 8610
rect 12866 8582 12871 8610
rect 9473 8470 9478 8498
rect 9506 8470 9982 8498
rect 10010 8470 10015 8498
rect 11657 8470 11662 8498
rect 11690 8470 12950 8498
rect 12978 8470 12983 8498
rect 8185 8414 8190 8442
rect 8218 8414 9254 8442
rect 9282 8414 11886 8442
rect 11914 8414 11919 8442
rect 8689 8358 8694 8386
rect 8722 8358 9590 8386
rect 9618 8358 9623 8386
rect 9697 8358 9702 8386
rect 9730 8358 10486 8386
rect 10514 8358 10519 8386
rect 10705 8358 10710 8386
rect 10738 8358 11830 8386
rect 11858 8358 11863 8386
rect 12329 8358 12334 8386
rect 12362 8358 12670 8386
rect 12698 8358 12703 8386
rect 11830 8330 11858 8358
rect 9977 8302 9982 8330
rect 10010 8302 11326 8330
rect 11354 8302 11359 8330
rect 11830 8302 12614 8330
rect 12642 8302 12647 8330
rect 2233 8218 2238 8246
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2370 8218 2375 8246
rect 17593 8218 17598 8246
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17730 8218 17735 8246
rect 20600 8106 21000 8120
rect 20001 8078 20006 8106
rect 20034 8078 21000 8106
rect 20600 8064 21000 8078
rect 9913 7826 9918 7854
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 10050 7826 10055 7854
rect 11769 7742 11774 7770
rect 11802 7742 12838 7770
rect 12866 7742 12871 7770
rect 9697 7630 9702 7658
rect 9730 7630 10598 7658
rect 10626 7630 10934 7658
rect 10962 7630 10967 7658
rect 10873 7574 10878 7602
rect 10906 7574 11382 7602
rect 11410 7574 11415 7602
rect 12217 7574 12222 7602
rect 12250 7574 12670 7602
rect 12698 7574 12703 7602
rect 13113 7574 13118 7602
rect 13146 7574 13398 7602
rect 13426 7574 18830 7602
rect 18858 7574 18863 7602
rect 2233 7434 2238 7462
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2370 7434 2375 7462
rect 17593 7434 17598 7462
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17730 7434 17735 7462
rect 8353 7238 8358 7266
rect 8386 7238 8750 7266
rect 8778 7238 9982 7266
rect 10010 7238 10015 7266
rect 9913 7042 9918 7070
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 10050 7042 10055 7070
rect 9865 6846 9870 6874
rect 9898 6846 11158 6874
rect 11186 6846 11494 6874
rect 11522 6846 11830 6874
rect 11858 6846 11863 6874
rect 11265 6734 11270 6762
rect 11298 6734 11494 6762
rect 11522 6734 11942 6762
rect 11970 6734 11975 6762
rect 2233 6650 2238 6678
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2370 6650 2375 6678
rect 17593 6650 17598 6678
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17730 6650 17735 6678
rect 9913 6258 9918 6286
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 10050 6258 10055 6286
rect 2233 5866 2238 5894
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2370 5866 2375 5894
rect 17593 5866 17598 5894
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17730 5866 17735 5894
rect 9913 5474 9918 5502
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 10050 5474 10055 5502
rect 2233 5082 2238 5110
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2370 5082 2375 5110
rect 17593 5082 17598 5110
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17730 5082 17735 5110
rect 9913 4690 9918 4718
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 10050 4690 10055 4718
rect 2233 4298 2238 4326
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2370 4298 2375 4326
rect 17593 4298 17598 4326
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17730 4298 17735 4326
rect 9913 3906 9918 3934
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 10050 3906 10055 3934
rect 2233 3514 2238 3542
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2370 3514 2375 3542
rect 17593 3514 17598 3542
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17730 3514 17735 3542
rect 9913 3122 9918 3150
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 10050 3122 10055 3150
rect 2233 2730 2238 2758
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2370 2730 2375 2758
rect 17593 2730 17598 2758
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17730 2730 17735 2758
rect 9913 2338 9918 2366
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 10050 2338 10055 2366
rect 10761 2030 10766 2058
rect 10794 2030 11382 2058
rect 11410 2030 11415 2058
rect 13113 2030 13118 2058
rect 13146 2030 13734 2058
rect 13762 2030 13767 2058
rect 2233 1946 2238 1974
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2370 1946 2375 1974
rect 17593 1946 17598 1974
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17730 1946 17735 1974
rect 9913 1554 9918 1582
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 10050 1554 10055 1582
<< via3 >>
rect 2238 19194 2266 19222
rect 2290 19194 2318 19222
rect 2342 19194 2370 19222
rect 17598 19194 17626 19222
rect 17650 19194 17678 19222
rect 17702 19194 17730 19222
rect 9918 18802 9946 18830
rect 9970 18802 9998 18830
rect 10022 18802 10050 18830
rect 2238 18410 2266 18438
rect 2290 18410 2318 18438
rect 2342 18410 2370 18438
rect 17598 18410 17626 18438
rect 17650 18410 17678 18438
rect 17702 18410 17730 18438
rect 9918 18018 9946 18046
rect 9970 18018 9998 18046
rect 10022 18018 10050 18046
rect 2238 17626 2266 17654
rect 2290 17626 2318 17654
rect 2342 17626 2370 17654
rect 17598 17626 17626 17654
rect 17650 17626 17678 17654
rect 17702 17626 17730 17654
rect 9918 17234 9946 17262
rect 9970 17234 9998 17262
rect 10022 17234 10050 17262
rect 2238 16842 2266 16870
rect 2290 16842 2318 16870
rect 2342 16842 2370 16870
rect 17598 16842 17626 16870
rect 17650 16842 17678 16870
rect 17702 16842 17730 16870
rect 9918 16450 9946 16478
rect 9970 16450 9998 16478
rect 10022 16450 10050 16478
rect 2238 16058 2266 16086
rect 2290 16058 2318 16086
rect 2342 16058 2370 16086
rect 17598 16058 17626 16086
rect 17650 16058 17678 16086
rect 17702 16058 17730 16086
rect 9918 15666 9946 15694
rect 9970 15666 9998 15694
rect 10022 15666 10050 15694
rect 2238 15274 2266 15302
rect 2290 15274 2318 15302
rect 2342 15274 2370 15302
rect 17598 15274 17626 15302
rect 17650 15274 17678 15302
rect 17702 15274 17730 15302
rect 9918 14882 9946 14910
rect 9970 14882 9998 14910
rect 10022 14882 10050 14910
rect 2238 14490 2266 14518
rect 2290 14490 2318 14518
rect 2342 14490 2370 14518
rect 17598 14490 17626 14518
rect 17650 14490 17678 14518
rect 17702 14490 17730 14518
rect 9918 14098 9946 14126
rect 9970 14098 9998 14126
rect 10022 14098 10050 14126
rect 2238 13706 2266 13734
rect 2290 13706 2318 13734
rect 2342 13706 2370 13734
rect 17598 13706 17626 13734
rect 17650 13706 17678 13734
rect 17702 13706 17730 13734
rect 9918 13314 9946 13342
rect 9970 13314 9998 13342
rect 10022 13314 10050 13342
rect 2238 12922 2266 12950
rect 2290 12922 2318 12950
rect 2342 12922 2370 12950
rect 17598 12922 17626 12950
rect 17650 12922 17678 12950
rect 17702 12922 17730 12950
rect 9918 12530 9946 12558
rect 9970 12530 9998 12558
rect 10022 12530 10050 12558
rect 2238 12138 2266 12166
rect 2290 12138 2318 12166
rect 2342 12138 2370 12166
rect 17598 12138 17626 12166
rect 17650 12138 17678 12166
rect 17702 12138 17730 12166
rect 9918 11746 9946 11774
rect 9970 11746 9998 11774
rect 10022 11746 10050 11774
rect 2238 11354 2266 11382
rect 2290 11354 2318 11382
rect 2342 11354 2370 11382
rect 17598 11354 17626 11382
rect 17650 11354 17678 11382
rect 17702 11354 17730 11382
rect 9142 10990 9170 11018
rect 9918 10962 9946 10990
rect 9970 10962 9998 10990
rect 10022 10962 10050 10990
rect 9142 10710 9170 10738
rect 2238 10570 2266 10598
rect 2290 10570 2318 10598
rect 2342 10570 2370 10598
rect 17598 10570 17626 10598
rect 17650 10570 17678 10598
rect 17702 10570 17730 10598
rect 9918 10178 9946 10206
rect 9970 10178 9998 10206
rect 10022 10178 10050 10206
rect 2238 9786 2266 9814
rect 2290 9786 2318 9814
rect 2342 9786 2370 9814
rect 17598 9786 17626 9814
rect 17650 9786 17678 9814
rect 17702 9786 17730 9814
rect 9918 9394 9946 9422
rect 9970 9394 9998 9422
rect 10022 9394 10050 9422
rect 2238 9002 2266 9030
rect 2290 9002 2318 9030
rect 2342 9002 2370 9030
rect 17598 9002 17626 9030
rect 17650 9002 17678 9030
rect 17702 9002 17730 9030
rect 9918 8610 9946 8638
rect 9970 8610 9998 8638
rect 10022 8610 10050 8638
rect 2238 8218 2266 8246
rect 2290 8218 2318 8246
rect 2342 8218 2370 8246
rect 17598 8218 17626 8246
rect 17650 8218 17678 8246
rect 17702 8218 17730 8246
rect 9918 7826 9946 7854
rect 9970 7826 9998 7854
rect 10022 7826 10050 7854
rect 2238 7434 2266 7462
rect 2290 7434 2318 7462
rect 2342 7434 2370 7462
rect 17598 7434 17626 7462
rect 17650 7434 17678 7462
rect 17702 7434 17730 7462
rect 9918 7042 9946 7070
rect 9970 7042 9998 7070
rect 10022 7042 10050 7070
rect 2238 6650 2266 6678
rect 2290 6650 2318 6678
rect 2342 6650 2370 6678
rect 17598 6650 17626 6678
rect 17650 6650 17678 6678
rect 17702 6650 17730 6678
rect 9918 6258 9946 6286
rect 9970 6258 9998 6286
rect 10022 6258 10050 6286
rect 2238 5866 2266 5894
rect 2290 5866 2318 5894
rect 2342 5866 2370 5894
rect 17598 5866 17626 5894
rect 17650 5866 17678 5894
rect 17702 5866 17730 5894
rect 9918 5474 9946 5502
rect 9970 5474 9998 5502
rect 10022 5474 10050 5502
rect 2238 5082 2266 5110
rect 2290 5082 2318 5110
rect 2342 5082 2370 5110
rect 17598 5082 17626 5110
rect 17650 5082 17678 5110
rect 17702 5082 17730 5110
rect 9918 4690 9946 4718
rect 9970 4690 9998 4718
rect 10022 4690 10050 4718
rect 2238 4298 2266 4326
rect 2290 4298 2318 4326
rect 2342 4298 2370 4326
rect 17598 4298 17626 4326
rect 17650 4298 17678 4326
rect 17702 4298 17730 4326
rect 9918 3906 9946 3934
rect 9970 3906 9998 3934
rect 10022 3906 10050 3934
rect 2238 3514 2266 3542
rect 2290 3514 2318 3542
rect 2342 3514 2370 3542
rect 17598 3514 17626 3542
rect 17650 3514 17678 3542
rect 17702 3514 17730 3542
rect 9918 3122 9946 3150
rect 9970 3122 9998 3150
rect 10022 3122 10050 3150
rect 2238 2730 2266 2758
rect 2290 2730 2318 2758
rect 2342 2730 2370 2758
rect 17598 2730 17626 2758
rect 17650 2730 17678 2758
rect 17702 2730 17730 2758
rect 9918 2338 9946 2366
rect 9970 2338 9998 2366
rect 10022 2338 10050 2366
rect 2238 1946 2266 1974
rect 2290 1946 2318 1974
rect 2342 1946 2370 1974
rect 17598 1946 17626 1974
rect 17650 1946 17678 1974
rect 17702 1946 17730 1974
rect 9918 1554 9946 1582
rect 9970 1554 9998 1582
rect 10022 1554 10050 1582
<< metal4 >>
rect 2224 19222 2384 19238
rect 2224 19194 2238 19222
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2370 19194 2384 19222
rect 2224 18438 2384 19194
rect 2224 18410 2238 18438
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2370 18410 2384 18438
rect 2224 17654 2384 18410
rect 2224 17626 2238 17654
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2370 17626 2384 17654
rect 2224 16870 2384 17626
rect 2224 16842 2238 16870
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2370 16842 2384 16870
rect 2224 16086 2384 16842
rect 2224 16058 2238 16086
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2370 16058 2384 16086
rect 2224 15302 2384 16058
rect 2224 15274 2238 15302
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2370 15274 2384 15302
rect 2224 14518 2384 15274
rect 2224 14490 2238 14518
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2370 14490 2384 14518
rect 2224 13734 2384 14490
rect 2224 13706 2238 13734
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2370 13706 2384 13734
rect 2224 12950 2384 13706
rect 2224 12922 2238 12950
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2370 12922 2384 12950
rect 2224 12166 2384 12922
rect 2224 12138 2238 12166
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2370 12138 2384 12166
rect 2224 11382 2384 12138
rect 2224 11354 2238 11382
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2370 11354 2384 11382
rect 2224 10598 2384 11354
rect 9904 18830 10064 19238
rect 9904 18802 9918 18830
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 10050 18802 10064 18830
rect 9904 18046 10064 18802
rect 9904 18018 9918 18046
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 10050 18018 10064 18046
rect 9904 17262 10064 18018
rect 9904 17234 9918 17262
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 10050 17234 10064 17262
rect 9904 16478 10064 17234
rect 9904 16450 9918 16478
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 10050 16450 10064 16478
rect 9904 15694 10064 16450
rect 9904 15666 9918 15694
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 10050 15666 10064 15694
rect 9904 14910 10064 15666
rect 9904 14882 9918 14910
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 10050 14882 10064 14910
rect 9904 14126 10064 14882
rect 9904 14098 9918 14126
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 10050 14098 10064 14126
rect 9904 13342 10064 14098
rect 9904 13314 9918 13342
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 10050 13314 10064 13342
rect 9904 12558 10064 13314
rect 9904 12530 9918 12558
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 10050 12530 10064 12558
rect 9904 11774 10064 12530
rect 9904 11746 9918 11774
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 10050 11746 10064 11774
rect 9142 11018 9170 11023
rect 9142 10738 9170 10990
rect 9142 10705 9170 10710
rect 9904 10990 10064 11746
rect 9904 10962 9918 10990
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 10050 10962 10064 10990
rect 2224 10570 2238 10598
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2370 10570 2384 10598
rect 2224 9814 2384 10570
rect 2224 9786 2238 9814
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2370 9786 2384 9814
rect 2224 9030 2384 9786
rect 2224 9002 2238 9030
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2370 9002 2384 9030
rect 2224 8246 2384 9002
rect 2224 8218 2238 8246
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2370 8218 2384 8246
rect 2224 7462 2384 8218
rect 2224 7434 2238 7462
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2370 7434 2384 7462
rect 2224 6678 2384 7434
rect 2224 6650 2238 6678
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2370 6650 2384 6678
rect 2224 5894 2384 6650
rect 2224 5866 2238 5894
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2370 5866 2384 5894
rect 2224 5110 2384 5866
rect 2224 5082 2238 5110
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2370 5082 2384 5110
rect 2224 4326 2384 5082
rect 2224 4298 2238 4326
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2370 4298 2384 4326
rect 2224 3542 2384 4298
rect 2224 3514 2238 3542
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2370 3514 2384 3542
rect 2224 2758 2384 3514
rect 2224 2730 2238 2758
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2370 2730 2384 2758
rect 2224 1974 2384 2730
rect 2224 1946 2238 1974
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2370 1946 2384 1974
rect 2224 1538 2384 1946
rect 9904 10206 10064 10962
rect 9904 10178 9918 10206
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 10050 10178 10064 10206
rect 9904 9422 10064 10178
rect 9904 9394 9918 9422
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 10050 9394 10064 9422
rect 9904 8638 10064 9394
rect 9904 8610 9918 8638
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 10050 8610 10064 8638
rect 9904 7854 10064 8610
rect 9904 7826 9918 7854
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 10050 7826 10064 7854
rect 9904 7070 10064 7826
rect 9904 7042 9918 7070
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 10050 7042 10064 7070
rect 9904 6286 10064 7042
rect 9904 6258 9918 6286
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 10050 6258 10064 6286
rect 9904 5502 10064 6258
rect 9904 5474 9918 5502
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 10050 5474 10064 5502
rect 9904 4718 10064 5474
rect 9904 4690 9918 4718
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 10050 4690 10064 4718
rect 9904 3934 10064 4690
rect 9904 3906 9918 3934
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 10050 3906 10064 3934
rect 9904 3150 10064 3906
rect 9904 3122 9918 3150
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 10050 3122 10064 3150
rect 9904 2366 10064 3122
rect 9904 2338 9918 2366
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 10050 2338 10064 2366
rect 9904 1582 10064 2338
rect 9904 1554 9918 1582
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 10050 1554 10064 1582
rect 9904 1538 10064 1554
rect 17584 19222 17744 19238
rect 17584 19194 17598 19222
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17730 19194 17744 19222
rect 17584 18438 17744 19194
rect 17584 18410 17598 18438
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17730 18410 17744 18438
rect 17584 17654 17744 18410
rect 17584 17626 17598 17654
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17730 17626 17744 17654
rect 17584 16870 17744 17626
rect 17584 16842 17598 16870
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17730 16842 17744 16870
rect 17584 16086 17744 16842
rect 17584 16058 17598 16086
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17730 16058 17744 16086
rect 17584 15302 17744 16058
rect 17584 15274 17598 15302
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17730 15274 17744 15302
rect 17584 14518 17744 15274
rect 17584 14490 17598 14518
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17730 14490 17744 14518
rect 17584 13734 17744 14490
rect 17584 13706 17598 13734
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17730 13706 17744 13734
rect 17584 12950 17744 13706
rect 17584 12922 17598 12950
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17730 12922 17744 12950
rect 17584 12166 17744 12922
rect 17584 12138 17598 12166
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17730 12138 17744 12166
rect 17584 11382 17744 12138
rect 17584 11354 17598 11382
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17730 11354 17744 11382
rect 17584 10598 17744 11354
rect 17584 10570 17598 10598
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17730 10570 17744 10598
rect 17584 9814 17744 10570
rect 17584 9786 17598 9814
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17730 9786 17744 9814
rect 17584 9030 17744 9786
rect 17584 9002 17598 9030
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17730 9002 17744 9030
rect 17584 8246 17744 9002
rect 17584 8218 17598 8246
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17730 8218 17744 8246
rect 17584 7462 17744 8218
rect 17584 7434 17598 7462
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17730 7434 17744 7462
rect 17584 6678 17744 7434
rect 17584 6650 17598 6678
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17730 6650 17744 6678
rect 17584 5894 17744 6650
rect 17584 5866 17598 5894
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17730 5866 17744 5894
rect 17584 5110 17744 5866
rect 17584 5082 17598 5110
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17730 5082 17744 5110
rect 17584 4326 17744 5082
rect 17584 4298 17598 4326
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17730 4298 17744 4326
rect 17584 3542 17744 4298
rect 17584 3514 17598 3542
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17730 3514 17744 3542
rect 17584 2758 17744 3514
rect 17584 2730 17598 2758
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17730 2730 17744 2758
rect 17584 1974 17744 2730
rect 17584 1946 17598 1974
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17730 1946 17744 1974
rect 17584 1538 17744 1946
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _105_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 9128 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _106_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8736 0 -1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _107_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9072 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _108_
timestamp 1698175906
transform -1 0 9632 0 1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _109_
timestamp 1698175906
transform -1 0 8288 0 -1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _110_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10528 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _111_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9240 0 -1 12544
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _112_
timestamp 1698175906
transform 1 0 10584 0 1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _113_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 9912 0 -1 12544
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _114_
timestamp 1698175906
transform -1 0 7952 0 -1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _115_
timestamp 1698175906
transform 1 0 8624 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _116_
timestamp 1698175906
transform -1 0 8232 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _117_
timestamp 1698175906
transform 1 0 8288 0 1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _118_
timestamp 1698175906
transform 1 0 8624 0 1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _119_
timestamp 1698175906
transform 1 0 8904 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _120_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9632 0 1 10192
box -43 -43 883 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _121_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 7504 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _122_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 7616 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _123_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8176 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _124_
timestamp 1698175906
transform 1 0 10976 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _125_
timestamp 1698175906
transform -1 0 12208 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _126_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 8008 0 -1 10192
box -43 -43 771 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _127_
timestamp 1698175906
transform -1 0 8344 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _128_
timestamp 1698175906
transform 1 0 8288 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _129_
timestamp 1698175906
transform 1 0 8960 0 1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _130_
timestamp 1698175906
transform 1 0 9632 0 1 12544
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _131_
timestamp 1698175906
transform 1 0 11424 0 -1 12544
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _132_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 6944 0 1 11760
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _133_
timestamp 1698175906
transform -1 0 6440 0 -1 11760
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _134_
timestamp 1698175906
transform 1 0 12824 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _135_
timestamp 1698175906
transform 1 0 11648 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _136_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9856 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _137_
timestamp 1698175906
transform 1 0 12152 0 -1 10192
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _138_
timestamp 1698175906
transform -1 0 11536 0 -1 9408
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _139_
timestamp 1698175906
transform -1 0 14392 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _140_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 13104 0 1 9408
box -43 -43 715 435
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _141_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10584 0 1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _142_
timestamp 1698175906
transform 1 0 6664 0 1 12544
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _143_
timestamp 1698175906
transform 1 0 7056 0 -1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _144_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9856 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _145_
timestamp 1698175906
transform 1 0 13776 0 1 11760
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _146_
timestamp 1698175906
transform 1 0 12768 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _147_
timestamp 1698175906
transform -1 0 9632 0 -1 13328
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _148_
timestamp 1698175906
transform -1 0 11424 0 -1 14112
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _149_
timestamp 1698175906
transform 1 0 9408 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _150_
timestamp 1698175906
transform 1 0 8904 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _151_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10080 0 1 11760
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _152_
timestamp 1698175906
transform 1 0 10640 0 -1 14112
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _153_
timestamp 1698175906
transform -1 0 9576 0 1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _154_
timestamp 1698175906
transform 1 0 9016 0 1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _155_
timestamp 1698175906
transform 1 0 9352 0 1 11760
box -43 -43 771 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _156_
timestamp 1698175906
transform -1 0 9296 0 1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _157_
timestamp 1698175906
transform -1 0 10248 0 -1 12544
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _158_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9688 0 -1 13328
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _159_
timestamp 1698175906
transform -1 0 9800 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _160_
timestamp 1698175906
transform 1 0 8624 0 -1 13328
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _161_
timestamp 1698175906
transform -1 0 8064 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _162_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 11536 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _163_
timestamp 1698175906
transform 1 0 12824 0 -1 12544
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _164_
timestamp 1698175906
transform -1 0 14000 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _165_
timestamp 1698175906
transform -1 0 12936 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _166_
timestamp 1698175906
transform 1 0 10584 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _167_
timestamp 1698175906
transform -1 0 8904 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _168_
timestamp 1698175906
transform -1 0 11256 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _169_
timestamp 1698175906
transform 1 0 10976 0 -1 9408
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _170_
timestamp 1698175906
transform 1 0 12376 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _171_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 11648 0 1 9408
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _172_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 11704 0 -1 13328
box -43 -43 659 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _173_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 11872 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _174_
timestamp 1698175906
transform -1 0 11704 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _175_
timestamp 1698175906
transform -1 0 9408 0 -1 11760
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _176_
timestamp 1698175906
transform 1 0 9072 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _177_
timestamp 1698175906
transform 1 0 9744 0 -1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _178_
timestamp 1698175906
transform -1 0 7896 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _179_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 7448 0 1 10976
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _180_
timestamp 1698175906
transform -1 0 9800 0 1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _181_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 9744 0 -1 8624
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _182_
timestamp 1698175906
transform 1 0 9240 0 -1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _183_
timestamp 1698175906
transform -1 0 6216 0 1 10192
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _184_
timestamp 1698175906
transform 1 0 6384 0 -1 10192
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _185_
timestamp 1698175906
transform 1 0 11200 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _186_
timestamp 1698175906
transform -1 0 12096 0 -1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _187_
timestamp 1698175906
transform 1 0 11256 0 -1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _188_
timestamp 1698175906
transform -1 0 10976 0 1 7056
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _189_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9296 0 1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _190_
timestamp 1698175906
transform -1 0 7392 0 1 8624
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _191_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 7672 0 1 9408
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _192_
timestamp 1698175906
transform -1 0 7448 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _193_
timestamp 1698175906
transform -1 0 6440 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _194_
timestamp 1698175906
transform -1 0 14056 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _195_
timestamp 1698175906
transform -1 0 12880 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _196_
timestamp 1698175906
transform 1 0 12880 0 -1 9408
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _197_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 12096 0 1 8624
box -43 -43 715 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _198_
timestamp 1698175906
transform 1 0 8680 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _199_
timestamp 1698175906
transform 1 0 10584 0 1 9408
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _200_
timestamp 1698175906
transform 1 0 10416 0 -1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _201_
timestamp 1698175906
transform -1 0 11256 0 1 8624
box -43 -43 715 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _202_
timestamp 1698175906
transform -1 0 13216 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _203_
timestamp 1698175906
transform 1 0 11200 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _204_
timestamp 1698175906
transform 1 0 12544 0 -1 8624
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _205_
timestamp 1698175906
transform -1 0 12992 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _206_
timestamp 1698175906
transform 1 0 11648 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _207_
timestamp 1698175906
transform 1 0 12544 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _208_
timestamp 1698175906
transform -1 0 14672 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _209_
timestamp 1698175906
transform 1 0 12544 0 -1 10192
box -43 -43 715 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _210_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 13160 0 1 11760
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _211_
timestamp 1698175906
transform 1 0 7168 0 1 11760
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _212_
timestamp 1698175906
transform 1 0 6888 0 -1 8624
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _213_
timestamp 1698175906
transform 1 0 6664 0 1 10192
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _214_
timestamp 1698175906
transform -1 0 6496 0 1 11760
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _215_
timestamp 1698175906
transform 1 0 13272 0 -1 9408
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _216_
timestamp 1698175906
transform -1 0 7056 0 -1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _217_
timestamp 1698175906
transform 1 0 13216 0 -1 11760
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _218_
timestamp 1698175906
transform 1 0 10584 0 1 14112
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _219_
timestamp 1698175906
transform 1 0 8008 0 1 14112
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _220_
timestamp 1698175906
transform 1 0 8792 0 -1 14112
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _221_
timestamp 1698175906
transform 1 0 6944 0 1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _222_
timestamp 1698175906
transform 1 0 13328 0 -1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _223_
timestamp 1698175906
transform 1 0 11704 0 1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _224_
timestamp 1698175906
transform 1 0 11256 0 1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _225_
timestamp 1698175906
transform -1 0 7224 0 -1 10976
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _226_
timestamp 1698175906
transform 1 0 8232 0 1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _227_
timestamp 1698175906
transform -1 0 6384 0 -1 10192
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _228_
timestamp 1698175906
transform 1 0 9744 0 -1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _229_
timestamp 1698175906
transform -1 0 7000 0 -1 9408
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _230_
timestamp 1698175906
transform 1 0 12768 0 1 8624
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _231_
timestamp 1698175906
transform -1 0 11256 0 -1 7840
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _232_
timestamp 1698175906
transform 1 0 11872 0 1 7840
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _233_
timestamp 1698175906
transform 1 0 11760 0 1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _234_
timestamp 1698175906
transform 1 0 13384 0 -1 10192
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _238_
timestamp 1698175906
transform -1 0 7112 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _239_
timestamp 1698175906
transform 1 0 14504 0 1 12544
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__132__A2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 7056 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__142__A2
timestamp 1698175906
transform -1 0 7168 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__183__A2
timestamp 1698175906
transform 1 0 6328 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__209__A2
timestamp 1698175906
transform 1 0 12656 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__210__CLK
timestamp 1698175906
transform 1 0 13272 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__211__CLK
timestamp 1698175906
transform 1 0 8904 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__212__CLK
timestamp 1698175906
transform 1 0 8736 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__213__CLK
timestamp 1698175906
transform 1 0 8344 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__214__CLK
timestamp 1698175906
transform 1 0 6496 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__215__CLK
timestamp 1698175906
transform 1 0 12320 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__216__CLK
timestamp 1698175906
transform 1 0 7448 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__217__CLK
timestamp 1698175906
transform 1 0 12656 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__218__CLK
timestamp 1698175906
transform 1 0 12320 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__219__CLK
timestamp 1698175906
transform 1 0 9744 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__220__CLK
timestamp 1698175906
transform 1 0 8400 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__221__CLK
timestamp 1698175906
transform 1 0 8680 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__222__CLK
timestamp 1698175906
transform 1 0 13216 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__223__CLK
timestamp 1698175906
transform 1 0 13440 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__224__CLK
timestamp 1698175906
transform 1 0 12992 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__225__CLK
timestamp 1698175906
transform 1 0 7336 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__226__CLK
timestamp 1698175906
transform 1 0 9968 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__227__CLK
timestamp 1698175906
transform 1 0 6776 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__228__CLK
timestamp 1698175906
transform 1 0 11480 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__229__CLK
timestamp 1698175906
transform 1 0 7000 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__230__CLK
timestamp 1698175906
transform 1 0 14616 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__231__CLK
timestamp 1698175906
transform 1 0 11704 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__232__CLK
timestamp 1698175906
transform 1 0 13608 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__233__CLK
timestamp 1698175906
transform 1 0 13496 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__234__CLK
timestamp 1698175906
transform 1 0 13272 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1698175906
transform 1 0 10696 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9520 0 -1 10976
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1698175906
transform -1 0 10472 0 1 10976
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1698175906
transform 1 0 11256 0 1 10192
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 784 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698175906
transform 1 0 2688 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698175906
transform 1 0 4592 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698175906
transform 1 0 6496 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_138 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8400 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_146 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8848 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_150 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9072 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_155
timestamp 1698175906
transform 1 0 9352 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_163
timestamp 1698175906
transform 1 0 9800 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_167 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10024 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_169
timestamp 1698175906
transform 1 0 10136 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_172
timestamp 1698175906
transform 1 0 10304 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_176
timestamp 1698175906
transform 1 0 10528 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_206
timestamp 1698175906
transform 1 0 12208 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_240
timestamp 1698175906
transform 1 0 14112 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_274
timestamp 1698175906
transform 1 0 16016 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_308
timestamp 1698175906
transform 1 0 17920 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_342
timestamp 1698175906
transform 1 0 19824 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_346
timestamp 1698175906
transform 1 0 20048 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_348
timestamp 1698175906
transform 1 0 20160 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 784 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698175906
transform 1 0 4368 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698175906
transform 1 0 4704 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698175906
transform 1 0 8288 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_142
timestamp 1698175906
transform 1 0 8624 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_150
timestamp 1698175906
transform 1 0 9072 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_154
timestamp 1698175906
transform 1 0 9296 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_207
timestamp 1698175906
transform 1 0 12264 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_209
timestamp 1698175906
transform 1 0 12376 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_212
timestamp 1698175906
transform 1 0 12544 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_220
timestamp 1698175906
transform 1 0 12992 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_222
timestamp 1698175906
transform 1 0 13104 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_249 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 14616 0 -1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_265
timestamp 1698175906
transform 1 0 15512 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_273
timestamp 1698175906
transform 1 0 15960 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_277
timestamp 1698175906
transform 1 0 16184 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_279
timestamp 1698175906
transform 1 0 16296 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_282
timestamp 1698175906
transform 1 0 16464 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_346
timestamp 1698175906
transform 1 0 20048 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_348
timestamp 1698175906
transform 1 0 20160 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698175906
transform 1 0 784 0 1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698175906
transform 1 0 2576 0 1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698175906
transform 1 0 2744 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698175906
transform 1 0 6328 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_107
timestamp 1698175906
transform 1 0 6664 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_171
timestamp 1698175906
transform 1 0 10248 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_177
timestamp 1698175906
transform 1 0 10584 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_241
timestamp 1698175906
transform 1 0 14168 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698175906
transform 1 0 14504 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698175906
transform 1 0 18088 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_317
timestamp 1698175906
transform 1 0 18424 0 1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698175906
transform 1 0 784 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698175906
transform 1 0 4368 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698175906
transform 1 0 4704 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698175906
transform 1 0 8288 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_142
timestamp 1698175906
transform 1 0 8624 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_206
timestamp 1698175906
transform 1 0 12208 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_212
timestamp 1698175906
transform 1 0 12544 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_276
timestamp 1698175906
transform 1 0 16128 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_282
timestamp 1698175906
transform 1 0 16464 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_346
timestamp 1698175906
transform 1 0 20048 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_348
timestamp 1698175906
transform 1 0 20160 0 -1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698175906
transform 1 0 784 0 1 3136
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698175906
transform 1 0 2576 0 1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698175906
transform 1 0 2744 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698175906
transform 1 0 6328 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_107
timestamp 1698175906
transform 1 0 6664 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698175906
transform 1 0 10248 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_177
timestamp 1698175906
transform 1 0 10584 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_241
timestamp 1698175906
transform 1 0 14168 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698175906
transform 1 0 14504 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698175906
transform 1 0 18088 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_317
timestamp 1698175906
transform 1 0 18424 0 1 3136
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698175906
transform 1 0 784 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698175906
transform 1 0 4368 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698175906
transform 1 0 4704 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698175906
transform 1 0 8288 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_142
timestamp 1698175906
transform 1 0 8624 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_206
timestamp 1698175906
transform 1 0 12208 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_212
timestamp 1698175906
transform 1 0 12544 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698175906
transform 1 0 16128 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_282
timestamp 1698175906
transform 1 0 16464 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_346
timestamp 1698175906
transform 1 0 20048 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_348
timestamp 1698175906
transform 1 0 20160 0 -1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698175906
transform 1 0 784 0 1 3920
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698175906
transform 1 0 2576 0 1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698175906
transform 1 0 2744 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698175906
transform 1 0 6328 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_107
timestamp 1698175906
transform 1 0 6664 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_171
timestamp 1698175906
transform 1 0 10248 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_177
timestamp 1698175906
transform 1 0 10584 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_241
timestamp 1698175906
transform 1 0 14168 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_247
timestamp 1698175906
transform 1 0 14504 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_311
timestamp 1698175906
transform 1 0 18088 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_317
timestamp 1698175906
transform 1 0 18424 0 1 3920
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698175906
transform 1 0 784 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698175906
transform 1 0 4368 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_72
timestamp 1698175906
transform 1 0 4704 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698175906
transform 1 0 8288 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_142
timestamp 1698175906
transform 1 0 8624 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_206
timestamp 1698175906
transform 1 0 12208 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_212
timestamp 1698175906
transform 1 0 12544 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_276
timestamp 1698175906
transform 1 0 16128 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_282
timestamp 1698175906
transform 1 0 16464 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_346
timestamp 1698175906
transform 1 0 20048 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_348
timestamp 1698175906
transform 1 0 20160 0 -1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698175906
transform 1 0 784 0 1 4704
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698175906
transform 1 0 2576 0 1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_37
timestamp 1698175906
transform 1 0 2744 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_101
timestamp 1698175906
transform 1 0 6328 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_107
timestamp 1698175906
transform 1 0 6664 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_171
timestamp 1698175906
transform 1 0 10248 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_177
timestamp 1698175906
transform 1 0 10584 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_241
timestamp 1698175906
transform 1 0 14168 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_247
timestamp 1698175906
transform 1 0 14504 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_311
timestamp 1698175906
transform 1 0 18088 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_317
timestamp 1698175906
transform 1 0 18424 0 1 4704
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698175906
transform 1 0 784 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698175906
transform 1 0 4368 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_72
timestamp 1698175906
transform 1 0 4704 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_136
timestamp 1698175906
transform 1 0 8288 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_142
timestamp 1698175906
transform 1 0 8624 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_206
timestamp 1698175906
transform 1 0 12208 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_212
timestamp 1698175906
transform 1 0 12544 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_276
timestamp 1698175906
transform 1 0 16128 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_282
timestamp 1698175906
transform 1 0 16464 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_346
timestamp 1698175906
transform 1 0 20048 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_348
timestamp 1698175906
transform 1 0 20160 0 -1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698175906
transform 1 0 784 0 1 5488
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698175906
transform 1 0 2576 0 1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_37
timestamp 1698175906
transform 1 0 2744 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698175906
transform 1 0 6328 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_107
timestamp 1698175906
transform 1 0 6664 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_171
timestamp 1698175906
transform 1 0 10248 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_177
timestamp 1698175906
transform 1 0 10584 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_241
timestamp 1698175906
transform 1 0 14168 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_247
timestamp 1698175906
transform 1 0 14504 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_311
timestamp 1698175906
transform 1 0 18088 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_317
timestamp 1698175906
transform 1 0 18424 0 1 5488
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2
timestamp 1698175906
transform 1 0 784 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698175906
transform 1 0 4368 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_72
timestamp 1698175906
transform 1 0 4704 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698175906
transform 1 0 8288 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_142
timestamp 1698175906
transform 1 0 8624 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_206
timestamp 1698175906
transform 1 0 12208 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_212
timestamp 1698175906
transform 1 0 12544 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_276
timestamp 1698175906
transform 1 0 16128 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_282
timestamp 1698175906
transform 1 0 16464 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_346
timestamp 1698175906
transform 1 0 20048 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_348
timestamp 1698175906
transform 1 0 20160 0 -1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698175906
transform 1 0 784 0 1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698175906
transform 1 0 2576 0 1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_37
timestamp 1698175906
transform 1 0 2744 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698175906
transform 1 0 6328 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_107
timestamp 1698175906
transform 1 0 6664 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_171
timestamp 1698175906
transform 1 0 10248 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_177
timestamp 1698175906
transform 1 0 10584 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_241
timestamp 1698175906
transform 1 0 14168 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_247
timestamp 1698175906
transform 1 0 14504 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_311
timestamp 1698175906
transform 1 0 18088 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_317
timestamp 1698175906
transform 1 0 18424 0 1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_2
timestamp 1698175906
transform 1 0 784 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_66
timestamp 1698175906
transform 1 0 4368 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_72
timestamp 1698175906
transform 1 0 4704 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_136
timestamp 1698175906
transform 1 0 8288 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_142
timestamp 1698175906
transform 1 0 8624 0 -1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_158
timestamp 1698175906
transform 1 0 9520 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_191
timestamp 1698175906
transform 1 0 11368 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_195
timestamp 1698175906
transform 1 0 11592 0 -1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_203
timestamp 1698175906
transform 1 0 12040 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_207
timestamp 1698175906
transform 1 0 12264 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_209
timestamp 1698175906
transform 1 0 12376 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_212
timestamp 1698175906
transform 1 0 12544 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_220
timestamp 1698175906
transform 1 0 12992 0 -1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_252
timestamp 1698175906
transform 1 0 14784 0 -1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_268
timestamp 1698175906
transform 1 0 15680 0 -1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_276
timestamp 1698175906
transform 1 0 16128 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_282
timestamp 1698175906
transform 1 0 16464 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_346
timestamp 1698175906
transform 1 0 20048 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_348
timestamp 1698175906
transform 1 0 20160 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698175906
transform 1 0 784 0 1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698175906
transform 1 0 2576 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_37
timestamp 1698175906
transform 1 0 2744 0 1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_101
timestamp 1698175906
transform 1 0 6328 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_107
timestamp 1698175906
transform 1 0 6664 0 1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_123
timestamp 1698175906
transform 1 0 7560 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_131
timestamp 1698175906
transform 1 0 8008 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_164
timestamp 1698175906
transform 1 0 9856 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_168
timestamp 1698175906
transform 1 0 10080 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_172
timestamp 1698175906
transform 1 0 10304 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_174
timestamp 1698175906
transform 1 0 10416 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_177
timestamp 1698175906
transform 1 0 10584 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_184
timestamp 1698175906
transform 1 0 10976 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_192
timestamp 1698175906
transform 1 0 11424 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_196
timestamp 1698175906
transform 1 0 11648 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_227
timestamp 1698175906
transform 1 0 13384 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_231
timestamp 1698175906
transform 1 0 13608 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_239
timestamp 1698175906
transform 1 0 14056 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_243
timestamp 1698175906
transform 1 0 14280 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_247
timestamp 1698175906
transform 1 0 14504 0 1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_311
timestamp 1698175906
transform 1 0 18088 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_317
timestamp 1698175906
transform 1 0 18424 0 1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_2
timestamp 1698175906
transform 1 0 784 0 -1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_66
timestamp 1698175906
transform 1 0 4368 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_72
timestamp 1698175906
transform 1 0 4704 0 -1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_136
timestamp 1698175906
transform 1 0 8288 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_142
timestamp 1698175906
transform 1 0 8624 0 -1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_158
timestamp 1698175906
transform 1 0 9520 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_195
timestamp 1698175906
transform 1 0 11592 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_199
timestamp 1698175906
transform 1 0 11816 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_207
timestamp 1698175906
transform 1 0 12264 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_209
timestamp 1698175906
transform 1 0 12376 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_224
timestamp 1698175906
transform 1 0 13216 0 -1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_256
timestamp 1698175906
transform 1 0 15008 0 -1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_272
timestamp 1698175906
transform 1 0 15904 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_282
timestamp 1698175906
transform 1 0 16464 0 -1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_346
timestamp 1698175906
transform 1 0 20048 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_348
timestamp 1698175906
transform 1 0 20160 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_2
timestamp 1698175906
transform 1 0 784 0 1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698175906
transform 1 0 2576 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_37
timestamp 1698175906
transform 1 0 2744 0 1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_101
timestamp 1698175906
transform 1 0 6328 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_107
timestamp 1698175906
transform 1 0 6664 0 1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_139
timestamp 1698175906
transform 1 0 8456 0 1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_155
timestamp 1698175906
transform 1 0 9352 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_163
timestamp 1698175906
transform 1 0 9800 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_171
timestamp 1698175906
transform 1 0 10248 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_177
timestamp 1698175906
transform 1 0 10584 0 1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_193
timestamp 1698175906
transform 1 0 11480 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_197
timestamp 1698175906
transform 1 0 11704 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_199
timestamp 1698175906
transform 1 0 11816 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_229
timestamp 1698175906
transform 1 0 13496 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_233
timestamp 1698175906
transform 1 0 13720 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_241
timestamp 1698175906
transform 1 0 14168 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_247
timestamp 1698175906
transform 1 0 14504 0 1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_311
timestamp 1698175906
transform 1 0 18088 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_317
timestamp 1698175906
transform 1 0 18424 0 1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_2
timestamp 1698175906
transform 1 0 784 0 -1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_66
timestamp 1698175906
transform 1 0 4368 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_72
timestamp 1698175906
transform 1 0 4704 0 -1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_104
timestamp 1698175906
transform 1 0 6496 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_108
timestamp 1698175906
transform 1 0 6720 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_110
timestamp 1698175906
transform 1 0 6832 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_142
timestamp 1698175906
transform 1 0 8624 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_146
timestamp 1698175906
transform 1 0 8848 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_150
timestamp 1698175906
transform 1 0 9072 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_168
timestamp 1698175906
transform 1 0 10080 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_172
timestamp 1698175906
transform 1 0 10304 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_180
timestamp 1698175906
transform 1 0 10752 0 -1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_196
timestamp 1698175906
transform 1 0 11648 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_204
timestamp 1698175906
transform 1 0 12096 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_208
timestamp 1698175906
transform 1 0 12320 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_222
timestamp 1698175906
transform 1 0 13104 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_230
timestamp 1698175906
transform 1 0 13552 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_234
timestamp 1698175906
transform 1 0 13776 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_239
timestamp 1698175906
transform 1 0 14056 0 -1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_271
timestamp 1698175906
transform 1 0 15848 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_279
timestamp 1698175906
transform 1 0 16296 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_282
timestamp 1698175906
transform 1 0 16464 0 -1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_314
timestamp 1698175906
transform 1 0 18256 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_322
timestamp 1698175906
transform 1 0 18704 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_28
timestamp 1698175906
transform 1 0 2240 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_32
timestamp 1698175906
transform 1 0 2464 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698175906
transform 1 0 2576 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_37
timestamp 1698175906
transform 1 0 2744 0 1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_69
timestamp 1698175906
transform 1 0 4536 0 1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_85
timestamp 1698175906
transform 1 0 5432 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_93
timestamp 1698175906
transform 1 0 5880 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_103
timestamp 1698175906
transform 1 0 6440 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_107
timestamp 1698175906
transform 1 0 6664 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_124
timestamp 1698175906
transform 1 0 7616 0 1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_156
timestamp 1698175906
transform 1 0 9408 0 1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_172
timestamp 1698175906
transform 1 0 10304 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_174
timestamp 1698175906
transform 1 0 10416 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_189
timestamp 1698175906
transform 1 0 11256 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_193
timestamp 1698175906
transform 1 0 11480 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_195
timestamp 1698175906
transform 1 0 11592 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_247
timestamp 1698175906
transform 1 0 14504 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_251
timestamp 1698175906
transform 1 0 14728 0 1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_317
timestamp 1698175906
transform 1 0 18424 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_321
timestamp 1698175906
transform 1 0 18648 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_28
timestamp 1698175906
transform 1 0 2240 0 -1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_60
timestamp 1698175906
transform 1 0 4032 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_68
timestamp 1698175906
transform 1 0 4480 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_72
timestamp 1698175906
transform 1 0 4704 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_80
timestamp 1698175906
transform 1 0 5152 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_121
timestamp 1698175906
transform 1 0 7448 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_130
timestamp 1698175906
transform 1 0 7952 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_134
timestamp 1698175906
transform 1 0 8176 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_148
timestamp 1698175906
transform 1 0 8960 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_158
timestamp 1698175906
transform 1 0 9520 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_162
timestamp 1698175906
transform 1 0 9744 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_172
timestamp 1698175906
transform 1 0 10304 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_180
timestamp 1698175906
transform 1 0 10752 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_194
timestamp 1698175906
transform 1 0 11536 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_198
timestamp 1698175906
transform 1 0 11760 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_206
timestamp 1698175906
transform 1 0 12208 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_223
timestamp 1698175906
transform 1 0 13160 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_254
timestamp 1698175906
transform 1 0 14896 0 -1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_270
timestamp 1698175906
transform 1 0 15792 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_278
timestamp 1698175906
transform 1 0 16240 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_282
timestamp 1698175906
transform 1 0 16464 0 -1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_346
timestamp 1698175906
transform 1 0 20048 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_348
timestamp 1698175906
transform 1 0 20160 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_2
timestamp 1698175906
transform 1 0 784 0 1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698175906
transform 1 0 2576 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_37
timestamp 1698175906
transform 1 0 2744 0 1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_101
timestamp 1698175906
transform 1 0 6328 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_107
timestamp 1698175906
transform 1 0 6664 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_111
timestamp 1698175906
transform 1 0 6888 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_125
timestamp 1698175906
transform 1 0 7672 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_135
timestamp 1698175906
transform 1 0 8232 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_139
timestamp 1698175906
transform 1 0 8456 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_153
timestamp 1698175906
transform 1 0 9240 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_170
timestamp 1698175906
transform 1 0 10192 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_174
timestamp 1698175906
transform 1 0 10416 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_184
timestamp 1698175906
transform 1 0 10976 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_234
timestamp 1698175906
transform 1 0 13776 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_238
timestamp 1698175906
transform 1 0 14000 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_240
timestamp 1698175906
transform 1 0 14112 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_247
timestamp 1698175906
transform 1 0 14504 0 1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_311
timestamp 1698175906
transform 1 0 18088 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_317
timestamp 1698175906
transform 1 0 18424 0 1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_2
timestamp 1698175906
transform 1 0 784 0 -1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_66
timestamp 1698175906
transform 1 0 4368 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_72
timestamp 1698175906
transform 1 0 4704 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_107
timestamp 1698175906
transform 1 0 6664 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_111
timestamp 1698175906
transform 1 0 6888 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_115
timestamp 1698175906
transform 1 0 7112 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_117
timestamp 1698175906
transform 1 0 7224 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_131
timestamp 1698175906
transform 1 0 8008 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_133
timestamp 1698175906
transform 1 0 8120 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_142
timestamp 1698175906
transform 1 0 8624 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_185
timestamp 1698175906
transform 1 0 11032 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_187
timestamp 1698175906
transform 1 0 11144 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_202
timestamp 1698175906
transform 1 0 11984 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_204
timestamp 1698175906
transform 1 0 12096 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_224
timestamp 1698175906
transform 1 0 13216 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_226
timestamp 1698175906
transform 1 0 13328 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_256
timestamp 1698175906
transform 1 0 15008 0 -1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_272
timestamp 1698175906
transform 1 0 15904 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_282
timestamp 1698175906
transform 1 0 16464 0 -1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_314
timestamp 1698175906
transform 1 0 18256 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_322
timestamp 1698175906
transform 1 0 18704 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_2
timestamp 1698175906
transform 1 0 784 0 1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698175906
transform 1 0 2576 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_37
timestamp 1698175906
transform 1 0 2744 0 1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_69
timestamp 1698175906
transform 1 0 4536 0 1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_85
timestamp 1698175906
transform 1 0 5432 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_93
timestamp 1698175906
transform 1 0 5880 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_99
timestamp 1698175906
transform 1 0 6216 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_103
timestamp 1698175906
transform 1 0 6440 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_177
timestamp 1698175906
transform 1 0 10584 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_239
timestamp 1698175906
transform 1 0 14056 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_243
timestamp 1698175906
transform 1 0 14280 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_247
timestamp 1698175906
transform 1 0 14504 0 1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_311
timestamp 1698175906
transform 1 0 18088 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_317
timestamp 1698175906
transform 1 0 18424 0 1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_333
timestamp 1698175906
transform 1 0 19320 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_341
timestamp 1698175906
transform 1 0 19768 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_28
timestamp 1698175906
transform 1 0 2240 0 -1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_60
timestamp 1698175906
transform 1 0 4032 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_68
timestamp 1698175906
transform 1 0 4480 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_72
timestamp 1698175906
transform 1 0 4704 0 -1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_117
timestamp 1698175906
transform 1 0 7224 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_137
timestamp 1698175906
transform 1 0 8344 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_139
timestamp 1698175906
transform 1 0 8456 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_142
timestamp 1698175906
transform 1 0 8624 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_208
timestamp 1698175906
transform 1 0 12320 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_212
timestamp 1698175906
transform 1 0 12544 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_216
timestamp 1698175906
transform 1 0 12768 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_224
timestamp 1698175906
transform 1 0 13216 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_227
timestamp 1698175906
transform 1 0 13384 0 -1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_243
timestamp 1698175906
transform 1 0 14280 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_245
timestamp 1698175906
transform 1 0 14392 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_250
timestamp 1698175906
transform 1 0 14672 0 -1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_266
timestamp 1698175906
transform 1 0 15568 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_274
timestamp 1698175906
transform 1 0 16016 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_278
timestamp 1698175906
transform 1 0 16240 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_282
timestamp 1698175906
transform 1 0 16464 0 -1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_314
timestamp 1698175906
transform 1 0 18256 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_322
timestamp 1698175906
transform 1 0 18704 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_28
timestamp 1698175906
transform 1 0 2240 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_32
timestamp 1698175906
transform 1 0 2464 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698175906
transform 1 0 2576 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_37
timestamp 1698175906
transform 1 0 2744 0 1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_101
timestamp 1698175906
transform 1 0 6328 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_107
timestamp 1698175906
transform 1 0 6664 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_111
timestamp 1698175906
transform 1 0 6888 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_121
timestamp 1698175906
transform 1 0 7448 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_223
timestamp 1698175906
transform 1 0 13160 0 1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_239
timestamp 1698175906
transform 1 0 14056 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_243
timestamp 1698175906
transform 1 0 14280 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_247
timestamp 1698175906
transform 1 0 14504 0 1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_311
timestamp 1698175906
transform 1 0 18088 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_317
timestamp 1698175906
transform 1 0 18424 0 1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_2
timestamp 1698175906
transform 1 0 784 0 -1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_66
timestamp 1698175906
transform 1 0 4368 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_72
timestamp 1698175906
transform 1 0 4704 0 -1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_88
timestamp 1698175906
transform 1 0 5600 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_96
timestamp 1698175906
transform 1 0 6048 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_103
timestamp 1698175906
transform 1 0 6440 0 -1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_119
timestamp 1698175906
transform 1 0 7336 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_123
timestamp 1698175906
transform 1 0 7560 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_136
timestamp 1698175906
transform 1 0 8288 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_142
timestamp 1698175906
transform 1 0 8624 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_146
timestamp 1698175906
transform 1 0 8848 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_172
timestamp 1698175906
transform 1 0 10304 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_192
timestamp 1698175906
transform 1 0 11424 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_202
timestamp 1698175906
transform 1 0 11984 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_212
timestamp 1698175906
transform 1 0 12544 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_253
timestamp 1698175906
transform 1 0 14840 0 -1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_269
timestamp 1698175906
transform 1 0 15736 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_277
timestamp 1698175906
transform 1 0 16184 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_279
timestamp 1698175906
transform 1 0 16296 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_282
timestamp 1698175906
transform 1 0 16464 0 -1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_346
timestamp 1698175906
transform 1 0 20048 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_348
timestamp 1698175906
transform 1 0 20160 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_28
timestamp 1698175906
transform 1 0 2240 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_32
timestamp 1698175906
transform 1 0 2464 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698175906
transform 1 0 2576 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_37
timestamp 1698175906
transform 1 0 2744 0 1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_69
timestamp 1698175906
transform 1 0 4536 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_73
timestamp 1698175906
transform 1 0 4760 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_104
timestamp 1698175906
transform 1 0 6496 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_112
timestamp 1698175906
transform 1 0 6944 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_145
timestamp 1698175906
transform 1 0 8792 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_183
timestamp 1698175906
transform 1 0 10920 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_191
timestamp 1698175906
transform 1 0 11368 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_193
timestamp 1698175906
transform 1 0 11480 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_223
timestamp 1698175906
transform 1 0 13160 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_227
timestamp 1698175906
transform 1 0 13384 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_231
timestamp 1698175906
transform 1 0 13608 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_233
timestamp 1698175906
transform 1 0 13720 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_239
timestamp 1698175906
transform 1 0 14056 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_243
timestamp 1698175906
transform 1 0 14280 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_247
timestamp 1698175906
transform 1 0 14504 0 1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_311
timestamp 1698175906
transform 1 0 18088 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_317
timestamp 1698175906
transform 1 0 18424 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_321
timestamp 1698175906
transform 1 0 18648 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_2
timestamp 1698175906
transform 1 0 784 0 -1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_66
timestamp 1698175906
transform 1 0 4368 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_72
timestamp 1698175906
transform 1 0 4704 0 -1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_106
timestamp 1698175906
transform 1 0 6608 0 -1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_138
timestamp 1698175906
transform 1 0 8400 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_142
timestamp 1698175906
transform 1 0 8624 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_150
timestamp 1698175906
transform 1 0 9072 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_152
timestamp 1698175906
transform 1 0 9184 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_171
timestamp 1698175906
transform 1 0 10248 0 -1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_187
timestamp 1698175906
transform 1 0 11144 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_191
timestamp 1698175906
transform 1 0 11368 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_198
timestamp 1698175906
transform 1 0 11760 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_208
timestamp 1698175906
transform 1 0 12320 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_212
timestamp 1698175906
transform 1 0 12544 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_216
timestamp 1698175906
transform 1 0 12768 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_255
timestamp 1698175906
transform 1 0 14952 0 -1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_271
timestamp 1698175906
transform 1 0 15848 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_279
timestamp 1698175906
transform 1 0 16296 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_282
timestamp 1698175906
transform 1 0 16464 0 -1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_346
timestamp 1698175906
transform 1 0 20048 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_348
timestamp 1698175906
transform 1 0 20160 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_2
timestamp 1698175906
transform 1 0 784 0 1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698175906
transform 1 0 2576 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_37
timestamp 1698175906
transform 1 0 2744 0 1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_101
timestamp 1698175906
transform 1 0 6328 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_112
timestamp 1698175906
transform 1 0 6944 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_116
timestamp 1698175906
transform 1 0 7168 0 1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_148
timestamp 1698175906
transform 1 0 8960 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_156
timestamp 1698175906
transform 1 0 9408 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_166
timestamp 1698175906
transform 1 0 9968 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_174
timestamp 1698175906
transform 1 0 10416 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_185
timestamp 1698175906
transform 1 0 11032 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_218
timestamp 1698175906
transform 1 0 12880 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_222
timestamp 1698175906
transform 1 0 13104 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_226
timestamp 1698175906
transform 1 0 13328 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_238
timestamp 1698175906
transform 1 0 14000 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_242
timestamp 1698175906
transform 1 0 14224 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_244
timestamp 1698175906
transform 1 0 14336 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_253
timestamp 1698175906
transform 1 0 14840 0 1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_285
timestamp 1698175906
transform 1 0 16632 0 1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_301
timestamp 1698175906
transform 1 0 17528 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_309
timestamp 1698175906
transform 1 0 17976 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_313
timestamp 1698175906
transform 1 0 18200 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_317
timestamp 1698175906
transform 1 0 18424 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_321
timestamp 1698175906
transform 1 0 18648 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_28
timestamp 1698175906
transform 1 0 2240 0 -1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_60
timestamp 1698175906
transform 1 0 4032 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_68
timestamp 1698175906
transform 1 0 4480 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_72
timestamp 1698175906
transform 1 0 4704 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_80
timestamp 1698175906
transform 1 0 5152 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_84
timestamp 1698175906
transform 1 0 5376 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_119
timestamp 1698175906
transform 1 0 7336 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_123
timestamp 1698175906
transform 1 0 7560 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_127
timestamp 1698175906
transform 1 0 7784 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_132
timestamp 1698175906
transform 1 0 8064 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_151
timestamp 1698175906
transform 1 0 9128 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_153
timestamp 1698175906
transform 1 0 9240 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_160
timestamp 1698175906
transform 1 0 9632 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_170
timestamp 1698175906
transform 1 0 10192 0 -1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_186
timestamp 1698175906
transform 1 0 11088 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_188
timestamp 1698175906
transform 1 0 11200 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_208
timestamp 1698175906
transform 1 0 12320 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_212
timestamp 1698175906
transform 1 0 12544 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_214
timestamp 1698175906
transform 1 0 12656 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_219
timestamp 1698175906
transform 1 0 12936 0 -1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_251
timestamp 1698175906
transform 1 0 14728 0 -1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_267
timestamp 1698175906
transform 1 0 15624 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_275
timestamp 1698175906
transform 1 0 16072 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_279
timestamp 1698175906
transform 1 0 16296 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_282
timestamp 1698175906
transform 1 0 16464 0 -1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_314
timestamp 1698175906
transform 1 0 18256 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_322
timestamp 1698175906
transform 1 0 18704 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_2
timestamp 1698175906
transform 1 0 784 0 1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698175906
transform 1 0 2576 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_37
timestamp 1698175906
transform 1 0 2744 0 1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_101
timestamp 1698175906
transform 1 0 6328 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_107
timestamp 1698175906
transform 1 0 6664 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_111
timestamp 1698175906
transform 1 0 6888 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_141
timestamp 1698175906
transform 1 0 8568 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_145
timestamp 1698175906
transform 1 0 8792 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_163
timestamp 1698175906
transform 1 0 9800 0 1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_171
timestamp 1698175906
transform 1 0 10248 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_177
timestamp 1698175906
transform 1 0 10584 0 1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_193
timestamp 1698175906
transform 1 0 11480 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_226
timestamp 1698175906
transform 1 0 13328 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_230
timestamp 1698175906
transform 1 0 13552 0 1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_238
timestamp 1698175906
transform 1 0 14000 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_242
timestamp 1698175906
transform 1 0 14224 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_244
timestamp 1698175906
transform 1 0 14336 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_247
timestamp 1698175906
transform 1 0 14504 0 1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_311
timestamp 1698175906
transform 1 0 18088 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_317
timestamp 1698175906
transform 1 0 18424 0 1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_2
timestamp 1698175906
transform 1 0 784 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_66
timestamp 1698175906
transform 1 0 4368 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_72
timestamp 1698175906
transform 1 0 4704 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_136
timestamp 1698175906
transform 1 0 8288 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_142
timestamp 1698175906
transform 1 0 8624 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_144
timestamp 1698175906
transform 1 0 8736 0 -1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_174
timestamp 1698175906
transform 1 0 10416 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_183
timestamp 1698175906
transform 1 0 10920 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_192
timestamp 1698175906
transform 1 0 11424 0 -1 14112
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_208
timestamp 1698175906
transform 1 0 12320 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_212
timestamp 1698175906
transform 1 0 12544 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_276
timestamp 1698175906
transform 1 0 16128 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_282
timestamp 1698175906
transform 1 0 16464 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_346
timestamp 1698175906
transform 1 0 20048 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_348
timestamp 1698175906
transform 1 0 20160 0 -1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_2
timestamp 1698175906
transform 1 0 784 0 1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698175906
transform 1 0 2576 0 1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_37
timestamp 1698175906
transform 1 0 2744 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_101
timestamp 1698175906
transform 1 0 6328 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_107
timestamp 1698175906
transform 1 0 6664 0 1 14112
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_123
timestamp 1698175906
transform 1 0 7560 0 1 14112
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_160
timestamp 1698175906
transform 1 0 9632 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_164
timestamp 1698175906
transform 1 0 9856 0 1 14112
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_172
timestamp 1698175906
transform 1 0 10304 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_174
timestamp 1698175906
transform 1 0 10416 0 1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_206
timestamp 1698175906
transform 1 0 12208 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_210
timestamp 1698175906
transform 1 0 12432 0 1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_242
timestamp 1698175906
transform 1 0 14224 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_244
timestamp 1698175906
transform 1 0 14336 0 1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_247
timestamp 1698175906
transform 1 0 14504 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_311
timestamp 1698175906
transform 1 0 18088 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_317
timestamp 1698175906
transform 1 0 18424 0 1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_2
timestamp 1698175906
transform 1 0 784 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_66
timestamp 1698175906
transform 1 0 4368 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_72
timestamp 1698175906
transform 1 0 4704 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_136
timestamp 1698175906
transform 1 0 8288 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_142
timestamp 1698175906
transform 1 0 8624 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_206
timestamp 1698175906
transform 1 0 12208 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_212
timestamp 1698175906
transform 1 0 12544 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_276
timestamp 1698175906
transform 1 0 16128 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_282
timestamp 1698175906
transform 1 0 16464 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_346
timestamp 1698175906
transform 1 0 20048 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_348
timestamp 1698175906
transform 1 0 20160 0 -1 14896
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698175906
transform 1 0 784 0 1 14896
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698175906
transform 1 0 2576 0 1 14896
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_37
timestamp 1698175906
transform 1 0 2744 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_101
timestamp 1698175906
transform 1 0 6328 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_107
timestamp 1698175906
transform 1 0 6664 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_171
timestamp 1698175906
transform 1 0 10248 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_177
timestamp 1698175906
transform 1 0 10584 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_241
timestamp 1698175906
transform 1 0 14168 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_247
timestamp 1698175906
transform 1 0 14504 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_311
timestamp 1698175906
transform 1 0 18088 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_317
timestamp 1698175906
transform 1 0 18424 0 1 14896
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2
timestamp 1698175906
transform 1 0 784 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_66
timestamp 1698175906
transform 1 0 4368 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_72
timestamp 1698175906
transform 1 0 4704 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_136
timestamp 1698175906
transform 1 0 8288 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_142
timestamp 1698175906
transform 1 0 8624 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_206
timestamp 1698175906
transform 1 0 12208 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_212
timestamp 1698175906
transform 1 0 12544 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_276
timestamp 1698175906
transform 1 0 16128 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_282
timestamp 1698175906
transform 1 0 16464 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_346
timestamp 1698175906
transform 1 0 20048 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_348
timestamp 1698175906
transform 1 0 20160 0 -1 15680
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_2
timestamp 1698175906
transform 1 0 784 0 1 15680
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698175906
transform 1 0 2576 0 1 15680
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_37
timestamp 1698175906
transform 1 0 2744 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_101
timestamp 1698175906
transform 1 0 6328 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_107
timestamp 1698175906
transform 1 0 6664 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_171
timestamp 1698175906
transform 1 0 10248 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_177
timestamp 1698175906
transform 1 0 10584 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_241
timestamp 1698175906
transform 1 0 14168 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_247
timestamp 1698175906
transform 1 0 14504 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_311
timestamp 1698175906
transform 1 0 18088 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_317
timestamp 1698175906
transform 1 0 18424 0 1 15680
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2
timestamp 1698175906
transform 1 0 784 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_66
timestamp 1698175906
transform 1 0 4368 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_72
timestamp 1698175906
transform 1 0 4704 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_136
timestamp 1698175906
transform 1 0 8288 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_142
timestamp 1698175906
transform 1 0 8624 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_206
timestamp 1698175906
transform 1 0 12208 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_212
timestamp 1698175906
transform 1 0 12544 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_276
timestamp 1698175906
transform 1 0 16128 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_282
timestamp 1698175906
transform 1 0 16464 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_346
timestamp 1698175906
transform 1 0 20048 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_348
timestamp 1698175906
transform 1 0 20160 0 -1 16464
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698175906
transform 1 0 784 0 1 16464
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698175906
transform 1 0 2576 0 1 16464
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_37
timestamp 1698175906
transform 1 0 2744 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_101
timestamp 1698175906
transform 1 0 6328 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_107
timestamp 1698175906
transform 1 0 6664 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_171
timestamp 1698175906
transform 1 0 10248 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_177
timestamp 1698175906
transform 1 0 10584 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_241
timestamp 1698175906
transform 1 0 14168 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_247
timestamp 1698175906
transform 1 0 14504 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_311
timestamp 1698175906
transform 1 0 18088 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_317
timestamp 1698175906
transform 1 0 18424 0 1 16464
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_2
timestamp 1698175906
transform 1 0 784 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_66
timestamp 1698175906
transform 1 0 4368 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_72
timestamp 1698175906
transform 1 0 4704 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_136
timestamp 1698175906
transform 1 0 8288 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_142
timestamp 1698175906
transform 1 0 8624 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_206
timestamp 1698175906
transform 1 0 12208 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_212
timestamp 1698175906
transform 1 0 12544 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_276
timestamp 1698175906
transform 1 0 16128 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_282
timestamp 1698175906
transform 1 0 16464 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_346
timestamp 1698175906
transform 1 0 20048 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_348
timestamp 1698175906
transform 1 0 20160 0 -1 17248
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698175906
transform 1 0 784 0 1 17248
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698175906
transform 1 0 2576 0 1 17248
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_37
timestamp 1698175906
transform 1 0 2744 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_101
timestamp 1698175906
transform 1 0 6328 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_107
timestamp 1698175906
transform 1 0 6664 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_171
timestamp 1698175906
transform 1 0 10248 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_177
timestamp 1698175906
transform 1 0 10584 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_241
timestamp 1698175906
transform 1 0 14168 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_247
timestamp 1698175906
transform 1 0 14504 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_311
timestamp 1698175906
transform 1 0 18088 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_317
timestamp 1698175906
transform 1 0 18424 0 1 17248
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2
timestamp 1698175906
transform 1 0 784 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1698175906
transform 1 0 4368 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_72
timestamp 1698175906
transform 1 0 4704 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_136
timestamp 1698175906
transform 1 0 8288 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_142
timestamp 1698175906
transform 1 0 8624 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_206
timestamp 1698175906
transform 1 0 12208 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_212
timestamp 1698175906
transform 1 0 12544 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_276
timestamp 1698175906
transform 1 0 16128 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_282
timestamp 1698175906
transform 1 0 16464 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_346
timestamp 1698175906
transform 1 0 20048 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_348
timestamp 1698175906
transform 1 0 20160 0 -1 18032
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_2
timestamp 1698175906
transform 1 0 784 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698175906
transform 1 0 2576 0 1 18032
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_37
timestamp 1698175906
transform 1 0 2744 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_101
timestamp 1698175906
transform 1 0 6328 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_107
timestamp 1698175906
transform 1 0 6664 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_171
timestamp 1698175906
transform 1 0 10248 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_177
timestamp 1698175906
transform 1 0 10584 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_241
timestamp 1698175906
transform 1 0 14168 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_247
timestamp 1698175906
transform 1 0 14504 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_311
timestamp 1698175906
transform 1 0 18088 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_317
timestamp 1698175906
transform 1 0 18424 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_2
timestamp 1698175906
transform 1 0 784 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_66
timestamp 1698175906
transform 1 0 4368 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_72
timestamp 1698175906
transform 1 0 4704 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_136
timestamp 1698175906
transform 1 0 8288 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_142
timestamp 1698175906
transform 1 0 8624 0 -1 18816
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_150
timestamp 1698175906
transform 1 0 9072 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_154
timestamp 1698175906
transform 1 0 9296 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_156
timestamp 1698175906
transform 1 0 9408 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_183
timestamp 1698175906
transform 1 0 10920 0 -1 18816
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_199
timestamp 1698175906
transform 1 0 11816 0 -1 18816
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_207
timestamp 1698175906
transform 1 0 12264 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_209
timestamp 1698175906
transform 1 0 12376 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_216
timestamp 1698175906
transform 1 0 12768 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_243
timestamp 1698175906
transform 1 0 14280 0 -1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_275
timestamp 1698175906
transform 1 0 16072 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_279
timestamp 1698175906
transform 1 0 16296 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_282
timestamp 1698175906
transform 1 0 16464 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_346
timestamp 1698175906
transform 1 0 20048 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_348
timestamp 1698175906
transform 1 0 20160 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_2
timestamp 1698175906
transform 1 0 784 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_36
timestamp 1698175906
transform 1 0 2688 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_70
timestamp 1698175906
transform 1 0 4592 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_104
timestamp 1698175906
transform 1 0 6496 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_138
timestamp 1698175906
transform 1 0 8400 0 1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_165
timestamp 1698175906
transform 1 0 9912 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_169
timestamp 1698175906
transform 1 0 10136 0 1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_198
timestamp 1698175906
transform 1 0 11760 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_202
timestamp 1698175906
transform 1 0 11984 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_232
timestamp 1698175906
transform 1 0 13664 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_236
timestamp 1698175906
transform 1 0 13888 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_266
timestamp 1698175906
transform 1 0 15568 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_270
timestamp 1698175906
transform 1 0 15792 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_274
timestamp 1698175906
transform 1 0 16016 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_308
timestamp 1698175906
transform 1 0 17920 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_342
timestamp 1698175906
transform 1 0 19824 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_346
timestamp 1698175906
transform 1 0 20048 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_348
timestamp 1698175906
transform 1 0 20160 0 1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita27_24 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19992 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita27_25
timestamp 1698175906
transform -1 0 9352 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita27_26
timestamp 1698175906
transform -1 0 12768 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18760 0 -1 8624
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output2
timestamp 1698175906
transform 1 0 13160 0 -1 2352
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output3
timestamp 1698175906
transform 1 0 18760 0 -1 10976
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output4
timestamp 1698175906
transform -1 0 2240 0 1 10976
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output5
timestamp 1698175906
transform -1 0 2240 0 1 8624
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output6
timestamp 1698175906
transform 1 0 18760 0 1 12544
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output7
timestamp 1698175906
transform -1 0 2240 0 -1 9408
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output8
timestamp 1698175906
transform 1 0 14112 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output9
timestamp 1698175906
transform 1 0 12824 0 -1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output10
timestamp 1698175906
transform 1 0 18760 0 1 8624
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output11
timestamp 1698175906
transform 1 0 10808 0 -1 2352
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output12
timestamp 1698175906
transform 1 0 8456 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output13
timestamp 1698175906
transform -1 0 2240 0 -1 10976
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output14
timestamp 1698175906
transform -1 0 12096 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output15
timestamp 1698175906
transform 1 0 10304 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output16
timestamp 1698175906
transform 1 0 9464 0 -1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output17
timestamp 1698175906
transform 1 0 12208 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output18
timestamp 1698175906
transform 1 0 18760 0 1 11760
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output19
timestamp 1698175906
transform -1 0 2240 0 -1 13328
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output20
timestamp 1698175906
transform 1 0 18760 0 -1 10192
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output21
timestamp 1698175906
transform -1 0 2240 0 1 11760
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output22
timestamp 1698175906
transform 1 0 9352 0 -1 2352
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output23
timestamp 1698175906
transform 1 0 18760 0 -1 13328
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_45 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 672 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698175906
transform -1 0 20328 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_46
timestamp 1698175906
transform 1 0 672 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698175906
transform -1 0 20328 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_47
timestamp 1698175906
transform 1 0 672 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698175906
transform -1 0 20328 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_48
timestamp 1698175906
transform 1 0 672 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698175906
transform -1 0 20328 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_49
timestamp 1698175906
transform 1 0 672 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698175906
transform -1 0 20328 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_50
timestamp 1698175906
transform 1 0 672 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698175906
transform -1 0 20328 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_51
timestamp 1698175906
transform 1 0 672 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698175906
transform -1 0 20328 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_52
timestamp 1698175906
transform 1 0 672 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698175906
transform -1 0 20328 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_53
timestamp 1698175906
transform 1 0 672 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698175906
transform -1 0 20328 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_54
timestamp 1698175906
transform 1 0 672 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698175906
transform -1 0 20328 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_55
timestamp 1698175906
transform 1 0 672 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698175906
transform -1 0 20328 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_56
timestamp 1698175906
transform 1 0 672 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698175906
transform -1 0 20328 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_57
timestamp 1698175906
transform 1 0 672 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698175906
transform -1 0 20328 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_58
timestamp 1698175906
transform 1 0 672 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698175906
transform -1 0 20328 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_59
timestamp 1698175906
transform 1 0 672 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698175906
transform -1 0 20328 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_60
timestamp 1698175906
transform 1 0 672 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698175906
transform -1 0 20328 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_61
timestamp 1698175906
transform 1 0 672 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698175906
transform -1 0 20328 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_62
timestamp 1698175906
transform 1 0 672 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698175906
transform -1 0 20328 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_63
timestamp 1698175906
transform 1 0 672 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698175906
transform -1 0 20328 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_64
timestamp 1698175906
transform 1 0 672 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698175906
transform -1 0 20328 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_65
timestamp 1698175906
transform 1 0 672 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698175906
transform -1 0 20328 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_66
timestamp 1698175906
transform 1 0 672 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698175906
transform -1 0 20328 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_67
timestamp 1698175906
transform 1 0 672 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698175906
transform -1 0 20328 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_68
timestamp 1698175906
transform 1 0 672 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698175906
transform -1 0 20328 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_69
timestamp 1698175906
transform 1 0 672 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698175906
transform -1 0 20328 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_70
timestamp 1698175906
transform 1 0 672 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698175906
transform -1 0 20328 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_71
timestamp 1698175906
transform 1 0 672 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698175906
transform -1 0 20328 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_72
timestamp 1698175906
transform 1 0 672 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698175906
transform -1 0 20328 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_73
timestamp 1698175906
transform 1 0 672 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698175906
transform -1 0 20328 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_74
timestamp 1698175906
transform 1 0 672 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698175906
transform -1 0 20328 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_75
timestamp 1698175906
transform 1 0 672 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698175906
transform -1 0 20328 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_76
timestamp 1698175906
transform 1 0 672 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698175906
transform -1 0 20328 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_77
timestamp 1698175906
transform 1 0 672 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698175906
transform -1 0 20328 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_78
timestamp 1698175906
transform 1 0 672 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698175906
transform -1 0 20328 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_79
timestamp 1698175906
transform 1 0 672 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698175906
transform -1 0 20328 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_80
timestamp 1698175906
transform 1 0 672 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698175906
transform -1 0 20328 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_81
timestamp 1698175906
transform 1 0 672 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698175906
transform -1 0 20328 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_82
timestamp 1698175906
transform 1 0 672 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698175906
transform -1 0 20328 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_83
timestamp 1698175906
transform 1 0 672 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698175906
transform -1 0 20328 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_84
timestamp 1698175906
transform 1 0 672 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698175906
transform -1 0 20328 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_85
timestamp 1698175906
transform 1 0 672 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698175906
transform -1 0 20328 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_86
timestamp 1698175906
transform 1 0 672 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698175906
transform -1 0 20328 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_87
timestamp 1698175906
transform 1 0 672 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698175906
transform -1 0 20328 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_88
timestamp 1698175906
transform 1 0 672 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698175906
transform -1 0 20328 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_89
timestamp 1698175906
transform 1 0 672 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698175906
transform -1 0 20328 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_90 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 2576 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_91
timestamp 1698175906
transform 1 0 4480 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_92
timestamp 1698175906
transform 1 0 6384 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_93
timestamp 1698175906
transform 1 0 8288 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_94
timestamp 1698175906
transform 1 0 10192 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_95
timestamp 1698175906
transform 1 0 12096 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_96
timestamp 1698175906
transform 1 0 14000 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_97
timestamp 1698175906
transform 1 0 15904 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_98
timestamp 1698175906
transform 1 0 17808 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_99
timestamp 1698175906
transform 1 0 19712 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_100
timestamp 1698175906
transform 1 0 4592 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_101
timestamp 1698175906
transform 1 0 8512 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_102
timestamp 1698175906
transform 1 0 12432 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_103
timestamp 1698175906
transform 1 0 16352 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_104
timestamp 1698175906
transform 1 0 2632 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_105
timestamp 1698175906
transform 1 0 6552 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_106
timestamp 1698175906
transform 1 0 10472 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_107
timestamp 1698175906
transform 1 0 14392 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_108
timestamp 1698175906
transform 1 0 18312 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_109
timestamp 1698175906
transform 1 0 4592 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_110
timestamp 1698175906
transform 1 0 8512 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_111
timestamp 1698175906
transform 1 0 12432 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_112
timestamp 1698175906
transform 1 0 16352 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_113
timestamp 1698175906
transform 1 0 2632 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_114
timestamp 1698175906
transform 1 0 6552 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_115
timestamp 1698175906
transform 1 0 10472 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_116
timestamp 1698175906
transform 1 0 14392 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_117
timestamp 1698175906
transform 1 0 18312 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_118
timestamp 1698175906
transform 1 0 4592 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_119
timestamp 1698175906
transform 1 0 8512 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_120
timestamp 1698175906
transform 1 0 12432 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_121
timestamp 1698175906
transform 1 0 16352 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_122
timestamp 1698175906
transform 1 0 2632 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_123
timestamp 1698175906
transform 1 0 6552 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_124
timestamp 1698175906
transform 1 0 10472 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_125
timestamp 1698175906
transform 1 0 14392 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_126
timestamp 1698175906
transform 1 0 18312 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_127
timestamp 1698175906
transform 1 0 4592 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_128
timestamp 1698175906
transform 1 0 8512 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_129
timestamp 1698175906
transform 1 0 12432 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_130
timestamp 1698175906
transform 1 0 16352 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_131
timestamp 1698175906
transform 1 0 2632 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_132
timestamp 1698175906
transform 1 0 6552 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_133
timestamp 1698175906
transform 1 0 10472 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_134
timestamp 1698175906
transform 1 0 14392 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_135
timestamp 1698175906
transform 1 0 18312 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_136
timestamp 1698175906
transform 1 0 4592 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_137
timestamp 1698175906
transform 1 0 8512 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_138
timestamp 1698175906
transform 1 0 12432 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_139
timestamp 1698175906
transform 1 0 16352 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_140
timestamp 1698175906
transform 1 0 2632 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_141
timestamp 1698175906
transform 1 0 6552 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_142
timestamp 1698175906
transform 1 0 10472 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_143
timestamp 1698175906
transform 1 0 14392 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_144
timestamp 1698175906
transform 1 0 18312 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_145
timestamp 1698175906
transform 1 0 4592 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_146
timestamp 1698175906
transform 1 0 8512 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_147
timestamp 1698175906
transform 1 0 12432 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_148
timestamp 1698175906
transform 1 0 16352 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_149
timestamp 1698175906
transform 1 0 2632 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_150
timestamp 1698175906
transform 1 0 6552 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_151
timestamp 1698175906
transform 1 0 10472 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_152
timestamp 1698175906
transform 1 0 14392 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_153
timestamp 1698175906
transform 1 0 18312 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_154
timestamp 1698175906
transform 1 0 4592 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_155
timestamp 1698175906
transform 1 0 8512 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_156
timestamp 1698175906
transform 1 0 12432 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_157
timestamp 1698175906
transform 1 0 16352 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_158
timestamp 1698175906
transform 1 0 2632 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_159
timestamp 1698175906
transform 1 0 6552 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_160
timestamp 1698175906
transform 1 0 10472 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_161
timestamp 1698175906
transform 1 0 14392 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_162
timestamp 1698175906
transform 1 0 18312 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_163
timestamp 1698175906
transform 1 0 4592 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_164
timestamp 1698175906
transform 1 0 8512 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_165
timestamp 1698175906
transform 1 0 12432 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_166
timestamp 1698175906
transform 1 0 16352 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_167
timestamp 1698175906
transform 1 0 2632 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_168
timestamp 1698175906
transform 1 0 6552 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_169
timestamp 1698175906
transform 1 0 10472 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_170
timestamp 1698175906
transform 1 0 14392 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_171
timestamp 1698175906
transform 1 0 18312 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_172
timestamp 1698175906
transform 1 0 4592 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_173
timestamp 1698175906
transform 1 0 8512 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_174
timestamp 1698175906
transform 1 0 12432 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_175
timestamp 1698175906
transform 1 0 16352 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_176
timestamp 1698175906
transform 1 0 2632 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_177
timestamp 1698175906
transform 1 0 6552 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_178
timestamp 1698175906
transform 1 0 10472 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_179
timestamp 1698175906
transform 1 0 14392 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_180
timestamp 1698175906
transform 1 0 18312 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_181
timestamp 1698175906
transform 1 0 4592 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_182
timestamp 1698175906
transform 1 0 8512 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_183
timestamp 1698175906
transform 1 0 12432 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_184
timestamp 1698175906
transform 1 0 16352 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_185
timestamp 1698175906
transform 1 0 2632 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_186
timestamp 1698175906
transform 1 0 6552 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_187
timestamp 1698175906
transform 1 0 10472 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_188
timestamp 1698175906
transform 1 0 14392 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_189
timestamp 1698175906
transform 1 0 18312 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_190
timestamp 1698175906
transform 1 0 4592 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_191
timestamp 1698175906
transform 1 0 8512 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_192
timestamp 1698175906
transform 1 0 12432 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_193
timestamp 1698175906
transform 1 0 16352 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_194
timestamp 1698175906
transform 1 0 2632 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_195
timestamp 1698175906
transform 1 0 6552 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_196
timestamp 1698175906
transform 1 0 10472 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_197
timestamp 1698175906
transform 1 0 14392 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_198
timestamp 1698175906
transform 1 0 18312 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_199
timestamp 1698175906
transform 1 0 4592 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_200
timestamp 1698175906
transform 1 0 8512 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_201
timestamp 1698175906
transform 1 0 12432 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_202
timestamp 1698175906
transform 1 0 16352 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_203
timestamp 1698175906
transform 1 0 2632 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_204
timestamp 1698175906
transform 1 0 6552 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_205
timestamp 1698175906
transform 1 0 10472 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_206
timestamp 1698175906
transform 1 0 14392 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_207
timestamp 1698175906
transform 1 0 18312 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_208
timestamp 1698175906
transform 1 0 4592 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_209
timestamp 1698175906
transform 1 0 8512 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_210
timestamp 1698175906
transform 1 0 12432 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_211
timestamp 1698175906
transform 1 0 16352 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_212
timestamp 1698175906
transform 1 0 2632 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_213
timestamp 1698175906
transform 1 0 6552 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_214
timestamp 1698175906
transform 1 0 10472 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_215
timestamp 1698175906
transform 1 0 14392 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_216
timestamp 1698175906
transform 1 0 18312 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_217
timestamp 1698175906
transform 1 0 4592 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_218
timestamp 1698175906
transform 1 0 8512 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_219
timestamp 1698175906
transform 1 0 12432 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_220
timestamp 1698175906
transform 1 0 16352 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_221
timestamp 1698175906
transform 1 0 2632 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_222
timestamp 1698175906
transform 1 0 6552 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_223
timestamp 1698175906
transform 1 0 10472 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_224
timestamp 1698175906
transform 1 0 14392 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_225
timestamp 1698175906
transform 1 0 18312 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_226
timestamp 1698175906
transform 1 0 4592 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_227
timestamp 1698175906
transform 1 0 8512 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_228
timestamp 1698175906
transform 1 0 12432 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_229
timestamp 1698175906
transform 1 0 16352 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_230
timestamp 1698175906
transform 1 0 2632 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_231
timestamp 1698175906
transform 1 0 6552 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_232
timestamp 1698175906
transform 1 0 10472 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_233
timestamp 1698175906
transform 1 0 14392 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_234
timestamp 1698175906
transform 1 0 18312 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_235
timestamp 1698175906
transform 1 0 4592 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_236
timestamp 1698175906
transform 1 0 8512 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_237
timestamp 1698175906
transform 1 0 12432 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_238
timestamp 1698175906
transform 1 0 16352 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_239
timestamp 1698175906
transform 1 0 2632 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_240
timestamp 1698175906
transform 1 0 6552 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_241
timestamp 1698175906
transform 1 0 10472 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_242
timestamp 1698175906
transform 1 0 14392 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_243
timestamp 1698175906
transform 1 0 18312 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_244
timestamp 1698175906
transform 1 0 4592 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_245
timestamp 1698175906
transform 1 0 8512 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_246
timestamp 1698175906
transform 1 0 12432 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_247
timestamp 1698175906
transform 1 0 16352 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_248
timestamp 1698175906
transform 1 0 2632 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_249
timestamp 1698175906
transform 1 0 6552 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_250
timestamp 1698175906
transform 1 0 10472 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_251
timestamp 1698175906
transform 1 0 14392 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_252
timestamp 1698175906
transform 1 0 18312 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_253
timestamp 1698175906
transform 1 0 4592 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_254
timestamp 1698175906
transform 1 0 8512 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_255
timestamp 1698175906
transform 1 0 12432 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_256
timestamp 1698175906
transform 1 0 16352 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_257
timestamp 1698175906
transform 1 0 2632 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_258
timestamp 1698175906
transform 1 0 6552 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_259
timestamp 1698175906
transform 1 0 10472 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_260
timestamp 1698175906
transform 1 0 14392 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_261
timestamp 1698175906
transform 1 0 18312 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_262
timestamp 1698175906
transform 1 0 4592 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_263
timestamp 1698175906
transform 1 0 8512 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_264
timestamp 1698175906
transform 1 0 12432 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_265
timestamp 1698175906
transform 1 0 16352 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_266
timestamp 1698175906
transform 1 0 2632 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_267
timestamp 1698175906
transform 1 0 6552 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_268
timestamp 1698175906
transform 1 0 10472 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_269
timestamp 1698175906
transform 1 0 14392 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_270
timestamp 1698175906
transform 1 0 18312 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_271
timestamp 1698175906
transform 1 0 4592 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_272
timestamp 1698175906
transform 1 0 8512 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_273
timestamp 1698175906
transform 1 0 12432 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_274
timestamp 1698175906
transform 1 0 16352 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_275
timestamp 1698175906
transform 1 0 2632 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_276
timestamp 1698175906
transform 1 0 6552 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_277
timestamp 1698175906
transform 1 0 10472 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_278
timestamp 1698175906
transform 1 0 14392 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_279
timestamp 1698175906
transform 1 0 18312 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_280
timestamp 1698175906
transform 1 0 4592 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_281
timestamp 1698175906
transform 1 0 8512 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_282
timestamp 1698175906
transform 1 0 12432 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_283
timestamp 1698175906
transform 1 0 16352 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_284
timestamp 1698175906
transform 1 0 2632 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_285
timestamp 1698175906
transform 1 0 6552 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_286
timestamp 1698175906
transform 1 0 10472 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_287
timestamp 1698175906
transform 1 0 14392 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_288
timestamp 1698175906
transform 1 0 18312 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_289
timestamp 1698175906
transform 1 0 4592 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_290
timestamp 1698175906
transform 1 0 8512 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_291
timestamp 1698175906
transform 1 0 12432 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_292
timestamp 1698175906
transform 1 0 16352 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_293
timestamp 1698175906
transform 1 0 2576 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_294
timestamp 1698175906
transform 1 0 4480 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_295
timestamp 1698175906
transform 1 0 6384 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_296
timestamp 1698175906
transform 1 0 8288 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_297
timestamp 1698175906
transform 1 0 10192 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_298
timestamp 1698175906
transform 1 0 12096 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_299
timestamp 1698175906
transform 1 0 14000 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_300
timestamp 1698175906
transform 1 0 15904 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_301
timestamp 1698175906
transform 1 0 17808 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_302
timestamp 1698175906
transform 1 0 19712 0 1 18816
box -43 -43 155 435
<< labels >>
flabel metal3 s 0 14112 400 14168 0 FreeSans 224 0 0 0 clk
port 0 nsew signal input
flabel metal3 s 20600 10080 21000 10136 0 FreeSans 224 0 0 0 segm[0]
port 1 nsew signal tristate
flabel metal3 s 20600 8064 21000 8120 0 FreeSans 224 0 0 0 segm[10]
port 2 nsew signal tristate
flabel metal2 s 13104 0 13160 400 0 FreeSans 224 90 0 0 segm[11]
port 3 nsew signal tristate
flabel metal3 s 20600 10416 21000 10472 0 FreeSans 224 0 0 0 segm[12]
port 4 nsew signal tristate
flabel metal3 s 0 11088 400 11144 0 FreeSans 224 0 0 0 segm[13]
port 5 nsew signal tristate
flabel metal3 s 0 8736 400 8792 0 FreeSans 224 0 0 0 segm[1]
port 6 nsew signal tristate
flabel metal3 s 20600 12432 21000 12488 0 FreeSans 224 0 0 0 segm[2]
port 7 nsew signal tristate
flabel metal2 s 9072 0 9128 400 0 FreeSans 224 90 0 0 segm[3]
port 8 nsew signal tristate
flabel metal3 s 0 9072 400 9128 0 FreeSans 224 0 0 0 segm[4]
port 9 nsew signal tristate
flabel metal2 s 12432 20600 12488 21000 0 FreeSans 224 90 0 0 segm[5]
port 10 nsew signal tristate
flabel metal2 s 13104 20600 13160 21000 0 FreeSans 224 90 0 0 segm[6]
port 11 nsew signal tristate
flabel metal2 s 12768 20600 12824 21000 0 FreeSans 224 90 0 0 segm[7]
port 12 nsew signal tristate
flabel metal3 s 20600 8736 21000 8792 0 FreeSans 224 0 0 0 segm[8]
port 13 nsew signal tristate
flabel metal2 s 10752 0 10808 400 0 FreeSans 224 90 0 0 segm[9]
port 14 nsew signal tristate
flabel metal2 s 8400 20600 8456 21000 0 FreeSans 224 90 0 0 sel[0]
port 15 nsew signal tristate
flabel metal3 s 0 10416 400 10472 0 FreeSans 224 0 0 0 sel[10]
port 16 nsew signal tristate
flabel metal2 s 11088 0 11144 400 0 FreeSans 224 90 0 0 sel[11]
port 17 nsew signal tristate
flabel metal2 s 10080 20600 10136 21000 0 FreeSans 224 90 0 0 sel[1]
port 18 nsew signal tristate
flabel metal2 s 9408 20600 9464 21000 0 FreeSans 224 90 0 0 sel[2]
port 19 nsew signal tristate
flabel metal2 s 11424 20600 11480 21000 0 FreeSans 224 90 0 0 sel[3]
port 20 nsew signal tristate
flabel metal3 s 20600 11760 21000 11816 0 FreeSans 224 0 0 0 sel[4]
port 21 nsew signal tristate
flabel metal3 s 0 12768 400 12824 0 FreeSans 224 0 0 0 sel[5]
port 22 nsew signal tristate
flabel metal3 s 20600 9744 21000 9800 0 FreeSans 224 0 0 0 sel[6]
port 23 nsew signal tristate
flabel metal3 s 0 11760 400 11816 0 FreeSans 224 0 0 0 sel[7]
port 24 nsew signal tristate
flabel metal2 s 9744 0 9800 400 0 FreeSans 224 90 0 0 sel[8]
port 25 nsew signal tristate
flabel metal3 s 20600 12768 21000 12824 0 FreeSans 224 0 0 0 sel[9]
port 26 nsew signal tristate
flabel metal4 s 2224 1538 2384 19238 0 FreeSans 640 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 17584 1538 17744 19238 0 FreeSans 640 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 9904 1538 10064 19238 0 FreeSans 640 90 0 0 vss
port 28 nsew ground bidirectional
rlabel metal1 10500 19208 10500 19208 0 vdd
rlabel metal1 10500 18816 10500 18816 0 vss
rlabel metal2 6188 11788 6188 11788 0 _000_
rlabel metal2 13748 9296 13748 9296 0 _001_
rlabel metal2 6580 13048 6580 13048 0 _002_
rlabel metal3 13300 11508 13300 11508 0 _003_
rlabel metal2 10892 14168 10892 14168 0 _004_
rlabel metal2 9044 13888 9044 13888 0 _005_
rlabel metal2 9660 13748 9660 13748 0 _006_
rlabel metal2 7420 13356 7420 13356 0 _007_
rlabel metal2 13804 12516 13804 12516 0 _008_
rlabel metal2 12180 13356 12180 13356 0 _009_
rlabel metal2 11732 12852 11732 12852 0 _010_
rlabel metal2 6748 10948 6748 10948 0 _011_
rlabel metal3 9156 8372 9156 8372 0 _012_
rlabel metal2 5908 9912 5908 9912 0 _013_
rlabel metal2 10220 7112 10220 7112 0 _014_
rlabel metal2 6188 8988 6188 8988 0 _015_
rlabel metal3 12964 8876 12964 8876 0 _016_
rlabel metal2 10780 8204 10780 8204 0 _017_
rlabel metal2 12348 8232 12348 8232 0 _018_
rlabel metal3 12460 7588 12460 7588 0 _019_
rlabel metal3 13440 9940 13440 9940 0 _020_
rlabel metal2 12656 11900 12656 11900 0 _021_
rlabel metal2 7700 11704 7700 11704 0 _022_
rlabel metal2 7364 8596 7364 8596 0 _023_
rlabel metal2 7140 10500 7140 10500 0 _024_
rlabel metal3 9408 13132 9408 13132 0 _025_
rlabel metal2 9660 11228 9660 11228 0 _026_
rlabel metal2 9996 12376 9996 12376 0 _027_
rlabel metal2 9772 13468 9772 13468 0 _028_
rlabel metal3 8428 13076 8428 13076 0 _029_
rlabel metal3 12068 12348 12068 12348 0 _030_
rlabel metal2 13076 12488 13076 12488 0 _031_
rlabel metal3 12516 13132 12516 13132 0 _032_
rlabel metal2 11452 12992 11452 12992 0 _033_
rlabel metal2 7532 10164 7532 10164 0 _034_
rlabel metal3 11788 10444 11788 10444 0 _035_
rlabel metal2 11620 10080 11620 10080 0 _036_
rlabel metal3 12292 12684 12292 12684 0 _037_
rlabel metal3 11704 13076 11704 13076 0 _038_
rlabel metal2 12012 12488 12012 12488 0 _039_
rlabel metal2 7252 11004 7252 11004 0 _040_
rlabel metal2 9436 9632 9436 9632 0 _041_
rlabel metal2 9492 8736 9492 8736 0 _042_
rlabel metal2 7364 11004 7364 11004 0 _043_
rlabel metal2 9548 8232 9548 8232 0 _044_
rlabel metal2 6580 9996 6580 9996 0 _045_
rlabel metal2 6272 10500 6272 10500 0 _046_
rlabel metal2 12516 9408 12516 9408 0 _047_
rlabel metal2 10780 7378 10780 7378 0 _048_
rlabel metal3 11144 7588 11144 7588 0 _049_
rlabel metal3 7364 9184 7364 9184 0 _050_
rlabel metal2 7280 8932 7280 8932 0 _051_
rlabel metal2 7224 9212 7224 9212 0 _052_
rlabel metal2 6356 8960 6356 8960 0 _053_
rlabel metal2 13916 8652 13916 8652 0 _054_
rlabel metal2 12180 9016 12180 9016 0 _055_
rlabel metal2 12880 8428 12880 8428 0 _056_
rlabel metal2 11032 8932 11032 8932 0 _057_
rlabel metal3 11004 8932 11004 8932 0 _058_
rlabel metal2 10668 8596 10668 8596 0 _059_
rlabel metal2 13076 7896 13076 7896 0 _060_
rlabel metal2 12964 8456 12964 8456 0 _061_
rlabel metal2 12852 7266 12852 7266 0 _062_
rlabel metal3 12320 7756 12320 7756 0 _063_
rlabel metal2 13076 10360 13076 10360 0 _064_
rlabel metal2 8904 10780 8904 10780 0 _065_
rlabel metal2 9492 10528 9492 10528 0 _066_
rlabel metal2 7952 9996 7952 9996 0 _067_
rlabel metal2 7588 9408 7588 9408 0 _068_
rlabel metal2 10892 11312 10892 11312 0 _069_
rlabel metal2 10724 11872 10724 11872 0 _070_
rlabel metal2 11844 11368 11844 11368 0 _071_
rlabel metal3 8876 12236 8876 12236 0 _072_
rlabel metal2 8876 9240 8876 9240 0 _073_
rlabel metal2 7420 9044 7420 9044 0 _074_
rlabel metal2 9156 10024 9156 10024 0 _075_
rlabel metal2 10108 10360 10108 10360 0 _076_
rlabel metal2 10836 10472 10836 10472 0 _077_
rlabel metal2 9380 9464 9380 9464 0 _078_
rlabel metal2 7644 9016 7644 9016 0 _079_
rlabel metal3 8736 10276 8736 10276 0 _080_
rlabel metal3 11536 11508 11536 11508 0 _081_
rlabel metal2 7756 10080 7756 10080 0 _082_
rlabel metal2 7028 11396 7028 11396 0 _083_
rlabel metal2 9100 9212 9100 9212 0 _084_
rlabel metal2 9772 12236 9772 12236 0 _085_
rlabel metal2 13860 12152 13860 12152 0 _086_
rlabel metal2 7140 12516 7140 12516 0 _087_
rlabel metal2 6356 11732 6356 11732 0 _088_
rlabel metal2 13020 9352 13020 9352 0 _089_
rlabel metal2 11900 10612 11900 10612 0 _090_
rlabel metal3 10808 9492 10808 9492 0 _091_
rlabel metal3 12628 10052 12628 10052 0 _092_
rlabel metal2 13524 9380 13524 9380 0 _093_
rlabel metal2 13944 9492 13944 9492 0 _094_
rlabel metal2 7224 13188 7224 13188 0 _095_
rlabel metal2 6916 12824 6916 12824 0 _096_
rlabel metal2 12656 9212 12656 9212 0 _097_
rlabel metal2 13076 11760 13076 11760 0 _098_
rlabel metal3 11732 13916 11732 13916 0 _099_
rlabel metal3 10976 13972 10976 13972 0 _100_
rlabel metal2 9772 11200 9772 11200 0 _101_
rlabel metal2 9100 11368 9100 11368 0 _102_
rlabel metal2 10724 13678 10724 13678 0 _103_
rlabel metal2 9156 13524 9156 13524 0 _104_
rlabel metal3 1239 14140 1239 14140 0 clk
rlabel metal2 11340 10556 11340 10556 0 clknet_0_clk
rlabel metal2 8932 14112 8932 14112 0 clknet_1_0__leaf_clk
rlabel metal3 11536 14308 11536 14308 0 clknet_1_1__leaf_clk
rlabel metal2 11620 11788 11620 11788 0 dut27.count\[0\]
rlabel metal2 9324 12096 9324 12096 0 dut27.count\[1\]
rlabel metal2 8372 9044 8372 9044 0 dut27.count\[2\]
rlabel metal2 8372 10416 8372 10416 0 dut27.count\[3\]
rlabel metal2 18844 8008 18844 8008 0 net1
rlabel metal2 13972 8680 13972 8680 0 net10
rlabel metal3 10332 7644 10332 7644 0 net11
rlabel metal2 8512 13580 8512 13580 0 net12
rlabel metal2 2156 10556 2156 10556 0 net13
rlabel metal2 11284 6776 11284 6776 0 net14
rlabel metal2 10332 14910 10332 14910 0 net15
rlabel metal2 9436 13552 9436 13552 0 net16
rlabel metal3 11704 14028 11704 14028 0 net17
rlabel metal2 14756 11732 14756 11732 0 net18
rlabel metal2 5516 13104 5516 13104 0 net19
rlabel metal2 13244 3178 13244 3178 0 net2
rlabel metal2 14812 9352 14812 9352 0 net20
rlabel metal3 3178 11956 3178 11956 0 net21
rlabel metal2 9436 3178 9436 3178 0 net22
rlabel metal2 18732 12908 18732 12908 0 net23
rlabel metal2 20132 10192 20132 10192 0 net24
rlabel metal2 9100 1015 9100 1015 0 net25
rlabel metal2 12628 19012 12628 19012 0 net26
rlabel metal2 14588 10402 14588 10402 0 net3
rlabel metal2 5684 10948 5684 10948 0 net4
rlabel metal2 6860 8792 6860 8792 0 net5
rlabel metal2 14644 12684 14644 12684 0 net6
rlabel metal2 5460 9184 5460 9184 0 net7
rlabel metal2 13244 13888 13244 13888 0 net8
rlabel metal2 12824 15960 12824 15960 0 net9
rlabel metal2 20020 8204 20020 8204 0 segm[10]
rlabel metal2 13132 1211 13132 1211 0 segm[11]
rlabel metal2 20020 10556 20020 10556 0 segm[12]
rlabel metal3 679 11116 679 11116 0 segm[13]
rlabel metal3 679 8764 679 8764 0 segm[1]
rlabel metal2 20020 12628 20020 12628 0 segm[2]
rlabel metal3 679 9100 679 9100 0 segm[4]
rlabel metal2 13132 19873 13132 19873 0 segm[6]
rlabel metal2 12796 19957 12796 19957 0 segm[7]
rlabel metal2 20020 8820 20020 8820 0 segm[8]
rlabel metal2 10780 1211 10780 1211 0 segm[9]
rlabel metal2 8428 19873 8428 19873 0 sel[0]
rlabel metal3 679 10444 679 10444 0 sel[10]
rlabel metal2 11116 1043 11116 1043 0 sel[11]
rlabel metal2 10108 19873 10108 19873 0 sel[1]
rlabel metal3 9744 18732 9744 18732 0 sel[2]
rlabel metal2 11452 19873 11452 19873 0 sel[3]
rlabel metal2 20020 11900 20020 11900 0 sel[4]
rlabel metal3 679 12796 679 12796 0 sel[5]
rlabel metal2 20020 9828 20020 9828 0 sel[6]
rlabel metal3 679 11788 679 11788 0 sel[7]
rlabel metal2 9772 1211 9772 1211 0 sel[8]
rlabel metal2 19964 12936 19964 12936 0 sel[9]
<< properties >>
string FIXED_BBOX 0 0 21000 21000
<< end >>
