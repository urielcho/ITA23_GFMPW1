magic
tech gf180mcuD
magscale 1 5
timestamp 1699641671
<< metal1 >>
rect 672 19221 20328 19238
rect 672 19195 2239 19221
rect 2265 19195 2291 19221
rect 2317 19195 2343 19221
rect 2369 19195 17599 19221
rect 17625 19195 17651 19221
rect 17677 19195 17703 19221
rect 17729 19195 20328 19221
rect 672 19178 20328 19195
rect 7687 19137 7713 19143
rect 7687 19105 7713 19111
rect 9311 19137 9337 19143
rect 9311 19105 9337 19111
rect 11215 19137 11241 19143
rect 11215 19105 11241 19111
rect 12783 19137 12809 19143
rect 12783 19105 12809 19111
rect 7961 18999 7967 19025
rect 7993 18999 7999 19025
rect 8969 18999 8975 19025
rect 9001 18999 9007 19025
rect 10873 18999 10879 19025
rect 10905 18999 10911 19025
rect 12273 18999 12279 19025
rect 12305 18999 12311 19025
rect 672 18829 20328 18846
rect 672 18803 9919 18829
rect 9945 18803 9971 18829
rect 9997 18803 10023 18829
rect 10049 18803 20328 18829
rect 672 18786 20328 18803
rect 9367 18745 9393 18751
rect 9367 18713 9393 18719
rect 11047 18745 11073 18751
rect 11047 18713 11073 18719
rect 8857 18607 8863 18633
rect 8889 18607 8895 18633
rect 10593 18607 10599 18633
rect 10625 18607 10631 18633
rect 672 18437 20328 18454
rect 672 18411 2239 18437
rect 2265 18411 2291 18437
rect 2317 18411 2343 18437
rect 2369 18411 17599 18437
rect 17625 18411 17651 18437
rect 17677 18411 17703 18437
rect 17729 18411 20328 18437
rect 672 18394 20328 18411
rect 9031 18353 9057 18359
rect 9031 18321 9057 18327
rect 8521 18215 8527 18241
rect 8553 18215 8559 18241
rect 672 18045 20328 18062
rect 672 18019 9919 18045
rect 9945 18019 9971 18045
rect 9997 18019 10023 18045
rect 10049 18019 20328 18045
rect 672 18002 20328 18019
rect 672 17653 20328 17670
rect 672 17627 2239 17653
rect 2265 17627 2291 17653
rect 2317 17627 2343 17653
rect 2369 17627 17599 17653
rect 17625 17627 17651 17653
rect 17677 17627 17703 17653
rect 17729 17627 20328 17653
rect 672 17610 20328 17627
rect 672 17261 20328 17278
rect 672 17235 9919 17261
rect 9945 17235 9971 17261
rect 9997 17235 10023 17261
rect 10049 17235 20328 17261
rect 672 17218 20328 17235
rect 672 16869 20328 16886
rect 672 16843 2239 16869
rect 2265 16843 2291 16869
rect 2317 16843 2343 16869
rect 2369 16843 17599 16869
rect 17625 16843 17651 16869
rect 17677 16843 17703 16869
rect 17729 16843 20328 16869
rect 672 16826 20328 16843
rect 672 16477 20328 16494
rect 672 16451 9919 16477
rect 9945 16451 9971 16477
rect 9997 16451 10023 16477
rect 10049 16451 20328 16477
rect 672 16434 20328 16451
rect 672 16085 20328 16102
rect 672 16059 2239 16085
rect 2265 16059 2291 16085
rect 2317 16059 2343 16085
rect 2369 16059 17599 16085
rect 17625 16059 17651 16085
rect 17677 16059 17703 16085
rect 17729 16059 20328 16085
rect 672 16042 20328 16059
rect 672 15693 20328 15710
rect 672 15667 9919 15693
rect 9945 15667 9971 15693
rect 9997 15667 10023 15693
rect 10049 15667 20328 15693
rect 672 15650 20328 15667
rect 672 15301 20328 15318
rect 672 15275 2239 15301
rect 2265 15275 2291 15301
rect 2317 15275 2343 15301
rect 2369 15275 17599 15301
rect 17625 15275 17651 15301
rect 17677 15275 17703 15301
rect 17729 15275 20328 15301
rect 672 15258 20328 15275
rect 672 14909 20328 14926
rect 672 14883 9919 14909
rect 9945 14883 9971 14909
rect 9997 14883 10023 14909
rect 10049 14883 20328 14909
rect 672 14866 20328 14883
rect 672 14517 20328 14534
rect 672 14491 2239 14517
rect 2265 14491 2291 14517
rect 2317 14491 2343 14517
rect 2369 14491 17599 14517
rect 17625 14491 17651 14517
rect 17677 14491 17703 14517
rect 17729 14491 20328 14517
rect 672 14474 20328 14491
rect 672 14125 20328 14142
rect 672 14099 9919 14125
rect 9945 14099 9971 14125
rect 9997 14099 10023 14125
rect 10049 14099 20328 14125
rect 672 14082 20328 14099
rect 8695 14041 8721 14047
rect 8857 14015 8863 14041
rect 8889 14015 8895 14041
rect 8695 14009 8721 14015
rect 9137 13903 9143 13929
rect 9169 13903 9175 13929
rect 10879 13873 10905 13879
rect 9529 13847 9535 13873
rect 9561 13847 9567 13873
rect 10593 13847 10599 13873
rect 10625 13847 10631 13873
rect 10879 13841 10905 13847
rect 12391 13873 12417 13879
rect 12391 13841 12417 13847
rect 672 13733 20328 13750
rect 672 13707 2239 13733
rect 2265 13707 2291 13733
rect 2317 13707 2343 13733
rect 2369 13707 17599 13733
rect 17625 13707 17651 13733
rect 17677 13707 17703 13733
rect 17729 13707 20328 13733
rect 672 13690 20328 13707
rect 7351 13593 7377 13599
rect 20007 13593 20033 13599
rect 12217 13567 12223 13593
rect 12249 13567 12255 13593
rect 13841 13567 13847 13593
rect 13873 13567 13879 13593
rect 7351 13561 7377 13567
rect 20007 13561 20033 13567
rect 8801 13511 8807 13537
rect 8833 13511 8839 13537
rect 9081 13511 9087 13537
rect 9113 13511 9119 13537
rect 10817 13511 10823 13537
rect 10849 13511 10855 13537
rect 12385 13511 12391 13537
rect 12417 13511 12423 13537
rect 18937 13511 18943 13537
rect 18969 13511 18975 13537
rect 9535 13481 9561 13487
rect 8409 13455 8415 13481
rect 8441 13455 8447 13481
rect 8969 13455 8975 13481
rect 9001 13455 9007 13481
rect 9535 13449 9561 13455
rect 9703 13481 9729 13487
rect 14071 13481 14097 13487
rect 11153 13455 11159 13481
rect 11185 13455 11191 13481
rect 12777 13455 12783 13481
rect 12809 13455 12815 13481
rect 9703 13449 9729 13455
rect 14071 13449 14097 13455
rect 9367 13425 9393 13431
rect 9367 13393 9393 13399
rect 672 13341 20328 13358
rect 672 13315 9919 13341
rect 9945 13315 9971 13341
rect 9997 13315 10023 13341
rect 10049 13315 20328 13341
rect 672 13298 20328 13315
rect 10375 13257 10401 13263
rect 9697 13231 9703 13257
rect 9729 13231 9735 13257
rect 10375 13225 10401 13231
rect 12279 13257 12305 13263
rect 12279 13225 12305 13231
rect 14295 13257 14321 13263
rect 14295 13225 14321 13231
rect 11103 13201 11129 13207
rect 11103 13169 11129 13175
rect 11719 13201 11745 13207
rect 11719 13169 11745 13175
rect 12167 13201 12193 13207
rect 12167 13169 12193 13175
rect 12223 13201 12249 13207
rect 12223 13169 12249 13175
rect 8807 13145 8833 13151
rect 6953 13119 6959 13145
rect 6985 13119 6991 13145
rect 8689 13119 8695 13145
rect 8721 13119 8727 13145
rect 8807 13113 8833 13119
rect 8919 13145 8945 13151
rect 10263 13145 10289 13151
rect 9025 13119 9031 13145
rect 9057 13119 9063 13145
rect 8919 13113 8945 13119
rect 10263 13113 10289 13119
rect 10431 13145 10457 13151
rect 12335 13145 12361 13151
rect 11937 13119 11943 13145
rect 11969 13119 11975 13145
rect 12665 13119 12671 13145
rect 12697 13119 12703 13145
rect 18825 13119 18831 13145
rect 18857 13119 18863 13145
rect 10431 13113 10457 13119
rect 12335 13113 12361 13119
rect 9255 13089 9281 13095
rect 7345 13063 7351 13089
rect 7377 13063 7383 13089
rect 8409 13063 8415 13089
rect 8441 13063 8447 13089
rect 8745 13063 8751 13089
rect 8777 13063 8783 13089
rect 9255 13057 9281 13063
rect 9423 13089 9449 13095
rect 13001 13063 13007 13089
rect 13033 13063 13039 13089
rect 14065 13063 14071 13089
rect 14097 13063 14103 13089
rect 19945 13063 19951 13089
rect 19977 13063 19983 13089
rect 9423 13057 9449 13063
rect 9535 13033 9561 13039
rect 9535 13001 9561 13007
rect 10991 13033 11017 13039
rect 10991 13001 11017 13007
rect 11159 13033 11185 13039
rect 11159 13001 11185 13007
rect 11663 13033 11689 13039
rect 11663 13001 11689 13007
rect 672 12949 20328 12966
rect 672 12923 2239 12949
rect 2265 12923 2291 12949
rect 2317 12923 2343 12949
rect 2369 12923 17599 12949
rect 17625 12923 17651 12949
rect 17677 12923 17703 12949
rect 17729 12923 20328 12949
rect 672 12906 20328 12923
rect 7855 12865 7881 12871
rect 7855 12833 7881 12839
rect 11663 12865 11689 12871
rect 11663 12833 11689 12839
rect 12335 12865 12361 12871
rect 12335 12833 12361 12839
rect 13679 12865 13705 12871
rect 13679 12833 13705 12839
rect 10039 12809 10065 12815
rect 13511 12809 13537 12815
rect 11209 12783 11215 12809
rect 11241 12783 11247 12809
rect 12833 12783 12839 12809
rect 12865 12783 12871 12809
rect 10039 12777 10065 12783
rect 13511 12777 13537 12783
rect 13735 12809 13761 12815
rect 13735 12777 13761 12783
rect 9031 12753 9057 12759
rect 8913 12727 8919 12753
rect 8945 12727 8951 12753
rect 9031 12721 9057 12727
rect 10095 12753 10121 12759
rect 10655 12753 10681 12759
rect 10257 12727 10263 12753
rect 10289 12727 10295 12753
rect 10095 12721 10121 12727
rect 10655 12721 10681 12727
rect 10767 12753 10793 12759
rect 10767 12721 10793 12727
rect 10935 12753 10961 12759
rect 11607 12753 11633 12759
rect 11153 12727 11159 12753
rect 11185 12727 11191 12753
rect 10935 12721 10961 12727
rect 11607 12721 11633 12727
rect 12391 12753 12417 12759
rect 12391 12721 12417 12727
rect 12783 12753 12809 12759
rect 12783 12721 12809 12727
rect 13455 12753 13481 12759
rect 13455 12721 13481 12727
rect 7911 12697 7937 12703
rect 7911 12665 7937 12671
rect 8583 12697 8609 12703
rect 8583 12665 8609 12671
rect 8695 12697 8721 12703
rect 8695 12665 8721 12671
rect 9143 12697 9169 12703
rect 9143 12665 9169 12671
rect 9199 12697 9225 12703
rect 11439 12697 11465 12703
rect 11321 12671 11327 12697
rect 11353 12671 11359 12697
rect 9199 12665 9225 12671
rect 11439 12665 11465 12671
rect 12503 12697 12529 12703
rect 12665 12671 12671 12697
rect 12697 12671 12703 12697
rect 12503 12665 12529 12671
rect 8527 12641 8553 12647
rect 8527 12609 8553 12615
rect 8639 12641 8665 12647
rect 8639 12609 8665 12615
rect 9983 12641 10009 12647
rect 9983 12609 10009 12615
rect 10599 12641 10625 12647
rect 10599 12609 10625 12615
rect 10879 12641 10905 12647
rect 10879 12609 10905 12615
rect 672 12557 20328 12574
rect 672 12531 9919 12557
rect 9945 12531 9971 12557
rect 9997 12531 10023 12557
rect 10049 12531 20328 12557
rect 672 12514 20328 12531
rect 10033 12391 10039 12417
rect 10065 12391 10071 12417
rect 11327 12361 11353 12367
rect 9641 12335 9647 12361
rect 9673 12335 9679 12361
rect 11327 12329 11353 12335
rect 11097 12279 11103 12305
rect 11129 12279 11135 12305
rect 672 12165 20328 12182
rect 672 12139 2239 12165
rect 2265 12139 2291 12165
rect 2317 12139 2343 12165
rect 2369 12139 17599 12165
rect 17625 12139 17651 12165
rect 17677 12139 17703 12165
rect 17729 12139 20328 12165
rect 672 12122 20328 12139
rect 967 12025 993 12031
rect 20007 12025 20033 12031
rect 10817 11999 10823 12025
rect 10849 11999 10855 12025
rect 967 11993 993 11999
rect 20007 11993 20033 11999
rect 13063 11969 13089 11975
rect 2137 11943 2143 11969
rect 2169 11943 2175 11969
rect 11041 11943 11047 11969
rect 11073 11943 11079 11969
rect 18825 11943 18831 11969
rect 18857 11943 18863 11969
rect 13063 11937 13089 11943
rect 9143 11913 9169 11919
rect 7457 11887 7463 11913
rect 7489 11887 7495 11913
rect 9143 11881 9169 11887
rect 9311 11913 9337 11919
rect 9311 11881 9337 11887
rect 10823 11913 10849 11919
rect 10823 11881 10849 11887
rect 12671 11913 12697 11919
rect 12671 11881 12697 11887
rect 12727 11913 12753 11919
rect 12727 11881 12753 11887
rect 12839 11913 12865 11919
rect 12839 11881 12865 11887
rect 12951 11913 12977 11919
rect 12951 11881 12977 11887
rect 13231 11913 13257 11919
rect 13231 11881 13257 11887
rect 7631 11857 7657 11863
rect 7631 11825 7657 11831
rect 10655 11857 10681 11863
rect 10655 11825 10681 11831
rect 10767 11857 10793 11863
rect 10767 11825 10793 11831
rect 13007 11857 13033 11863
rect 13007 11825 13033 11831
rect 672 11773 20328 11790
rect 672 11747 9919 11773
rect 9945 11747 9971 11773
rect 9997 11747 10023 11773
rect 10049 11747 20328 11773
rect 672 11730 20328 11747
rect 9753 11663 9759 11689
rect 9785 11663 9791 11689
rect 9143 11633 9169 11639
rect 13001 11607 13007 11633
rect 13033 11607 13039 11633
rect 9143 11601 9169 11607
rect 7687 11577 7713 11583
rect 2137 11551 2143 11577
rect 2169 11551 2175 11577
rect 7401 11551 7407 11577
rect 7433 11551 7439 11577
rect 7687 11545 7713 11551
rect 7743 11577 7769 11583
rect 7743 11545 7769 11551
rect 7855 11577 7881 11583
rect 9087 11577 9113 11583
rect 7961 11551 7967 11577
rect 7993 11551 7999 11577
rect 9641 11551 9647 11577
rect 9673 11551 9679 11577
rect 12609 11551 12615 11577
rect 12641 11551 12647 11577
rect 14289 11551 14295 11577
rect 14321 11551 14327 11577
rect 18937 11551 18943 11577
rect 18969 11551 18975 11577
rect 7855 11545 7881 11551
rect 9087 11545 9113 11551
rect 7799 11521 7825 11527
rect 6001 11495 6007 11521
rect 6033 11495 6039 11521
rect 7065 11495 7071 11521
rect 7097 11495 7103 11521
rect 7799 11489 7825 11495
rect 8191 11521 8217 11527
rect 15919 11521 15945 11527
rect 14065 11495 14071 11521
rect 14097 11495 14103 11521
rect 14625 11495 14631 11521
rect 14657 11495 14663 11521
rect 15689 11495 15695 11521
rect 15721 11495 15727 11521
rect 8191 11489 8217 11495
rect 15919 11489 15945 11495
rect 967 11465 993 11471
rect 967 11433 993 11439
rect 9143 11465 9169 11471
rect 9143 11433 9169 11439
rect 20007 11465 20033 11471
rect 20007 11433 20033 11439
rect 672 11381 20328 11398
rect 672 11355 2239 11381
rect 2265 11355 2291 11381
rect 2317 11355 2343 11381
rect 2369 11355 17599 11381
rect 17625 11355 17651 11381
rect 17677 11355 17703 11381
rect 17729 11355 20328 11381
rect 672 11338 20328 11355
rect 8639 11297 8665 11303
rect 8017 11271 8023 11297
rect 8049 11271 8055 11297
rect 8639 11265 8665 11271
rect 13959 11297 13985 11303
rect 13959 11265 13985 11271
rect 967 11241 993 11247
rect 967 11209 993 11215
rect 6791 11241 6817 11247
rect 14183 11241 14209 11247
rect 7121 11215 7127 11241
rect 7153 11215 7159 11241
rect 6791 11209 6817 11215
rect 14183 11209 14209 11215
rect 20007 11241 20033 11247
rect 20007 11209 20033 11215
rect 7743 11185 7769 11191
rect 2137 11159 2143 11185
rect 2169 11159 2175 11185
rect 7743 11153 7769 11159
rect 7855 11185 7881 11191
rect 7855 11153 7881 11159
rect 8807 11185 8833 11191
rect 8807 11153 8833 11159
rect 8919 11185 8945 11191
rect 8919 11153 8945 11159
rect 9031 11185 9057 11191
rect 12335 11185 12361 11191
rect 13343 11185 13369 11191
rect 9473 11159 9479 11185
rect 9505 11159 9511 11185
rect 11433 11159 11439 11185
rect 11465 11159 11471 11185
rect 12609 11159 12615 11185
rect 12641 11159 12647 11185
rect 13057 11159 13063 11185
rect 13089 11159 13095 11185
rect 18825 11159 18831 11185
rect 18857 11159 18863 11185
rect 9031 11153 9057 11159
rect 12335 11153 12361 11159
rect 13343 11153 13369 11159
rect 7183 11129 7209 11135
rect 7183 11097 7209 11103
rect 7407 11129 7433 11135
rect 7407 11097 7433 11103
rect 8303 11129 8329 11135
rect 8303 11097 8329 11103
rect 8471 11129 8497 11135
rect 8471 11097 8497 11103
rect 8751 11129 8777 11135
rect 11999 11129 12025 11135
rect 9585 11103 9591 11129
rect 9617 11103 9623 11129
rect 9753 11103 9759 11129
rect 9785 11103 9791 11129
rect 10705 11103 10711 11129
rect 10737 11103 10743 11129
rect 11545 11103 11551 11129
rect 11577 11103 11583 11129
rect 11713 11103 11719 11129
rect 11745 11103 11751 11129
rect 8751 11097 8777 11103
rect 11999 11097 12025 11103
rect 12391 11129 12417 11135
rect 13287 11129 13313 11135
rect 13001 11103 13007 11129
rect 13033 11103 13039 11129
rect 12391 11097 12417 11103
rect 13287 11097 13313 11103
rect 13399 11129 13425 11135
rect 13791 11129 13817 11135
rect 13617 11103 13623 11129
rect 13649 11103 13655 11129
rect 13399 11097 13425 11103
rect 13791 11097 13817 11103
rect 13903 11129 13929 11135
rect 13903 11097 13929 11103
rect 6735 11073 6761 11079
rect 6735 11041 6761 11047
rect 7127 11073 7153 11079
rect 7127 11041 7153 11047
rect 7295 11073 7321 11079
rect 10879 11073 10905 11079
rect 11215 11073 11241 11079
rect 9809 11047 9815 11073
rect 9841 11047 9847 11073
rect 11041 11047 11047 11073
rect 11073 11047 11079 11073
rect 7295 11041 7321 11047
rect 10879 11041 10905 11047
rect 11215 11041 11241 11047
rect 14743 11073 14769 11079
rect 14905 11047 14911 11073
rect 14937 11047 14943 11073
rect 14743 11041 14769 11047
rect 672 10989 20328 11006
rect 672 10963 9919 10989
rect 9945 10963 9971 10989
rect 9997 10963 10023 10989
rect 10049 10963 20328 10989
rect 672 10946 20328 10963
rect 7463 10905 7489 10911
rect 7463 10873 7489 10879
rect 7519 10905 7545 10911
rect 7519 10873 7545 10879
rect 7687 10905 7713 10911
rect 7687 10873 7713 10879
rect 7799 10905 7825 10911
rect 9311 10905 9337 10911
rect 13399 10905 13425 10911
rect 8913 10879 8919 10905
rect 8945 10879 8951 10905
rect 10537 10879 10543 10905
rect 10569 10879 10575 10905
rect 7799 10873 7825 10879
rect 9311 10873 9337 10879
rect 13399 10873 13425 10879
rect 13511 10905 13537 10911
rect 13511 10873 13537 10879
rect 7295 10849 7321 10855
rect 6673 10823 6679 10849
rect 6705 10823 6711 10849
rect 7295 10817 7321 10823
rect 7407 10793 7433 10799
rect 7065 10767 7071 10793
rect 7097 10767 7103 10793
rect 7407 10761 7433 10767
rect 7855 10793 7881 10799
rect 7855 10761 7881 10767
rect 9087 10793 9113 10799
rect 9087 10761 9113 10767
rect 9255 10793 9281 10799
rect 10711 10793 10737 10799
rect 13567 10793 13593 10799
rect 9809 10767 9815 10793
rect 9841 10767 9847 10793
rect 11153 10767 11159 10793
rect 11185 10767 11191 10793
rect 11489 10767 11495 10793
rect 11521 10767 11527 10793
rect 14065 10767 14071 10793
rect 14097 10767 14103 10793
rect 9255 10761 9281 10767
rect 10711 10761 10737 10767
rect 13567 10761 13593 10767
rect 8079 10737 8105 10743
rect 5609 10711 5615 10737
rect 5641 10711 5647 10737
rect 8079 10705 8105 10711
rect 9591 10737 9617 10743
rect 9591 10705 9617 10711
rect 10375 10737 10401 10743
rect 10375 10705 10401 10711
rect 11103 10737 11129 10743
rect 12111 10737 12137 10743
rect 11601 10711 11607 10737
rect 11633 10711 11639 10737
rect 11993 10711 11999 10737
rect 12025 10711 12031 10737
rect 11103 10705 11129 10711
rect 12111 10705 12137 10711
rect 12335 10737 12361 10743
rect 15695 10737 15721 10743
rect 14401 10711 14407 10737
rect 14433 10711 14439 10737
rect 15465 10711 15471 10737
rect 15497 10711 15503 10737
rect 12335 10705 12361 10711
rect 15695 10705 15721 10711
rect 12279 10681 12305 10687
rect 12279 10649 12305 10655
rect 672 10597 20328 10614
rect 672 10571 2239 10597
rect 2265 10571 2291 10597
rect 2317 10571 2343 10597
rect 2369 10571 17599 10597
rect 17625 10571 17651 10597
rect 17677 10571 17703 10597
rect 17729 10571 20328 10597
rect 672 10554 20328 10571
rect 7351 10513 7377 10519
rect 7351 10481 7377 10487
rect 967 10457 993 10463
rect 7183 10457 7209 10463
rect 4993 10431 4999 10457
rect 5025 10431 5031 10457
rect 967 10425 993 10431
rect 7183 10425 7209 10431
rect 8527 10457 8553 10463
rect 14015 10457 14041 10463
rect 20007 10457 20033 10463
rect 9753 10431 9759 10457
rect 9785 10431 9791 10457
rect 16025 10431 16031 10457
rect 16057 10431 16063 10457
rect 8527 10425 8553 10431
rect 14015 10425 14041 10431
rect 20007 10425 20033 10431
rect 7687 10401 7713 10407
rect 2137 10375 2143 10401
rect 2169 10375 2175 10401
rect 6449 10375 6455 10401
rect 6481 10375 6487 10401
rect 7687 10369 7713 10375
rect 8583 10401 8609 10407
rect 8913 10375 8919 10401
rect 8945 10375 8951 10401
rect 9585 10375 9591 10401
rect 9617 10375 9623 10401
rect 10649 10375 10655 10401
rect 10681 10375 10687 10401
rect 14569 10375 14575 10401
rect 14601 10375 14607 10401
rect 18825 10375 18831 10401
rect 18857 10375 18863 10401
rect 8583 10369 8609 10375
rect 6679 10345 6705 10351
rect 6057 10319 6063 10345
rect 6089 10319 6095 10345
rect 6679 10313 6705 10319
rect 6847 10345 6873 10351
rect 6847 10313 6873 10319
rect 8471 10345 8497 10351
rect 14127 10345 14153 10351
rect 9193 10319 9199 10345
rect 9225 10319 9231 10345
rect 9529 10319 9535 10345
rect 9561 10319 9567 10345
rect 12553 10319 12559 10345
rect 12585 10319 12591 10345
rect 8471 10313 8497 10319
rect 14127 10313 14153 10319
rect 14239 10345 14265 10351
rect 14239 10313 14265 10319
rect 14295 10345 14321 10351
rect 14961 10319 14967 10345
rect 14993 10319 14999 10345
rect 14295 10313 14321 10319
rect 6791 10289 6817 10295
rect 6791 10257 6817 10263
rect 7407 10289 7433 10295
rect 7407 10257 7433 10263
rect 7519 10289 7545 10295
rect 7519 10257 7545 10263
rect 672 10205 20328 10222
rect 672 10179 9919 10205
rect 9945 10179 9971 10205
rect 9997 10179 10023 10205
rect 10049 10179 20328 10205
rect 672 10162 20328 10179
rect 7575 10121 7601 10127
rect 7575 10089 7601 10095
rect 6343 10065 6369 10071
rect 6343 10033 6369 10039
rect 6791 10065 6817 10071
rect 6791 10033 6817 10039
rect 6903 10065 6929 10071
rect 6903 10033 6929 10039
rect 7127 10065 7153 10071
rect 7127 10033 7153 10039
rect 7855 10065 7881 10071
rect 7855 10033 7881 10039
rect 7911 10065 7937 10071
rect 7911 10033 7937 10039
rect 8415 10065 8441 10071
rect 12161 10039 12167 10065
rect 12193 10039 12199 10065
rect 14345 10039 14351 10065
rect 14377 10039 14383 10065
rect 8415 10033 8441 10039
rect 6735 10009 6761 10015
rect 6735 9977 6761 9983
rect 7183 10009 7209 10015
rect 7183 9977 7209 9983
rect 7463 10009 7489 10015
rect 7463 9977 7489 9983
rect 7631 10009 7657 10015
rect 7631 9977 7657 9983
rect 8023 10009 8049 10015
rect 8185 9983 8191 10009
rect 8217 9983 8223 10009
rect 11321 9983 11327 10009
rect 11353 9983 11359 10009
rect 12329 9983 12335 10009
rect 12361 9983 12367 10009
rect 12609 9983 12615 10009
rect 12641 9983 12647 10009
rect 18825 9983 18831 10009
rect 18857 9983 18863 10009
rect 8023 9977 8049 9983
rect 6567 9953 6593 9959
rect 8801 9927 8807 9953
rect 8833 9927 8839 9953
rect 6567 9921 6593 9927
rect 7127 9897 7153 9903
rect 7127 9865 7153 9871
rect 12279 9897 12305 9903
rect 12279 9865 12305 9871
rect 20007 9897 20033 9903
rect 20007 9865 20033 9871
rect 672 9813 20328 9830
rect 672 9787 2239 9813
rect 2265 9787 2291 9813
rect 2317 9787 2343 9813
rect 2369 9787 17599 9813
rect 17625 9787 17651 9813
rect 17677 9787 17703 9813
rect 17729 9787 20328 9813
rect 672 9770 20328 9787
rect 8639 9729 8665 9735
rect 8639 9697 8665 9703
rect 10991 9673 11017 9679
rect 7121 9647 7127 9673
rect 7153 9647 7159 9673
rect 8185 9647 8191 9673
rect 8217 9647 8223 9673
rect 13001 9647 13007 9673
rect 13033 9647 13039 9673
rect 13617 9647 13623 9673
rect 13649 9647 13655 9673
rect 10991 9641 11017 9647
rect 10431 9617 10457 9623
rect 6729 9591 6735 9617
rect 6761 9591 6767 9617
rect 9529 9591 9535 9617
rect 9561 9591 9567 9617
rect 9865 9591 9871 9617
rect 9897 9591 9903 9617
rect 10431 9585 10457 9591
rect 11159 9617 11185 9623
rect 11159 9585 11185 9591
rect 11383 9617 11409 9623
rect 14127 9617 14153 9623
rect 11601 9591 11607 9617
rect 11633 9591 11639 9617
rect 13225 9591 13231 9617
rect 13257 9591 13263 9617
rect 13449 9591 13455 9617
rect 13481 9591 13487 9617
rect 11383 9585 11409 9591
rect 14127 9585 14153 9591
rect 14519 9617 14545 9623
rect 14519 9585 14545 9591
rect 14799 9617 14825 9623
rect 14799 9585 14825 9591
rect 8583 9561 8609 9567
rect 10655 9561 10681 9567
rect 14295 9561 14321 9567
rect 9193 9535 9199 9561
rect 9225 9535 9231 9561
rect 9417 9535 9423 9561
rect 9449 9535 9455 9561
rect 10817 9535 10823 9561
rect 10849 9535 10855 9561
rect 11881 9535 11887 9561
rect 11913 9535 11919 9561
rect 12385 9535 12391 9561
rect 12417 9535 12423 9561
rect 8583 9529 8609 9535
rect 10655 9529 10681 9535
rect 14295 9529 14321 9535
rect 14687 9561 14713 9567
rect 14687 9529 14713 9535
rect 14911 9561 14937 9567
rect 14911 9529 14937 9535
rect 14967 9561 14993 9567
rect 14967 9529 14993 9535
rect 15135 9561 15161 9567
rect 15135 9529 15161 9535
rect 15303 9561 15329 9567
rect 15303 9529 15329 9535
rect 8415 9505 8441 9511
rect 8415 9473 8441 9479
rect 8695 9505 8721 9511
rect 8695 9473 8721 9479
rect 8807 9505 8833 9511
rect 10095 9505 10121 9511
rect 9025 9479 9031 9505
rect 9057 9479 9063 9505
rect 9753 9479 9759 9505
rect 9785 9479 9791 9505
rect 8807 9473 8833 9479
rect 10095 9473 10121 9479
rect 10151 9505 10177 9511
rect 10151 9473 10177 9479
rect 10207 9505 10233 9511
rect 10207 9473 10233 9479
rect 13847 9505 13873 9511
rect 14239 9505 14265 9511
rect 14009 9479 14015 9505
rect 14041 9479 14047 9505
rect 13847 9473 13873 9479
rect 14239 9473 14265 9479
rect 14631 9505 14657 9511
rect 14631 9473 14657 9479
rect 15191 9505 15217 9511
rect 15191 9473 15217 9479
rect 672 9421 20328 9438
rect 672 9395 9919 9421
rect 9945 9395 9971 9421
rect 9997 9395 10023 9421
rect 10049 9395 20328 9421
rect 672 9378 20328 9395
rect 7015 9337 7041 9343
rect 7015 9305 7041 9311
rect 8247 9337 8273 9343
rect 8247 9305 8273 9311
rect 8919 9337 8945 9343
rect 8919 9305 8945 9311
rect 10879 9337 10905 9343
rect 10879 9305 10905 9311
rect 12055 9337 12081 9343
rect 12055 9305 12081 9311
rect 14295 9337 14321 9343
rect 14295 9305 14321 9311
rect 8409 9255 8415 9281
rect 8441 9255 8447 9281
rect 8745 9255 8751 9281
rect 8777 9255 8783 9281
rect 9529 9255 9535 9281
rect 9561 9255 9567 9281
rect 7127 9225 7153 9231
rect 6841 9199 6847 9225
rect 6873 9199 6879 9225
rect 7127 9193 7153 9199
rect 9087 9225 9113 9231
rect 9087 9193 9113 9199
rect 9143 9225 9169 9231
rect 10599 9225 10625 9231
rect 11327 9225 11353 9231
rect 12111 9225 12137 9231
rect 9305 9199 9311 9225
rect 9337 9199 9343 9225
rect 9865 9199 9871 9225
rect 9897 9199 9903 9225
rect 10313 9199 10319 9225
rect 10345 9199 10351 9225
rect 10761 9199 10767 9225
rect 10793 9199 10799 9225
rect 11993 9199 11999 9225
rect 12025 9199 12031 9225
rect 14065 9199 14071 9225
rect 14097 9199 14103 9225
rect 9143 9193 9169 9199
rect 10599 9193 10625 9199
rect 11327 9193 11353 9199
rect 12111 9193 12137 9199
rect 7071 9169 7097 9175
rect 10431 9169 10457 9175
rect 9361 9143 9367 9169
rect 9393 9143 9399 9169
rect 7071 9137 7097 9143
rect 10431 9137 10457 9143
rect 11047 9169 11073 9175
rect 12609 9143 12615 9169
rect 12641 9143 12647 9169
rect 13673 9143 13679 9169
rect 13705 9143 13711 9169
rect 11047 9137 11073 9143
rect 10487 9113 10513 9119
rect 10487 9081 10513 9087
rect 10935 9113 10961 9119
rect 10935 9081 10961 9087
rect 672 9029 20328 9046
rect 672 9003 2239 9029
rect 2265 9003 2291 9029
rect 2317 9003 2343 9029
rect 2369 9003 17599 9029
rect 17625 9003 17651 9029
rect 17677 9003 17703 9029
rect 17729 9003 20328 9029
rect 672 8986 20328 9003
rect 6847 8945 6873 8951
rect 6847 8913 6873 8919
rect 12391 8945 12417 8951
rect 12391 8913 12417 8919
rect 967 8889 993 8895
rect 8751 8889 8777 8895
rect 7457 8863 7463 8889
rect 7489 8863 7495 8889
rect 8521 8863 8527 8889
rect 8553 8863 8559 8889
rect 967 8857 993 8863
rect 8751 8857 8777 8863
rect 9479 8889 9505 8895
rect 12727 8889 12753 8895
rect 11041 8863 11047 8889
rect 11073 8863 11079 8889
rect 12105 8863 12111 8889
rect 12137 8863 12143 8889
rect 9479 8857 9505 8863
rect 12727 8857 12753 8863
rect 20007 8889 20033 8895
rect 20007 8857 20033 8863
rect 9143 8833 9169 8839
rect 12279 8833 12305 8839
rect 2137 8807 2143 8833
rect 2169 8807 2175 8833
rect 7065 8807 7071 8833
rect 7097 8807 7103 8833
rect 9697 8807 9703 8833
rect 9729 8807 9735 8833
rect 10033 8807 10039 8833
rect 10065 8807 10071 8833
rect 10705 8807 10711 8833
rect 10737 8807 10743 8833
rect 9143 8801 9169 8807
rect 12279 8801 12305 8807
rect 12839 8833 12865 8839
rect 12839 8801 12865 8807
rect 13175 8833 13201 8839
rect 13175 8801 13201 8807
rect 13343 8833 13369 8839
rect 13343 8801 13369 8807
rect 13679 8833 13705 8839
rect 13679 8801 13705 8807
rect 14687 8833 14713 8839
rect 18825 8807 18831 8833
rect 18857 8807 18863 8833
rect 14687 8801 14713 8807
rect 6511 8777 6537 8783
rect 6511 8745 6537 8751
rect 6791 8777 6817 8783
rect 6791 8745 6817 8751
rect 6847 8777 6873 8783
rect 13231 8777 13257 8783
rect 9305 8751 9311 8777
rect 9337 8751 9343 8777
rect 9921 8751 9927 8777
rect 9953 8751 9959 8777
rect 6847 8745 6873 8751
rect 13231 8745 13257 8751
rect 14631 8777 14657 8783
rect 14631 8745 14657 8751
rect 14519 8721 14545 8727
rect 12553 8695 12559 8721
rect 12585 8695 12591 8721
rect 13001 8695 13007 8721
rect 13033 8695 13039 8721
rect 14519 8689 14545 8695
rect 672 8637 20328 8654
rect 672 8611 9919 8637
rect 9945 8611 9971 8637
rect 9997 8611 10023 8637
rect 10049 8611 20328 8637
rect 672 8594 20328 8611
rect 11047 8553 11073 8559
rect 11047 8521 11073 8527
rect 11159 8553 11185 8559
rect 11775 8553 11801 8559
rect 11601 8527 11607 8553
rect 11633 8527 11639 8553
rect 11159 8521 11185 8527
rect 11775 8521 11801 8527
rect 9087 8497 9113 8503
rect 6673 8471 6679 8497
rect 6705 8471 6711 8497
rect 9087 8465 9113 8471
rect 9143 8497 9169 8503
rect 9143 8465 9169 8471
rect 9255 8497 9281 8503
rect 9255 8465 9281 8471
rect 9423 8497 9449 8503
rect 9423 8465 9449 8471
rect 9479 8497 9505 8503
rect 10655 8497 10681 8503
rect 9809 8471 9815 8497
rect 9841 8471 9847 8497
rect 9479 8465 9505 8471
rect 10655 8465 10681 8471
rect 11215 8497 11241 8503
rect 11937 8471 11943 8497
rect 11969 8471 11975 8497
rect 11215 8465 11241 8471
rect 7295 8441 7321 8447
rect 10767 8441 10793 8447
rect 12335 8441 12361 8447
rect 15415 8441 15441 8447
rect 7065 8415 7071 8441
rect 7097 8415 7103 8441
rect 9921 8415 9927 8441
rect 9953 8415 9959 8441
rect 12049 8415 12055 8441
rect 12081 8415 12087 8441
rect 13729 8415 13735 8441
rect 13761 8415 13767 8441
rect 7295 8409 7321 8415
rect 10767 8409 10793 8415
rect 12335 8409 12361 8415
rect 15415 8409 15441 8415
rect 5609 8359 5615 8385
rect 5641 8359 5647 8385
rect 14121 8359 14127 8385
rect 14153 8359 14159 8385
rect 15185 8359 15191 8385
rect 15217 8359 15223 8385
rect 9423 8329 9449 8335
rect 9423 8297 9449 8303
rect 10935 8329 10961 8335
rect 10935 8297 10961 8303
rect 672 8245 20328 8262
rect 672 8219 2239 8245
rect 2265 8219 2291 8245
rect 2317 8219 2343 8245
rect 2369 8219 17599 8245
rect 17625 8219 17651 8245
rect 17677 8219 17703 8245
rect 17729 8219 20328 8245
rect 672 8202 20328 8219
rect 8807 8161 8833 8167
rect 8807 8129 8833 8135
rect 14071 8161 14097 8167
rect 14071 8129 14097 8135
rect 9871 8105 9897 8111
rect 9871 8073 9897 8079
rect 20007 8105 20033 8111
rect 20007 8073 20033 8079
rect 9759 8049 9785 8055
rect 8969 8023 8975 8049
rect 9001 8023 9007 8049
rect 9759 8017 9785 8023
rect 9983 8049 10009 8055
rect 10263 8049 10289 8055
rect 10089 8023 10095 8049
rect 10121 8023 10127 8049
rect 12721 8023 12727 8049
rect 12753 8023 12759 8049
rect 13057 8023 13063 8049
rect 13089 8023 13095 8049
rect 18825 8023 18831 8049
rect 18857 8023 18863 8049
rect 9983 8017 10009 8023
rect 10263 8017 10289 8023
rect 13511 7993 13537 7999
rect 14071 7993 14097 7999
rect 13511 7961 13537 7967
rect 14015 7965 14041 7971
rect 8863 7937 8889 7943
rect 12839 7937 12865 7943
rect 10033 7911 10039 7937
rect 10065 7911 10071 7937
rect 8863 7905 8889 7911
rect 12839 7905 12865 7911
rect 12895 7937 12921 7943
rect 12895 7905 12921 7911
rect 12951 7937 12977 7943
rect 12951 7905 12977 7911
rect 13455 7937 13481 7943
rect 14071 7961 14097 7967
rect 14015 7933 14041 7939
rect 13455 7905 13481 7911
rect 672 7853 20328 7870
rect 672 7827 9919 7853
rect 9945 7827 9971 7853
rect 9997 7827 10023 7853
rect 10049 7827 20328 7853
rect 672 7810 20328 7827
rect 10991 7769 11017 7775
rect 10991 7737 11017 7743
rect 14295 7769 14321 7775
rect 14295 7737 14321 7743
rect 8303 7713 8329 7719
rect 8303 7681 8329 7687
rect 8359 7713 8385 7719
rect 8359 7681 8385 7687
rect 11047 7713 11073 7719
rect 13001 7687 13007 7713
rect 13033 7687 13039 7713
rect 11047 7681 11073 7687
rect 8471 7657 8497 7663
rect 8471 7625 8497 7631
rect 8863 7657 8889 7663
rect 8863 7625 8889 7631
rect 8919 7657 8945 7663
rect 8919 7625 8945 7631
rect 9031 7657 9057 7663
rect 9031 7625 9057 7631
rect 9199 7657 9225 7663
rect 9199 7625 9225 7631
rect 9367 7657 9393 7663
rect 9367 7625 9393 7631
rect 9479 7657 9505 7663
rect 10873 7631 10879 7657
rect 10905 7631 10911 7657
rect 12665 7631 12671 7657
rect 12697 7631 12703 7657
rect 9479 7625 9505 7631
rect 9087 7601 9113 7607
rect 9087 7569 9113 7575
rect 9311 7601 9337 7607
rect 14065 7575 14071 7601
rect 14097 7575 14103 7601
rect 9311 7569 9337 7575
rect 672 7461 20328 7478
rect 672 7435 2239 7461
rect 2265 7435 2291 7461
rect 2317 7435 2343 7461
rect 2369 7435 17599 7461
rect 17625 7435 17651 7461
rect 17677 7435 17703 7461
rect 17729 7435 20328 7461
rect 672 7418 20328 7435
rect 13623 7321 13649 7327
rect 7905 7295 7911 7321
rect 7937 7295 7943 7321
rect 8969 7295 8975 7321
rect 9001 7295 9007 7321
rect 13337 7295 13343 7321
rect 13369 7295 13375 7321
rect 13623 7289 13649 7295
rect 9199 7265 9225 7271
rect 7569 7239 7575 7265
rect 7601 7239 7607 7265
rect 9199 7233 9225 7239
rect 10039 7265 10065 7271
rect 10039 7233 10065 7239
rect 10151 7265 10177 7271
rect 10151 7233 10177 7239
rect 10375 7265 10401 7271
rect 10375 7233 10401 7239
rect 10711 7265 10737 7271
rect 10711 7233 10737 7239
rect 10879 7265 10905 7271
rect 11937 7239 11943 7265
rect 11969 7239 11975 7265
rect 10879 7233 10905 7239
rect 12273 7183 12279 7209
rect 12305 7183 12311 7209
rect 10207 7153 10233 7159
rect 10207 7121 10233 7127
rect 10823 7153 10849 7159
rect 10823 7121 10849 7127
rect 672 7069 20328 7086
rect 672 7043 9919 7069
rect 9945 7043 9971 7069
rect 9997 7043 10023 7069
rect 10049 7043 20328 7069
rect 672 7026 20328 7043
rect 9591 6985 9617 6991
rect 9591 6953 9617 6959
rect 12671 6985 12697 6991
rect 12671 6953 12697 6959
rect 12727 6985 12753 6991
rect 12727 6953 12753 6959
rect 12951 6929 12977 6935
rect 10145 6903 10151 6929
rect 10177 6903 10183 6929
rect 12951 6897 12977 6903
rect 9753 6847 9759 6873
rect 9785 6847 9791 6873
rect 13113 6847 13119 6873
rect 13145 6847 13151 6873
rect 13007 6817 13033 6823
rect 11209 6791 11215 6817
rect 11241 6791 11247 6817
rect 13007 6785 13033 6791
rect 12783 6761 12809 6767
rect 12783 6729 12809 6735
rect 672 6677 20328 6694
rect 672 6651 2239 6677
rect 2265 6651 2291 6677
rect 2317 6651 2343 6677
rect 2369 6651 17599 6677
rect 17625 6651 17651 6677
rect 17677 6651 17703 6677
rect 17729 6651 20328 6677
rect 672 6634 20328 6651
rect 9143 6537 9169 6543
rect 7849 6511 7855 6537
rect 7881 6511 7887 6537
rect 8913 6511 8919 6537
rect 8945 6511 8951 6537
rect 9143 6505 9169 6511
rect 7513 6455 7519 6481
rect 7545 6455 7551 6481
rect 672 6285 20328 6302
rect 672 6259 9919 6285
rect 9945 6259 9971 6285
rect 9997 6259 10023 6285
rect 10049 6259 20328 6285
rect 672 6242 20328 6259
rect 9535 6201 9561 6207
rect 9535 6169 9561 6175
rect 10089 6119 10095 6145
rect 10121 6119 10127 6145
rect 9697 6063 9703 6089
rect 9729 6063 9735 6089
rect 11153 6007 11159 6033
rect 11185 6007 11191 6033
rect 672 5893 20328 5910
rect 672 5867 2239 5893
rect 2265 5867 2291 5893
rect 2317 5867 2343 5893
rect 2369 5867 17599 5893
rect 17625 5867 17651 5893
rect 17677 5867 17703 5893
rect 17729 5867 20328 5893
rect 672 5850 20328 5867
rect 672 5501 20328 5518
rect 672 5475 9919 5501
rect 9945 5475 9971 5501
rect 9997 5475 10023 5501
rect 10049 5475 20328 5501
rect 672 5458 20328 5475
rect 672 5109 20328 5126
rect 672 5083 2239 5109
rect 2265 5083 2291 5109
rect 2317 5083 2343 5109
rect 2369 5083 17599 5109
rect 17625 5083 17651 5109
rect 17677 5083 17703 5109
rect 17729 5083 20328 5109
rect 672 5066 20328 5083
rect 672 4717 20328 4734
rect 672 4691 9919 4717
rect 9945 4691 9971 4717
rect 9997 4691 10023 4717
rect 10049 4691 20328 4717
rect 672 4674 20328 4691
rect 672 4325 20328 4342
rect 672 4299 2239 4325
rect 2265 4299 2291 4325
rect 2317 4299 2343 4325
rect 2369 4299 17599 4325
rect 17625 4299 17651 4325
rect 17677 4299 17703 4325
rect 17729 4299 20328 4325
rect 672 4282 20328 4299
rect 672 3933 20328 3950
rect 672 3907 9919 3933
rect 9945 3907 9971 3933
rect 9997 3907 10023 3933
rect 10049 3907 20328 3933
rect 672 3890 20328 3907
rect 672 3541 20328 3558
rect 672 3515 2239 3541
rect 2265 3515 2291 3541
rect 2317 3515 2343 3541
rect 2369 3515 17599 3541
rect 17625 3515 17651 3541
rect 17677 3515 17703 3541
rect 17729 3515 20328 3541
rect 672 3498 20328 3515
rect 672 3149 20328 3166
rect 672 3123 9919 3149
rect 9945 3123 9971 3149
rect 9997 3123 10023 3149
rect 10049 3123 20328 3149
rect 672 3106 20328 3123
rect 672 2757 20328 2774
rect 672 2731 2239 2757
rect 2265 2731 2291 2757
rect 2317 2731 2343 2757
rect 2369 2731 17599 2757
rect 17625 2731 17651 2757
rect 17677 2731 17703 2757
rect 17729 2731 20328 2757
rect 672 2714 20328 2731
rect 672 2365 20328 2382
rect 672 2339 9919 2365
rect 9945 2339 9971 2365
rect 9997 2339 10023 2365
rect 10049 2339 20328 2365
rect 672 2322 20328 2339
rect 8913 2143 8919 2169
rect 8945 2143 8951 2169
rect 11097 2143 11103 2169
rect 11129 2143 11135 2169
rect 9367 2057 9393 2063
rect 9367 2025 9393 2031
rect 11383 2057 11409 2063
rect 11383 2025 11409 2031
rect 672 1973 20328 1990
rect 672 1947 2239 1973
rect 2265 1947 2291 1973
rect 2317 1947 2343 1973
rect 2369 1947 17599 1973
rect 17625 1947 17651 1973
rect 17677 1947 17703 1973
rect 17729 1947 20328 1973
rect 672 1930 20328 1947
rect 9311 1833 9337 1839
rect 12777 1807 12783 1833
rect 12809 1807 12815 1833
rect 9311 1801 9337 1807
rect 8969 1751 8975 1777
rect 9001 1751 9007 1777
rect 10705 1751 10711 1777
rect 10737 1751 10743 1777
rect 13673 1751 13679 1777
rect 13705 1751 13711 1777
rect 11215 1665 11241 1671
rect 11215 1633 11241 1639
rect 672 1581 20328 1598
rect 672 1555 9919 1581
rect 9945 1555 9971 1581
rect 9997 1555 10023 1581
rect 10049 1555 20328 1581
rect 672 1538 20328 1555
<< via1 >>
rect 2239 19195 2265 19221
rect 2291 19195 2317 19221
rect 2343 19195 2369 19221
rect 17599 19195 17625 19221
rect 17651 19195 17677 19221
rect 17703 19195 17729 19221
rect 7687 19111 7713 19137
rect 9311 19111 9337 19137
rect 11215 19111 11241 19137
rect 12783 19111 12809 19137
rect 7967 18999 7993 19025
rect 8975 18999 9001 19025
rect 10879 18999 10905 19025
rect 12279 18999 12305 19025
rect 9919 18803 9945 18829
rect 9971 18803 9997 18829
rect 10023 18803 10049 18829
rect 9367 18719 9393 18745
rect 11047 18719 11073 18745
rect 8863 18607 8889 18633
rect 10599 18607 10625 18633
rect 2239 18411 2265 18437
rect 2291 18411 2317 18437
rect 2343 18411 2369 18437
rect 17599 18411 17625 18437
rect 17651 18411 17677 18437
rect 17703 18411 17729 18437
rect 9031 18327 9057 18353
rect 8527 18215 8553 18241
rect 9919 18019 9945 18045
rect 9971 18019 9997 18045
rect 10023 18019 10049 18045
rect 2239 17627 2265 17653
rect 2291 17627 2317 17653
rect 2343 17627 2369 17653
rect 17599 17627 17625 17653
rect 17651 17627 17677 17653
rect 17703 17627 17729 17653
rect 9919 17235 9945 17261
rect 9971 17235 9997 17261
rect 10023 17235 10049 17261
rect 2239 16843 2265 16869
rect 2291 16843 2317 16869
rect 2343 16843 2369 16869
rect 17599 16843 17625 16869
rect 17651 16843 17677 16869
rect 17703 16843 17729 16869
rect 9919 16451 9945 16477
rect 9971 16451 9997 16477
rect 10023 16451 10049 16477
rect 2239 16059 2265 16085
rect 2291 16059 2317 16085
rect 2343 16059 2369 16085
rect 17599 16059 17625 16085
rect 17651 16059 17677 16085
rect 17703 16059 17729 16085
rect 9919 15667 9945 15693
rect 9971 15667 9997 15693
rect 10023 15667 10049 15693
rect 2239 15275 2265 15301
rect 2291 15275 2317 15301
rect 2343 15275 2369 15301
rect 17599 15275 17625 15301
rect 17651 15275 17677 15301
rect 17703 15275 17729 15301
rect 9919 14883 9945 14909
rect 9971 14883 9997 14909
rect 10023 14883 10049 14909
rect 2239 14491 2265 14517
rect 2291 14491 2317 14517
rect 2343 14491 2369 14517
rect 17599 14491 17625 14517
rect 17651 14491 17677 14517
rect 17703 14491 17729 14517
rect 9919 14099 9945 14125
rect 9971 14099 9997 14125
rect 10023 14099 10049 14125
rect 8695 14015 8721 14041
rect 8863 14015 8889 14041
rect 9143 13903 9169 13929
rect 9535 13847 9561 13873
rect 10599 13847 10625 13873
rect 10879 13847 10905 13873
rect 12391 13847 12417 13873
rect 2239 13707 2265 13733
rect 2291 13707 2317 13733
rect 2343 13707 2369 13733
rect 17599 13707 17625 13733
rect 17651 13707 17677 13733
rect 17703 13707 17729 13733
rect 7351 13567 7377 13593
rect 12223 13567 12249 13593
rect 13847 13567 13873 13593
rect 20007 13567 20033 13593
rect 8807 13511 8833 13537
rect 9087 13511 9113 13537
rect 10823 13511 10849 13537
rect 12391 13511 12417 13537
rect 18943 13511 18969 13537
rect 8415 13455 8441 13481
rect 8975 13455 9001 13481
rect 9535 13455 9561 13481
rect 9703 13455 9729 13481
rect 11159 13455 11185 13481
rect 12783 13455 12809 13481
rect 14071 13455 14097 13481
rect 9367 13399 9393 13425
rect 9919 13315 9945 13341
rect 9971 13315 9997 13341
rect 10023 13315 10049 13341
rect 9703 13231 9729 13257
rect 10375 13231 10401 13257
rect 12279 13231 12305 13257
rect 14295 13231 14321 13257
rect 11103 13175 11129 13201
rect 11719 13175 11745 13201
rect 12167 13175 12193 13201
rect 12223 13175 12249 13201
rect 6959 13119 6985 13145
rect 8695 13119 8721 13145
rect 8807 13119 8833 13145
rect 8919 13119 8945 13145
rect 9031 13119 9057 13145
rect 10263 13119 10289 13145
rect 10431 13119 10457 13145
rect 11943 13119 11969 13145
rect 12335 13119 12361 13145
rect 12671 13119 12697 13145
rect 18831 13119 18857 13145
rect 7351 13063 7377 13089
rect 8415 13063 8441 13089
rect 8751 13063 8777 13089
rect 9255 13063 9281 13089
rect 9423 13063 9449 13089
rect 13007 13063 13033 13089
rect 14071 13063 14097 13089
rect 19951 13063 19977 13089
rect 9535 13007 9561 13033
rect 10991 13007 11017 13033
rect 11159 13007 11185 13033
rect 11663 13007 11689 13033
rect 2239 12923 2265 12949
rect 2291 12923 2317 12949
rect 2343 12923 2369 12949
rect 17599 12923 17625 12949
rect 17651 12923 17677 12949
rect 17703 12923 17729 12949
rect 7855 12839 7881 12865
rect 11663 12839 11689 12865
rect 12335 12839 12361 12865
rect 13679 12839 13705 12865
rect 10039 12783 10065 12809
rect 11215 12783 11241 12809
rect 12839 12783 12865 12809
rect 13511 12783 13537 12809
rect 13735 12783 13761 12809
rect 8919 12727 8945 12753
rect 9031 12727 9057 12753
rect 10095 12727 10121 12753
rect 10263 12727 10289 12753
rect 10655 12727 10681 12753
rect 10767 12727 10793 12753
rect 10935 12727 10961 12753
rect 11159 12727 11185 12753
rect 11607 12727 11633 12753
rect 12391 12727 12417 12753
rect 12783 12727 12809 12753
rect 13455 12727 13481 12753
rect 7911 12671 7937 12697
rect 8583 12671 8609 12697
rect 8695 12671 8721 12697
rect 9143 12671 9169 12697
rect 9199 12671 9225 12697
rect 11327 12671 11353 12697
rect 11439 12671 11465 12697
rect 12503 12671 12529 12697
rect 12671 12671 12697 12697
rect 8527 12615 8553 12641
rect 8639 12615 8665 12641
rect 9983 12615 10009 12641
rect 10599 12615 10625 12641
rect 10879 12615 10905 12641
rect 9919 12531 9945 12557
rect 9971 12531 9997 12557
rect 10023 12531 10049 12557
rect 10039 12391 10065 12417
rect 9647 12335 9673 12361
rect 11327 12335 11353 12361
rect 11103 12279 11129 12305
rect 2239 12139 2265 12165
rect 2291 12139 2317 12165
rect 2343 12139 2369 12165
rect 17599 12139 17625 12165
rect 17651 12139 17677 12165
rect 17703 12139 17729 12165
rect 967 11999 993 12025
rect 10823 11999 10849 12025
rect 20007 11999 20033 12025
rect 2143 11943 2169 11969
rect 11047 11943 11073 11969
rect 13063 11943 13089 11969
rect 18831 11943 18857 11969
rect 7463 11887 7489 11913
rect 9143 11887 9169 11913
rect 9311 11887 9337 11913
rect 10823 11887 10849 11913
rect 12671 11887 12697 11913
rect 12727 11887 12753 11913
rect 12839 11887 12865 11913
rect 12951 11887 12977 11913
rect 13231 11887 13257 11913
rect 7631 11831 7657 11857
rect 10655 11831 10681 11857
rect 10767 11831 10793 11857
rect 13007 11831 13033 11857
rect 9919 11747 9945 11773
rect 9971 11747 9997 11773
rect 10023 11747 10049 11773
rect 9759 11663 9785 11689
rect 9143 11607 9169 11633
rect 13007 11607 13033 11633
rect 2143 11551 2169 11577
rect 7407 11551 7433 11577
rect 7687 11551 7713 11577
rect 7743 11551 7769 11577
rect 7855 11551 7881 11577
rect 7967 11551 7993 11577
rect 9087 11551 9113 11577
rect 9647 11551 9673 11577
rect 12615 11551 12641 11577
rect 14295 11551 14321 11577
rect 18943 11551 18969 11577
rect 6007 11495 6033 11521
rect 7071 11495 7097 11521
rect 7799 11495 7825 11521
rect 8191 11495 8217 11521
rect 14071 11495 14097 11521
rect 14631 11495 14657 11521
rect 15695 11495 15721 11521
rect 15919 11495 15945 11521
rect 967 11439 993 11465
rect 9143 11439 9169 11465
rect 20007 11439 20033 11465
rect 2239 11355 2265 11381
rect 2291 11355 2317 11381
rect 2343 11355 2369 11381
rect 17599 11355 17625 11381
rect 17651 11355 17677 11381
rect 17703 11355 17729 11381
rect 8023 11271 8049 11297
rect 8639 11271 8665 11297
rect 13959 11271 13985 11297
rect 967 11215 993 11241
rect 6791 11215 6817 11241
rect 7127 11215 7153 11241
rect 14183 11215 14209 11241
rect 20007 11215 20033 11241
rect 2143 11159 2169 11185
rect 7743 11159 7769 11185
rect 7855 11159 7881 11185
rect 8807 11159 8833 11185
rect 8919 11159 8945 11185
rect 9031 11159 9057 11185
rect 9479 11159 9505 11185
rect 11439 11159 11465 11185
rect 12335 11159 12361 11185
rect 12615 11159 12641 11185
rect 13063 11159 13089 11185
rect 13343 11159 13369 11185
rect 18831 11159 18857 11185
rect 7183 11103 7209 11129
rect 7407 11103 7433 11129
rect 8303 11103 8329 11129
rect 8471 11103 8497 11129
rect 8751 11103 8777 11129
rect 9591 11103 9617 11129
rect 9759 11103 9785 11129
rect 10711 11103 10737 11129
rect 11551 11103 11577 11129
rect 11719 11103 11745 11129
rect 11999 11103 12025 11129
rect 12391 11103 12417 11129
rect 13007 11103 13033 11129
rect 13287 11103 13313 11129
rect 13399 11103 13425 11129
rect 13623 11103 13649 11129
rect 13791 11103 13817 11129
rect 13903 11103 13929 11129
rect 6735 11047 6761 11073
rect 7127 11047 7153 11073
rect 7295 11047 7321 11073
rect 9815 11047 9841 11073
rect 10879 11047 10905 11073
rect 11047 11047 11073 11073
rect 11215 11047 11241 11073
rect 14743 11047 14769 11073
rect 14911 11047 14937 11073
rect 9919 10963 9945 10989
rect 9971 10963 9997 10989
rect 10023 10963 10049 10989
rect 7463 10879 7489 10905
rect 7519 10879 7545 10905
rect 7687 10879 7713 10905
rect 7799 10879 7825 10905
rect 8919 10879 8945 10905
rect 9311 10879 9337 10905
rect 10543 10879 10569 10905
rect 13399 10879 13425 10905
rect 13511 10879 13537 10905
rect 6679 10823 6705 10849
rect 7295 10823 7321 10849
rect 7071 10767 7097 10793
rect 7407 10767 7433 10793
rect 7855 10767 7881 10793
rect 9087 10767 9113 10793
rect 9255 10767 9281 10793
rect 9815 10767 9841 10793
rect 10711 10767 10737 10793
rect 11159 10767 11185 10793
rect 11495 10767 11521 10793
rect 13567 10767 13593 10793
rect 14071 10767 14097 10793
rect 5615 10711 5641 10737
rect 8079 10711 8105 10737
rect 9591 10711 9617 10737
rect 10375 10711 10401 10737
rect 11103 10711 11129 10737
rect 11607 10711 11633 10737
rect 11999 10711 12025 10737
rect 12111 10711 12137 10737
rect 12335 10711 12361 10737
rect 14407 10711 14433 10737
rect 15471 10711 15497 10737
rect 15695 10711 15721 10737
rect 12279 10655 12305 10681
rect 2239 10571 2265 10597
rect 2291 10571 2317 10597
rect 2343 10571 2369 10597
rect 17599 10571 17625 10597
rect 17651 10571 17677 10597
rect 17703 10571 17729 10597
rect 7351 10487 7377 10513
rect 967 10431 993 10457
rect 4999 10431 5025 10457
rect 7183 10431 7209 10457
rect 8527 10431 8553 10457
rect 9759 10431 9785 10457
rect 14015 10431 14041 10457
rect 16031 10431 16057 10457
rect 20007 10431 20033 10457
rect 2143 10375 2169 10401
rect 6455 10375 6481 10401
rect 7687 10375 7713 10401
rect 8583 10375 8609 10401
rect 8919 10375 8945 10401
rect 9591 10375 9617 10401
rect 10655 10375 10681 10401
rect 14575 10375 14601 10401
rect 18831 10375 18857 10401
rect 6063 10319 6089 10345
rect 6679 10319 6705 10345
rect 6847 10319 6873 10345
rect 8471 10319 8497 10345
rect 9199 10319 9225 10345
rect 9535 10319 9561 10345
rect 12559 10319 12585 10345
rect 14127 10319 14153 10345
rect 14239 10319 14265 10345
rect 14295 10319 14321 10345
rect 14967 10319 14993 10345
rect 6791 10263 6817 10289
rect 7407 10263 7433 10289
rect 7519 10263 7545 10289
rect 9919 10179 9945 10205
rect 9971 10179 9997 10205
rect 10023 10179 10049 10205
rect 7575 10095 7601 10121
rect 6343 10039 6369 10065
rect 6791 10039 6817 10065
rect 6903 10039 6929 10065
rect 7127 10039 7153 10065
rect 7855 10039 7881 10065
rect 7911 10039 7937 10065
rect 8415 10039 8441 10065
rect 12167 10039 12193 10065
rect 14351 10039 14377 10065
rect 6735 9983 6761 10009
rect 7183 9983 7209 10009
rect 7463 9983 7489 10009
rect 7631 9983 7657 10009
rect 8023 9983 8049 10009
rect 8191 9983 8217 10009
rect 11327 9983 11353 10009
rect 12335 9983 12361 10009
rect 12615 9983 12641 10009
rect 18831 9983 18857 10009
rect 6567 9927 6593 9953
rect 8807 9927 8833 9953
rect 7127 9871 7153 9897
rect 12279 9871 12305 9897
rect 20007 9871 20033 9897
rect 2239 9787 2265 9813
rect 2291 9787 2317 9813
rect 2343 9787 2369 9813
rect 17599 9787 17625 9813
rect 17651 9787 17677 9813
rect 17703 9787 17729 9813
rect 8639 9703 8665 9729
rect 7127 9647 7153 9673
rect 8191 9647 8217 9673
rect 10991 9647 11017 9673
rect 13007 9647 13033 9673
rect 13623 9647 13649 9673
rect 6735 9591 6761 9617
rect 9535 9591 9561 9617
rect 9871 9591 9897 9617
rect 10431 9591 10457 9617
rect 11159 9591 11185 9617
rect 11383 9591 11409 9617
rect 11607 9591 11633 9617
rect 13231 9591 13257 9617
rect 13455 9591 13481 9617
rect 14127 9591 14153 9617
rect 14519 9591 14545 9617
rect 14799 9591 14825 9617
rect 8583 9535 8609 9561
rect 9199 9535 9225 9561
rect 9423 9535 9449 9561
rect 10655 9535 10681 9561
rect 10823 9535 10849 9561
rect 11887 9535 11913 9561
rect 12391 9535 12417 9561
rect 14295 9535 14321 9561
rect 14687 9535 14713 9561
rect 14911 9535 14937 9561
rect 14967 9535 14993 9561
rect 15135 9535 15161 9561
rect 15303 9535 15329 9561
rect 8415 9479 8441 9505
rect 8695 9479 8721 9505
rect 8807 9479 8833 9505
rect 9031 9479 9057 9505
rect 9759 9479 9785 9505
rect 10095 9479 10121 9505
rect 10151 9479 10177 9505
rect 10207 9479 10233 9505
rect 13847 9479 13873 9505
rect 14015 9479 14041 9505
rect 14239 9479 14265 9505
rect 14631 9479 14657 9505
rect 15191 9479 15217 9505
rect 9919 9395 9945 9421
rect 9971 9395 9997 9421
rect 10023 9395 10049 9421
rect 7015 9311 7041 9337
rect 8247 9311 8273 9337
rect 8919 9311 8945 9337
rect 10879 9311 10905 9337
rect 12055 9311 12081 9337
rect 14295 9311 14321 9337
rect 8415 9255 8441 9281
rect 8751 9255 8777 9281
rect 9535 9255 9561 9281
rect 6847 9199 6873 9225
rect 7127 9199 7153 9225
rect 9087 9199 9113 9225
rect 9143 9199 9169 9225
rect 9311 9199 9337 9225
rect 9871 9199 9897 9225
rect 10319 9199 10345 9225
rect 10599 9199 10625 9225
rect 10767 9199 10793 9225
rect 11327 9199 11353 9225
rect 11999 9199 12025 9225
rect 12111 9199 12137 9225
rect 14071 9199 14097 9225
rect 7071 9143 7097 9169
rect 9367 9143 9393 9169
rect 10431 9143 10457 9169
rect 11047 9143 11073 9169
rect 12615 9143 12641 9169
rect 13679 9143 13705 9169
rect 10487 9087 10513 9113
rect 10935 9087 10961 9113
rect 2239 9003 2265 9029
rect 2291 9003 2317 9029
rect 2343 9003 2369 9029
rect 17599 9003 17625 9029
rect 17651 9003 17677 9029
rect 17703 9003 17729 9029
rect 6847 8919 6873 8945
rect 12391 8919 12417 8945
rect 967 8863 993 8889
rect 7463 8863 7489 8889
rect 8527 8863 8553 8889
rect 8751 8863 8777 8889
rect 9479 8863 9505 8889
rect 11047 8863 11073 8889
rect 12111 8863 12137 8889
rect 12727 8863 12753 8889
rect 20007 8863 20033 8889
rect 2143 8807 2169 8833
rect 7071 8807 7097 8833
rect 9143 8807 9169 8833
rect 9703 8807 9729 8833
rect 10039 8807 10065 8833
rect 10711 8807 10737 8833
rect 12279 8807 12305 8833
rect 12839 8807 12865 8833
rect 13175 8807 13201 8833
rect 13343 8807 13369 8833
rect 13679 8807 13705 8833
rect 14687 8807 14713 8833
rect 18831 8807 18857 8833
rect 6511 8751 6537 8777
rect 6791 8751 6817 8777
rect 6847 8751 6873 8777
rect 9311 8751 9337 8777
rect 9927 8751 9953 8777
rect 13231 8751 13257 8777
rect 14631 8751 14657 8777
rect 12559 8695 12585 8721
rect 13007 8695 13033 8721
rect 14519 8695 14545 8721
rect 9919 8611 9945 8637
rect 9971 8611 9997 8637
rect 10023 8611 10049 8637
rect 11047 8527 11073 8553
rect 11159 8527 11185 8553
rect 11607 8527 11633 8553
rect 11775 8527 11801 8553
rect 6679 8471 6705 8497
rect 9087 8471 9113 8497
rect 9143 8471 9169 8497
rect 9255 8471 9281 8497
rect 9423 8471 9449 8497
rect 9479 8471 9505 8497
rect 9815 8471 9841 8497
rect 10655 8471 10681 8497
rect 11215 8471 11241 8497
rect 11943 8471 11969 8497
rect 7071 8415 7097 8441
rect 7295 8415 7321 8441
rect 9927 8415 9953 8441
rect 10767 8415 10793 8441
rect 12055 8415 12081 8441
rect 12335 8415 12361 8441
rect 13735 8415 13761 8441
rect 15415 8415 15441 8441
rect 5615 8359 5641 8385
rect 14127 8359 14153 8385
rect 15191 8359 15217 8385
rect 9423 8303 9449 8329
rect 10935 8303 10961 8329
rect 2239 8219 2265 8245
rect 2291 8219 2317 8245
rect 2343 8219 2369 8245
rect 17599 8219 17625 8245
rect 17651 8219 17677 8245
rect 17703 8219 17729 8245
rect 8807 8135 8833 8161
rect 14071 8135 14097 8161
rect 9871 8079 9897 8105
rect 20007 8079 20033 8105
rect 8975 8023 9001 8049
rect 9759 8023 9785 8049
rect 9983 8023 10009 8049
rect 10095 8023 10121 8049
rect 10263 8023 10289 8049
rect 12727 8023 12753 8049
rect 13063 8023 13089 8049
rect 18831 8023 18857 8049
rect 13511 7967 13537 7993
rect 8863 7911 8889 7937
rect 10039 7911 10065 7937
rect 12839 7911 12865 7937
rect 12895 7911 12921 7937
rect 12951 7911 12977 7937
rect 13455 7911 13481 7937
rect 14015 7939 14041 7965
rect 14071 7967 14097 7993
rect 9919 7827 9945 7853
rect 9971 7827 9997 7853
rect 10023 7827 10049 7853
rect 10991 7743 11017 7769
rect 14295 7743 14321 7769
rect 8303 7687 8329 7713
rect 8359 7687 8385 7713
rect 11047 7687 11073 7713
rect 13007 7687 13033 7713
rect 8471 7631 8497 7657
rect 8863 7631 8889 7657
rect 8919 7631 8945 7657
rect 9031 7631 9057 7657
rect 9199 7631 9225 7657
rect 9367 7631 9393 7657
rect 9479 7631 9505 7657
rect 10879 7631 10905 7657
rect 12671 7631 12697 7657
rect 9087 7575 9113 7601
rect 9311 7575 9337 7601
rect 14071 7575 14097 7601
rect 2239 7435 2265 7461
rect 2291 7435 2317 7461
rect 2343 7435 2369 7461
rect 17599 7435 17625 7461
rect 17651 7435 17677 7461
rect 17703 7435 17729 7461
rect 7911 7295 7937 7321
rect 8975 7295 9001 7321
rect 13343 7295 13369 7321
rect 13623 7295 13649 7321
rect 7575 7239 7601 7265
rect 9199 7239 9225 7265
rect 10039 7239 10065 7265
rect 10151 7239 10177 7265
rect 10375 7239 10401 7265
rect 10711 7239 10737 7265
rect 10879 7239 10905 7265
rect 11943 7239 11969 7265
rect 12279 7183 12305 7209
rect 10207 7127 10233 7153
rect 10823 7127 10849 7153
rect 9919 7043 9945 7069
rect 9971 7043 9997 7069
rect 10023 7043 10049 7069
rect 9591 6959 9617 6985
rect 12671 6959 12697 6985
rect 12727 6959 12753 6985
rect 10151 6903 10177 6929
rect 12951 6903 12977 6929
rect 9759 6847 9785 6873
rect 13119 6847 13145 6873
rect 11215 6791 11241 6817
rect 13007 6791 13033 6817
rect 12783 6735 12809 6761
rect 2239 6651 2265 6677
rect 2291 6651 2317 6677
rect 2343 6651 2369 6677
rect 17599 6651 17625 6677
rect 17651 6651 17677 6677
rect 17703 6651 17729 6677
rect 7855 6511 7881 6537
rect 8919 6511 8945 6537
rect 9143 6511 9169 6537
rect 7519 6455 7545 6481
rect 9919 6259 9945 6285
rect 9971 6259 9997 6285
rect 10023 6259 10049 6285
rect 9535 6175 9561 6201
rect 10095 6119 10121 6145
rect 9703 6063 9729 6089
rect 11159 6007 11185 6033
rect 2239 5867 2265 5893
rect 2291 5867 2317 5893
rect 2343 5867 2369 5893
rect 17599 5867 17625 5893
rect 17651 5867 17677 5893
rect 17703 5867 17729 5893
rect 9919 5475 9945 5501
rect 9971 5475 9997 5501
rect 10023 5475 10049 5501
rect 2239 5083 2265 5109
rect 2291 5083 2317 5109
rect 2343 5083 2369 5109
rect 17599 5083 17625 5109
rect 17651 5083 17677 5109
rect 17703 5083 17729 5109
rect 9919 4691 9945 4717
rect 9971 4691 9997 4717
rect 10023 4691 10049 4717
rect 2239 4299 2265 4325
rect 2291 4299 2317 4325
rect 2343 4299 2369 4325
rect 17599 4299 17625 4325
rect 17651 4299 17677 4325
rect 17703 4299 17729 4325
rect 9919 3907 9945 3933
rect 9971 3907 9997 3933
rect 10023 3907 10049 3933
rect 2239 3515 2265 3541
rect 2291 3515 2317 3541
rect 2343 3515 2369 3541
rect 17599 3515 17625 3541
rect 17651 3515 17677 3541
rect 17703 3515 17729 3541
rect 9919 3123 9945 3149
rect 9971 3123 9997 3149
rect 10023 3123 10049 3149
rect 2239 2731 2265 2757
rect 2291 2731 2317 2757
rect 2343 2731 2369 2757
rect 17599 2731 17625 2757
rect 17651 2731 17677 2757
rect 17703 2731 17729 2757
rect 9919 2339 9945 2365
rect 9971 2339 9997 2365
rect 10023 2339 10049 2365
rect 8919 2143 8945 2169
rect 11103 2143 11129 2169
rect 9367 2031 9393 2057
rect 11383 2031 11409 2057
rect 2239 1947 2265 1973
rect 2291 1947 2317 1973
rect 2343 1947 2369 1973
rect 17599 1947 17625 1973
rect 17651 1947 17677 1973
rect 17703 1947 17729 1973
rect 9311 1807 9337 1833
rect 12783 1807 12809 1833
rect 8975 1751 9001 1777
rect 10711 1751 10737 1777
rect 13679 1751 13705 1777
rect 11215 1639 11241 1665
rect 9919 1555 9945 1581
rect 9971 1555 9997 1581
rect 10023 1555 10049 1581
<< metal2 >>
rect 8064 20600 8120 21000
rect 8400 20600 8456 21000
rect 8736 20600 8792 21000
rect 9072 20600 9128 21000
rect 10416 20600 10472 21000
rect 11088 20600 11144 21000
rect 12096 20600 12152 21000
rect 2238 19222 2370 19227
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2238 19189 2370 19194
rect 7686 19138 7714 19143
rect 7686 19091 7714 19110
rect 8078 19138 8106 20600
rect 8078 19105 8106 19110
rect 7966 19025 7994 19031
rect 7966 18999 7967 19025
rect 7993 18999 7994 19025
rect 2238 18438 2370 18443
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2238 18405 2370 18410
rect 2238 17654 2370 17659
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2238 17621 2370 17626
rect 2238 16870 2370 16875
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2238 16837 2370 16842
rect 2238 16086 2370 16091
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2238 16053 2370 16058
rect 2238 15302 2370 15307
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2238 15269 2370 15274
rect 2238 14518 2370 14523
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2238 14485 2370 14490
rect 7350 14042 7378 14047
rect 2238 13734 2370 13739
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2238 13701 2370 13706
rect 7350 13593 7378 14014
rect 7966 14042 7994 18999
rect 8414 18354 8442 20600
rect 8750 18746 8778 20600
rect 9086 19138 9114 20600
rect 9310 19138 9338 19143
rect 9086 19137 9338 19138
rect 9086 19111 9311 19137
rect 9337 19111 9338 19137
rect 9086 19110 9338 19111
rect 9310 19105 9338 19110
rect 8750 18713 8778 18718
rect 8974 19025 9002 19031
rect 8974 18999 8975 19025
rect 9001 18999 9002 19025
rect 8414 18321 8442 18326
rect 8862 18633 8890 18639
rect 8862 18607 8863 18633
rect 8889 18607 8890 18633
rect 8526 18241 8554 18247
rect 8526 18215 8527 18241
rect 8553 18215 8554 18241
rect 8526 15974 8554 18215
rect 7966 14009 7994 14014
rect 8414 15946 8554 15974
rect 8414 13594 8442 15946
rect 8694 14042 8722 14047
rect 8694 13995 8722 14014
rect 8862 14041 8890 18607
rect 8862 14015 8863 14041
rect 8889 14015 8890 14041
rect 8862 14009 8890 14015
rect 7350 13567 7351 13593
rect 7377 13567 7378 13593
rect 7350 13561 7378 13567
rect 8358 13566 8442 13594
rect 2086 13482 2114 13487
rect 966 12025 994 12031
rect 966 11999 967 12025
rect 993 11999 994 12025
rect 966 11802 994 11999
rect 966 11769 994 11774
rect 966 11466 994 11471
rect 966 11419 994 11438
rect 966 11242 994 11247
rect 966 11195 994 11214
rect 2086 10738 2114 13454
rect 8358 13370 8386 13566
rect 8806 13537 8834 13543
rect 8806 13511 8807 13537
rect 8833 13511 8834 13537
rect 8414 13482 8442 13487
rect 8806 13482 8834 13511
rect 8414 13481 8778 13482
rect 8414 13455 8415 13481
rect 8441 13455 8778 13481
rect 8414 13454 8778 13455
rect 8414 13449 8442 13454
rect 8358 13342 8442 13370
rect 6958 13145 6986 13151
rect 6958 13119 6959 13145
rect 6985 13119 6986 13145
rect 2238 12950 2370 12955
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2238 12917 2370 12922
rect 2238 12166 2370 12171
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2238 12133 2370 12138
rect 2142 11970 2170 11975
rect 2142 11923 2170 11942
rect 2142 11578 2170 11583
rect 2142 11531 2170 11550
rect 5614 11578 5642 11583
rect 2238 11382 2370 11387
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2238 11349 2370 11354
rect 2142 11186 2170 11191
rect 2142 11139 2170 11158
rect 2086 10705 2114 10710
rect 5614 11130 5642 11550
rect 6006 11522 6034 11527
rect 6006 11186 6034 11494
rect 6958 11410 6986 13119
rect 7350 13090 7378 13095
rect 7350 13043 7378 13062
rect 7854 13090 7882 13095
rect 7854 12865 7882 13062
rect 7854 12839 7855 12865
rect 7881 12839 7882 12865
rect 7854 12833 7882 12839
rect 8414 13089 8442 13342
rect 8414 13063 8415 13089
rect 8441 13063 8442 13089
rect 7910 12698 7938 12703
rect 7910 12651 7938 12670
rect 8414 12642 8442 13063
rect 8694 13145 8722 13151
rect 8694 13119 8695 13145
rect 8721 13119 8722 13145
rect 8694 12810 8722 13119
rect 8750 13089 8778 13454
rect 8806 13449 8834 13454
rect 8974 13481 9002 18999
rect 9918 18830 10050 18835
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 9918 18797 10050 18802
rect 9366 18746 9394 18751
rect 9366 18699 9394 18718
rect 10430 18746 10458 20600
rect 11102 19138 11130 20600
rect 11214 19138 11242 19143
rect 11102 19137 11242 19138
rect 11102 19111 11215 19137
rect 11241 19111 11242 19137
rect 11102 19110 11242 19111
rect 11214 19105 11242 19110
rect 12110 19138 12138 20600
rect 17598 19222 17730 19227
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17598 19189 17730 19194
rect 12110 19105 12138 19110
rect 12782 19138 12810 19143
rect 12782 19091 12810 19110
rect 10878 19026 10906 19031
rect 10878 19025 10962 19026
rect 10878 18999 10879 19025
rect 10905 18999 10962 19025
rect 10878 18998 10962 18999
rect 10878 18993 10906 18998
rect 10430 18713 10458 18718
rect 10598 18633 10626 18639
rect 10598 18607 10599 18633
rect 10625 18607 10626 18633
rect 9030 18354 9058 18359
rect 9030 18307 9058 18326
rect 9918 18046 10050 18051
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 9918 18013 10050 18018
rect 9918 17262 10050 17267
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 9918 17229 10050 17234
rect 9918 16478 10050 16483
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 9918 16445 10050 16450
rect 9918 15694 10050 15699
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 9918 15661 10050 15666
rect 9918 14910 10050 14915
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 9918 14877 10050 14882
rect 9918 14126 10050 14131
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 9918 14093 10050 14098
rect 9086 14042 9114 14047
rect 9086 13538 9114 14014
rect 9142 13929 9170 13935
rect 9142 13903 9143 13929
rect 9169 13903 9170 13929
rect 9142 13874 9170 13903
rect 9142 13841 9170 13846
rect 9366 13874 9394 13879
rect 9086 13537 9170 13538
rect 9086 13511 9087 13537
rect 9113 13511 9170 13537
rect 9086 13510 9170 13511
rect 9086 13505 9114 13510
rect 8974 13455 8975 13481
rect 9001 13455 9002 13481
rect 8974 13449 9002 13455
rect 8750 13063 8751 13089
rect 8777 13063 8778 13089
rect 8750 13057 8778 13063
rect 8806 13145 8834 13151
rect 8806 13119 8807 13145
rect 8833 13119 8834 13145
rect 8414 12609 8442 12614
rect 8526 12782 8722 12810
rect 8526 12641 8554 12782
rect 8806 12754 8834 13119
rect 8918 13146 8946 13151
rect 8974 13146 9002 13151
rect 8918 13145 8974 13146
rect 8918 13119 8919 13145
rect 8945 13119 8974 13145
rect 8918 13118 8974 13119
rect 8918 13113 8946 13118
rect 8918 12754 8946 12759
rect 8806 12753 8946 12754
rect 8806 12727 8919 12753
rect 8945 12727 8946 12753
rect 8806 12726 8946 12727
rect 8582 12698 8610 12703
rect 8582 12651 8610 12670
rect 8694 12697 8722 12703
rect 8694 12671 8695 12697
rect 8721 12671 8722 12697
rect 8526 12615 8527 12641
rect 8553 12615 8554 12641
rect 7462 11970 7490 11975
rect 7462 11913 7490 11942
rect 7462 11887 7463 11913
rect 7489 11887 7490 11913
rect 7462 11881 7490 11887
rect 7630 11857 7658 11863
rect 7630 11831 7631 11857
rect 7657 11831 7658 11857
rect 7630 11690 7658 11831
rect 8526 11802 8554 12615
rect 8638 12642 8666 12647
rect 8694 12642 8722 12671
rect 8918 12698 8946 12726
rect 8918 12665 8946 12670
rect 8694 12614 8778 12642
rect 8638 12595 8666 12614
rect 8526 11769 8554 11774
rect 7630 11662 7770 11690
rect 7406 11577 7434 11583
rect 7406 11551 7407 11577
rect 7433 11551 7434 11577
rect 7070 11522 7098 11527
rect 7070 11521 7378 11522
rect 7070 11495 7071 11521
rect 7097 11495 7378 11521
rect 7070 11494 7378 11495
rect 7070 11489 7098 11494
rect 6958 11377 6986 11382
rect 7238 11410 7266 11415
rect 6790 11242 6818 11247
rect 7126 11242 7154 11247
rect 6790 11241 7154 11242
rect 6790 11215 6791 11241
rect 6817 11215 7127 11241
rect 7153 11215 7154 11241
rect 6790 11214 7154 11215
rect 6790 11209 6818 11214
rect 7126 11209 7154 11214
rect 6006 11153 6034 11158
rect 5614 10737 5642 11102
rect 7182 11130 7210 11135
rect 7182 11083 7210 11102
rect 6734 11074 6762 11079
rect 6678 11073 6762 11074
rect 6678 11047 6735 11073
rect 6761 11047 6762 11073
rect 6678 11046 6762 11047
rect 6678 10849 6706 11046
rect 6734 11041 6762 11046
rect 7126 11073 7154 11079
rect 7126 11047 7127 11073
rect 7153 11047 7154 11073
rect 6678 10823 6679 10849
rect 6705 10823 6706 10849
rect 6678 10817 6706 10823
rect 5614 10711 5615 10737
rect 5641 10711 5642 10737
rect 5614 10705 5642 10711
rect 7070 10793 7098 10799
rect 7070 10767 7071 10793
rect 7097 10767 7098 10793
rect 2238 10598 2370 10603
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2238 10565 2370 10570
rect 966 10457 994 10463
rect 966 10431 967 10457
rect 993 10431 994 10457
rect 966 10122 994 10431
rect 4998 10458 5026 10463
rect 4998 10411 5026 10430
rect 6734 10458 6762 10463
rect 7070 10458 7098 10767
rect 7126 10626 7154 11047
rect 7238 11018 7266 11382
rect 7350 11242 7378 11494
rect 7406 11410 7434 11551
rect 7686 11578 7714 11583
rect 7686 11531 7714 11550
rect 7742 11577 7770 11662
rect 8302 11634 8330 11639
rect 7742 11551 7743 11577
rect 7769 11551 7770 11577
rect 7742 11522 7770 11551
rect 7854 11578 7882 11583
rect 7966 11578 7994 11583
rect 7854 11577 7938 11578
rect 7854 11551 7855 11577
rect 7881 11551 7938 11577
rect 7854 11550 7938 11551
rect 7854 11545 7882 11550
rect 7742 11489 7770 11494
rect 7798 11521 7826 11527
rect 7798 11495 7799 11521
rect 7825 11495 7826 11521
rect 7406 11377 7434 11382
rect 7798 11298 7826 11495
rect 7518 11270 7826 11298
rect 7350 11214 7490 11242
rect 7406 11130 7434 11135
rect 7406 11083 7434 11102
rect 7294 11074 7322 11079
rect 7294 11073 7378 11074
rect 7294 11047 7295 11073
rect 7321 11047 7378 11073
rect 7294 11046 7378 11047
rect 7294 11041 7322 11046
rect 7126 10593 7154 10598
rect 7182 10990 7266 11018
rect 7182 10458 7210 10990
rect 7350 10906 7378 11046
rect 7350 10873 7378 10878
rect 7462 10905 7490 11214
rect 7462 10879 7463 10905
rect 7489 10879 7490 10905
rect 7462 10873 7490 10879
rect 7518 10905 7546 11270
rect 7742 11186 7770 11191
rect 7518 10879 7519 10905
rect 7545 10879 7546 10905
rect 7518 10873 7546 10879
rect 7574 10962 7602 10967
rect 7294 10849 7322 10855
rect 7294 10823 7295 10849
rect 7321 10823 7322 10849
rect 7294 10514 7322 10823
rect 7406 10793 7434 10799
rect 7406 10767 7407 10793
rect 7433 10767 7434 10793
rect 7350 10514 7378 10519
rect 7070 10457 7210 10458
rect 7070 10431 7183 10457
rect 7209 10431 7210 10457
rect 7070 10430 7210 10431
rect 2142 10402 2170 10407
rect 2142 10355 2170 10374
rect 6454 10401 6482 10407
rect 6454 10375 6455 10401
rect 6481 10375 6482 10401
rect 6062 10346 6090 10351
rect 6062 10299 6090 10318
rect 6454 10094 6482 10375
rect 6678 10346 6706 10351
rect 6678 10299 6706 10318
rect 6734 10122 6762 10430
rect 7182 10425 7210 10430
rect 7238 10513 7378 10514
rect 7238 10487 7351 10513
rect 7377 10487 7378 10513
rect 7238 10486 7378 10487
rect 6846 10346 6874 10351
rect 7238 10346 7266 10486
rect 7350 10481 7378 10486
rect 7406 10514 7434 10767
rect 7406 10481 7434 10486
rect 6846 10345 7266 10346
rect 6846 10319 6847 10345
rect 6873 10319 7266 10345
rect 6846 10318 7266 10319
rect 6846 10313 6874 10318
rect 6790 10289 6818 10295
rect 6790 10263 6791 10289
rect 6817 10263 6818 10289
rect 6790 10178 6818 10263
rect 7406 10289 7434 10295
rect 7406 10263 7407 10289
rect 7433 10263 7434 10289
rect 6790 10150 6874 10178
rect 6734 10094 6818 10122
rect 966 10089 994 10094
rect 6342 10066 6706 10094
rect 6342 10065 6370 10066
rect 6342 10039 6343 10065
rect 6369 10039 6370 10065
rect 6342 10033 6370 10039
rect 6566 9954 6594 9959
rect 6510 9926 6566 9954
rect 2238 9814 2370 9819
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2238 9781 2370 9786
rect 2238 9030 2370 9035
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2238 8997 2370 9002
rect 966 8890 994 8895
rect 966 8843 994 8862
rect 2142 8834 2170 8839
rect 2142 8787 2170 8806
rect 5614 8834 5642 8839
rect 5614 8385 5642 8806
rect 6510 8778 6538 9926
rect 6566 9907 6594 9926
rect 6678 9618 6706 10066
rect 6790 10065 6818 10094
rect 6790 10039 6791 10065
rect 6817 10039 6818 10065
rect 6790 10033 6818 10039
rect 6846 10066 6874 10150
rect 6902 10066 6930 10071
rect 7126 10066 7154 10071
rect 6846 10065 6930 10066
rect 6846 10039 6903 10065
rect 6929 10039 6930 10065
rect 6846 10038 6930 10039
rect 6902 10033 6930 10038
rect 7070 10065 7154 10066
rect 7070 10039 7127 10065
rect 7153 10039 7154 10065
rect 7070 10038 7154 10039
rect 6734 10009 6762 10015
rect 6734 9983 6735 10009
rect 6761 9983 6762 10009
rect 6734 9954 6762 9983
rect 6734 9921 6762 9926
rect 7070 9898 7098 10038
rect 7126 10033 7154 10038
rect 7182 10010 7210 10015
rect 7182 9963 7210 9982
rect 7014 9870 7070 9898
rect 6734 9618 6762 9623
rect 6678 9617 6986 9618
rect 6678 9591 6735 9617
rect 6761 9591 6986 9617
rect 6678 9590 6986 9591
rect 6734 9585 6762 9590
rect 6958 9506 6986 9590
rect 6846 9225 6874 9231
rect 6846 9199 6847 9225
rect 6873 9199 6874 9225
rect 6510 8731 6538 8750
rect 6678 9170 6706 9175
rect 6678 8497 6706 9142
rect 6846 8945 6874 9199
rect 6846 8919 6847 8945
rect 6873 8919 6874 8945
rect 6846 8913 6874 8919
rect 6846 8834 6874 8839
rect 6958 8834 6986 9478
rect 7014 9337 7042 9870
rect 7070 9865 7098 9870
rect 7126 9897 7154 9903
rect 7126 9871 7127 9897
rect 7153 9871 7154 9897
rect 7126 9673 7154 9871
rect 7126 9647 7127 9673
rect 7153 9647 7154 9673
rect 7126 9641 7154 9647
rect 7014 9311 7015 9337
rect 7041 9311 7042 9337
rect 7014 9305 7042 9311
rect 7126 9225 7154 9231
rect 7126 9199 7127 9225
rect 7153 9199 7154 9225
rect 7070 9170 7098 9175
rect 7070 9123 7098 9142
rect 7070 8834 7098 8839
rect 6958 8833 7098 8834
rect 6958 8807 7071 8833
rect 7097 8807 7098 8833
rect 6958 8806 7098 8807
rect 6790 8778 6818 8783
rect 6790 8731 6818 8750
rect 6846 8777 6874 8806
rect 6846 8751 6847 8777
rect 6873 8751 6874 8777
rect 6846 8745 6874 8751
rect 6678 8471 6679 8497
rect 6705 8471 6706 8497
rect 6678 8465 6706 8471
rect 7070 8442 7098 8806
rect 7126 8722 7154 9199
rect 7406 9058 7434 10263
rect 7518 10289 7546 10295
rect 7518 10263 7519 10289
rect 7545 10263 7546 10289
rect 7462 10010 7490 10015
rect 7518 10010 7546 10263
rect 7574 10121 7602 10934
rect 7686 10906 7714 10911
rect 7742 10906 7770 11158
rect 7854 11185 7882 11191
rect 7854 11159 7855 11185
rect 7881 11159 7882 11185
rect 7798 10906 7826 10911
rect 7742 10905 7826 10906
rect 7742 10879 7799 10905
rect 7825 10879 7826 10905
rect 7742 10878 7826 10879
rect 7686 10859 7714 10878
rect 7686 10514 7714 10519
rect 7686 10401 7714 10486
rect 7686 10375 7687 10401
rect 7713 10375 7714 10401
rect 7686 10369 7714 10375
rect 7574 10095 7575 10121
rect 7601 10095 7602 10121
rect 7574 10089 7602 10095
rect 7798 10094 7826 10878
rect 7854 10794 7882 11159
rect 7910 10962 7938 11550
rect 7966 11577 8050 11578
rect 7966 11551 7967 11577
rect 7993 11551 8050 11577
rect 7966 11550 8050 11551
rect 7966 11545 7994 11550
rect 8022 11297 8050 11550
rect 8190 11521 8218 11527
rect 8190 11495 8191 11521
rect 8217 11495 8218 11521
rect 8190 11410 8218 11495
rect 8190 11377 8218 11382
rect 8022 11271 8023 11297
rect 8049 11271 8050 11297
rect 8022 11265 8050 11271
rect 8302 11186 8330 11606
rect 8638 11578 8666 11583
rect 8638 11297 8666 11550
rect 8638 11271 8639 11297
rect 8665 11271 8666 11297
rect 8638 11265 8666 11271
rect 8750 11298 8778 12614
rect 8974 12586 9002 13118
rect 9030 13145 9058 13151
rect 9030 13119 9031 13145
rect 9057 13119 9058 13145
rect 9030 12753 9058 13119
rect 9030 12727 9031 12753
rect 9057 12727 9058 12753
rect 9030 12721 9058 12727
rect 9086 12810 9114 12815
rect 8750 11265 8778 11270
rect 8862 12558 9002 12586
rect 8302 11129 8330 11158
rect 8806 11186 8834 11191
rect 8806 11139 8834 11158
rect 8302 11103 8303 11129
rect 8329 11103 8330 11129
rect 8302 11097 8330 11103
rect 8470 11129 8498 11135
rect 8470 11103 8471 11129
rect 8497 11103 8498 11129
rect 8470 11018 8498 11103
rect 8750 11129 8778 11135
rect 8750 11103 8751 11129
rect 8777 11103 8778 11129
rect 8750 11074 8778 11103
rect 8862 11074 8890 12558
rect 9086 11802 9114 12782
rect 9142 12697 9170 13510
rect 9366 13482 9394 13846
rect 9366 13425 9394 13454
rect 9534 13873 9562 13879
rect 10598 13874 10626 18607
rect 10934 15974 10962 18998
rect 12278 19025 12306 19031
rect 12278 18999 12279 19025
rect 12305 18999 12306 19025
rect 11046 18746 11074 18751
rect 11046 18699 11074 18718
rect 12278 15974 12306 18999
rect 17598 18438 17730 18443
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17598 18405 17730 18410
rect 17598 17654 17730 17659
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17598 17621 17730 17626
rect 17598 16870 17730 16875
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17598 16837 17730 16842
rect 17598 16086 17730 16091
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17598 16053 17730 16058
rect 10934 15946 11074 15974
rect 9534 13847 9535 13873
rect 9561 13847 9562 13873
rect 9534 13481 9562 13847
rect 10374 13873 10626 13874
rect 10374 13847 10599 13873
rect 10625 13847 10626 13873
rect 10374 13846 10626 13847
rect 9534 13455 9535 13481
rect 9561 13455 9562 13481
rect 9534 13449 9562 13455
rect 9702 13481 9730 13487
rect 9702 13455 9703 13481
rect 9729 13455 9730 13481
rect 9366 13399 9367 13425
rect 9393 13399 9394 13425
rect 9254 13090 9282 13095
rect 9366 13090 9394 13399
rect 9702 13257 9730 13455
rect 9918 13342 10050 13347
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 9918 13309 10050 13314
rect 9702 13231 9703 13257
rect 9729 13231 9730 13257
rect 9702 13225 9730 13231
rect 10374 13257 10402 13846
rect 10598 13841 10626 13846
rect 10878 13874 10906 13879
rect 10878 13827 10906 13846
rect 10822 13538 10850 13543
rect 10822 13491 10850 13510
rect 10374 13231 10375 13257
rect 10401 13231 10402 13257
rect 10374 13225 10402 13231
rect 10262 13145 10290 13151
rect 10262 13119 10263 13145
rect 10289 13119 10290 13145
rect 9254 13089 9394 13090
rect 9254 13063 9255 13089
rect 9281 13063 9394 13089
rect 9254 13062 9394 13063
rect 9422 13089 9450 13095
rect 9422 13063 9423 13089
rect 9449 13063 9450 13089
rect 9142 12671 9143 12697
rect 9169 12671 9170 12697
rect 9142 12665 9170 12671
rect 9198 12698 9226 12703
rect 9142 11914 9170 11919
rect 9198 11914 9226 12670
rect 9254 12362 9282 13062
rect 9422 12698 9450 13063
rect 9534 13034 9562 13039
rect 9534 12987 9562 13006
rect 10038 13034 10066 13039
rect 10038 12809 10066 13006
rect 10038 12783 10039 12809
rect 10065 12783 10066 12809
rect 10038 12777 10066 12783
rect 9422 12665 9450 12670
rect 9982 12754 10010 12759
rect 9982 12642 10010 12726
rect 10094 12754 10122 12759
rect 10094 12753 10234 12754
rect 10094 12727 10095 12753
rect 10121 12727 10234 12753
rect 10094 12726 10234 12727
rect 10094 12721 10122 12726
rect 10206 12698 10234 12726
rect 10262 12753 10290 13119
rect 10262 12727 10263 12753
rect 10289 12727 10290 12753
rect 10262 12721 10290 12727
rect 10430 13145 10458 13151
rect 10430 13119 10431 13145
rect 10457 13119 10458 13145
rect 9814 12641 10010 12642
rect 9814 12615 9983 12641
rect 10009 12615 10010 12641
rect 9814 12614 10010 12615
rect 9254 12329 9282 12334
rect 9646 12362 9674 12367
rect 9142 11913 9226 11914
rect 9142 11887 9143 11913
rect 9169 11887 9226 11913
rect 9142 11886 9226 11887
rect 9310 11914 9338 11919
rect 9310 11913 9450 11914
rect 9310 11887 9311 11913
rect 9337 11887 9450 11913
rect 9310 11886 9450 11887
rect 9142 11881 9170 11886
rect 9310 11881 9338 11886
rect 9366 11802 9394 11807
rect 9086 11774 9226 11802
rect 9142 11634 9170 11639
rect 9142 11587 9170 11606
rect 9086 11578 9114 11583
rect 8974 11577 9114 11578
rect 8974 11551 9087 11577
rect 9113 11551 9114 11577
rect 8974 11550 9114 11551
rect 8470 10985 8498 10990
rect 8638 11046 8750 11074
rect 7910 10929 7938 10934
rect 7854 10793 7994 10794
rect 7854 10767 7855 10793
rect 7881 10767 7994 10793
rect 7854 10766 7994 10767
rect 7854 10761 7882 10766
rect 7798 10066 7882 10094
rect 7854 10065 7882 10066
rect 7854 10039 7855 10065
rect 7881 10039 7882 10065
rect 7854 10033 7882 10039
rect 7910 10065 7938 10071
rect 7910 10039 7911 10065
rect 7937 10039 7938 10065
rect 7630 10010 7658 10015
rect 7518 10009 7658 10010
rect 7518 9983 7631 10009
rect 7657 9983 7658 10009
rect 7518 9982 7658 9983
rect 7462 9963 7490 9982
rect 7630 9562 7658 9982
rect 7910 9954 7938 10039
rect 7630 9529 7658 9534
rect 7854 9926 7938 9954
rect 7854 9450 7882 9926
rect 7966 9674 7994 10766
rect 8078 10737 8106 10743
rect 8078 10711 8079 10737
rect 8105 10711 8106 10737
rect 8078 10626 8106 10711
rect 8078 10593 8106 10598
rect 8526 10514 8554 10519
rect 8526 10457 8554 10486
rect 8526 10431 8527 10457
rect 8553 10431 8554 10457
rect 8526 10425 8554 10431
rect 8582 10402 8610 10407
rect 8582 10355 8610 10374
rect 8470 10346 8498 10351
rect 8470 10299 8498 10318
rect 8638 10094 8666 11046
rect 8750 11041 8778 11046
rect 8806 11046 8890 11074
rect 8918 11186 8946 11191
rect 8806 10290 8834 11046
rect 8806 10257 8834 10262
rect 8862 10962 8890 10967
rect 8414 10066 8442 10071
rect 8414 10019 8442 10038
rect 8470 10066 8666 10094
rect 8022 10009 8050 10015
rect 8022 9983 8023 10009
rect 8049 9983 8050 10009
rect 8022 9898 8050 9983
rect 8022 9865 8050 9870
rect 8190 10009 8218 10015
rect 8190 9983 8191 10009
rect 8217 9983 8218 10009
rect 7966 9641 7994 9646
rect 8190 9674 8218 9983
rect 8190 9673 8274 9674
rect 8190 9647 8191 9673
rect 8217 9647 8274 9673
rect 8190 9646 8274 9647
rect 8190 9641 8218 9646
rect 7854 9417 7882 9422
rect 8246 9337 8274 9646
rect 8414 9506 8442 9511
rect 8414 9459 8442 9478
rect 8246 9311 8247 9337
rect 8273 9311 8274 9337
rect 8246 9305 8274 9311
rect 8414 9281 8442 9287
rect 8414 9255 8415 9281
rect 8441 9255 8442 9281
rect 8414 9170 8442 9255
rect 8414 9137 8442 9142
rect 7462 9058 7490 9063
rect 7406 9030 7462 9058
rect 7462 8889 7490 9030
rect 7462 8863 7463 8889
rect 7489 8863 7490 8889
rect 7462 8857 7490 8863
rect 7126 8689 7154 8694
rect 8302 8498 8330 8503
rect 8470 8498 8498 10066
rect 8806 9954 8834 9959
rect 8638 9730 8666 9735
rect 8526 9729 8666 9730
rect 8526 9703 8639 9729
rect 8665 9703 8666 9729
rect 8526 9702 8666 9703
rect 8526 9338 8554 9702
rect 8638 9697 8666 9702
rect 8806 9618 8834 9926
rect 8638 9590 8834 9618
rect 8582 9562 8610 9567
rect 8582 9515 8610 9534
rect 8638 9506 8666 9590
rect 8862 9562 8890 10934
rect 8918 10906 8946 11158
rect 8918 10859 8946 10878
rect 8974 10514 9002 11550
rect 9086 11545 9114 11550
rect 9142 11466 9170 11471
rect 9198 11466 9226 11774
rect 9142 11465 9226 11466
rect 9142 11439 9143 11465
rect 9169 11439 9226 11465
rect 9142 11438 9226 11439
rect 9142 11433 9170 11438
rect 9254 11410 9282 11415
rect 9366 11410 9394 11774
rect 9282 11382 9394 11410
rect 9254 11377 9282 11382
rect 9030 11186 9058 11191
rect 9030 11185 9226 11186
rect 9030 11159 9031 11185
rect 9057 11159 9226 11185
rect 9030 11158 9226 11159
rect 9030 11153 9058 11158
rect 9142 11018 9170 11023
rect 9142 10850 9170 10990
rect 9198 10906 9226 11158
rect 9310 10906 9338 10911
rect 9198 10878 9310 10906
rect 9310 10859 9338 10878
rect 9142 10822 9282 10850
rect 8974 10481 9002 10486
rect 9086 10793 9114 10799
rect 9086 10767 9087 10793
rect 9113 10767 9114 10793
rect 8918 10401 8946 10407
rect 8918 10375 8919 10401
rect 8945 10375 8946 10401
rect 8918 9730 8946 10375
rect 8974 10290 9002 10295
rect 8974 10094 9002 10262
rect 8974 10066 9058 10094
rect 8918 9697 8946 9702
rect 8806 9534 9002 9562
rect 8526 9310 8610 9338
rect 8526 9226 8554 9231
rect 8526 8889 8554 9198
rect 8526 8863 8527 8889
rect 8553 8863 8554 8889
rect 8526 8857 8554 8863
rect 8526 8498 8554 8503
rect 8470 8470 8526 8498
rect 7294 8442 7322 8447
rect 7070 8441 7322 8442
rect 7070 8415 7071 8441
rect 7097 8415 7295 8441
rect 7321 8415 7322 8441
rect 7070 8414 7322 8415
rect 7070 8409 7098 8414
rect 7294 8409 7322 8414
rect 5614 8359 5615 8385
rect 5641 8359 5642 8385
rect 5614 8353 5642 8359
rect 2238 8246 2370 8251
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2238 8213 2370 8218
rect 8302 7713 8330 8470
rect 8526 8465 8554 8470
rect 8582 8274 8610 9310
rect 8638 8946 8666 9478
rect 8694 9505 8722 9511
rect 8694 9479 8695 9505
rect 8721 9479 8722 9505
rect 8694 9450 8722 9479
rect 8806 9505 8834 9534
rect 8806 9479 8807 9505
rect 8833 9479 8834 9505
rect 8806 9473 8834 9479
rect 8694 9417 8722 9422
rect 8918 9450 8946 9455
rect 8918 9337 8946 9422
rect 8918 9311 8919 9337
rect 8945 9311 8946 9337
rect 8918 9305 8946 9311
rect 8750 9281 8778 9287
rect 8750 9255 8751 9281
rect 8777 9255 8778 9281
rect 8750 9058 8778 9255
rect 8750 9025 8778 9030
rect 8638 8918 8778 8946
rect 8582 8241 8610 8246
rect 8750 8889 8778 8918
rect 8750 8863 8751 8889
rect 8777 8863 8778 8889
rect 8302 7687 8303 7713
rect 8329 7687 8330 7713
rect 8302 7681 8330 7687
rect 8358 7714 8386 7719
rect 8358 7667 8386 7686
rect 8470 7658 8498 7663
rect 8470 7611 8498 7630
rect 7910 7602 7938 7607
rect 2238 7462 2370 7467
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2238 7429 2370 7434
rect 7910 7321 7938 7574
rect 7910 7295 7911 7321
rect 7937 7295 7938 7321
rect 7910 7289 7938 7295
rect 7574 7266 7602 7271
rect 7518 7238 7574 7266
rect 2238 6678 2370 6683
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2238 6645 2370 6650
rect 7518 6481 7546 7238
rect 7574 7219 7602 7238
rect 8750 7266 8778 8863
rect 8974 8890 9002 9534
rect 9030 9505 9058 10066
rect 9086 9786 9114 10767
rect 9254 10794 9282 10822
rect 9254 10793 9338 10794
rect 9254 10767 9255 10793
rect 9281 10767 9338 10793
rect 9254 10766 9338 10767
rect 9254 10761 9282 10766
rect 9254 10682 9282 10687
rect 9198 10345 9226 10351
rect 9198 10319 9199 10345
rect 9225 10319 9226 10345
rect 9198 10066 9226 10319
rect 9198 10033 9226 10038
rect 9086 9753 9114 9758
rect 9030 9479 9031 9505
rect 9057 9479 9058 9505
rect 9030 8946 9058 9479
rect 9142 9730 9170 9735
rect 9086 9226 9114 9231
rect 9086 9179 9114 9198
rect 9142 9225 9170 9702
rect 9198 9561 9226 9567
rect 9198 9535 9199 9561
rect 9225 9535 9226 9561
rect 9198 9450 9226 9535
rect 9198 9417 9226 9422
rect 9142 9199 9143 9225
rect 9169 9199 9170 9225
rect 9142 9193 9170 9199
rect 9086 8946 9114 8951
rect 9030 8918 9086 8946
rect 9086 8913 9114 8918
rect 8974 8862 9058 8890
rect 9030 8834 9058 8862
rect 9142 8834 9170 8839
rect 9030 8833 9170 8834
rect 9030 8807 9143 8833
rect 9169 8807 9170 8833
rect 9030 8806 9170 8807
rect 8862 8778 8890 8783
rect 8806 8162 8834 8167
rect 8862 8162 8890 8750
rect 9086 8497 9114 8806
rect 9142 8801 9170 8806
rect 9254 8778 9282 10654
rect 9310 9225 9338 10766
rect 9366 9954 9394 11382
rect 9422 10738 9450 11886
rect 9646 11802 9674 12334
rect 9646 11769 9674 11774
rect 9758 11858 9786 11863
rect 9758 11689 9786 11830
rect 9758 11663 9759 11689
rect 9785 11663 9786 11689
rect 9758 11657 9786 11663
rect 9646 11577 9674 11583
rect 9646 11551 9647 11577
rect 9673 11551 9674 11577
rect 9478 11186 9506 11191
rect 9478 11139 9506 11158
rect 9590 11129 9618 11135
rect 9590 11103 9591 11129
rect 9617 11103 9618 11129
rect 9590 10962 9618 11103
rect 9646 11018 9674 11551
rect 9646 10985 9674 10990
rect 9702 11298 9730 11303
rect 9590 10929 9618 10934
rect 9646 10906 9674 10911
rect 9590 10850 9618 10855
rect 9590 10738 9618 10822
rect 9422 10737 9618 10738
rect 9422 10711 9591 10737
rect 9617 10711 9618 10737
rect 9422 10710 9618 10711
rect 9534 10346 9562 10710
rect 9590 10705 9618 10710
rect 9590 10402 9618 10407
rect 9590 10355 9618 10374
rect 9534 10299 9562 10318
rect 9366 9921 9394 9926
rect 9422 10066 9450 10071
rect 9422 9561 9450 10038
rect 9422 9535 9423 9561
rect 9449 9535 9450 9561
rect 9422 9529 9450 9535
rect 9478 9786 9506 9791
rect 9310 9199 9311 9225
rect 9337 9199 9338 9225
rect 9310 9170 9338 9199
rect 9478 9338 9506 9758
rect 9534 9674 9562 9679
rect 9534 9617 9562 9646
rect 9534 9591 9535 9617
rect 9561 9591 9562 9617
rect 9534 9585 9562 9591
rect 9310 9137 9338 9142
rect 9366 9169 9394 9175
rect 9366 9143 9367 9169
rect 9393 9143 9394 9169
rect 9366 9114 9394 9143
rect 9310 8778 9338 8783
rect 9282 8777 9338 8778
rect 9282 8751 9311 8777
rect 9337 8751 9338 8777
rect 9282 8750 9338 8751
rect 9254 8731 9282 8750
rect 9310 8745 9338 8750
rect 9366 8610 9394 9086
rect 9478 8889 9506 9310
rect 9478 8863 9479 8889
rect 9505 8863 9506 8889
rect 9478 8857 9506 8863
rect 9534 9281 9562 9287
rect 9534 9255 9535 9281
rect 9561 9255 9562 9281
rect 9534 9226 9562 9255
rect 9534 8834 9562 9198
rect 9646 9226 9674 10878
rect 9702 10738 9730 11270
rect 9758 11129 9786 11135
rect 9758 11103 9759 11129
rect 9785 11103 9786 11129
rect 9758 10850 9786 11103
rect 9814 11073 9842 12614
rect 9982 12609 10010 12614
rect 10150 12642 10178 12647
rect 9918 12558 10050 12563
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 9918 12525 10050 12530
rect 10150 12474 10178 12614
rect 10038 12446 10178 12474
rect 10038 12417 10066 12446
rect 10038 12391 10039 12417
rect 10065 12391 10066 12417
rect 10038 12385 10066 12391
rect 10206 11858 10234 12670
rect 10206 11825 10234 11830
rect 9918 11774 10050 11779
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 9918 11741 10050 11746
rect 10430 11746 10458 13119
rect 10766 13146 10794 13151
rect 10654 13034 10682 13039
rect 10654 12754 10682 13006
rect 10654 12707 10682 12726
rect 10766 12753 10794 13118
rect 10990 13034 11018 13039
rect 10990 12987 11018 13006
rect 10990 12810 11018 12815
rect 10934 12754 10962 12759
rect 10766 12727 10767 12753
rect 10793 12727 10794 12753
rect 10766 12721 10794 12727
rect 10822 12753 10962 12754
rect 10822 12727 10935 12753
rect 10961 12727 10962 12753
rect 10822 12726 10962 12727
rect 10598 12642 10626 12647
rect 10598 12595 10626 12614
rect 10822 12025 10850 12726
rect 10934 12721 10962 12726
rect 10878 12642 10906 12647
rect 10990 12642 11018 12782
rect 10878 12641 11018 12642
rect 10878 12615 10879 12641
rect 10905 12615 11018 12641
rect 10878 12614 11018 12615
rect 10878 12609 10906 12614
rect 10822 11999 10823 12025
rect 10849 11999 10850 12025
rect 10822 11993 10850 11999
rect 11046 12306 11074 15946
rect 12222 15946 12306 15974
rect 12222 13593 12250 15946
rect 17598 15302 17730 15307
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17598 15269 17730 15274
rect 17598 14518 17730 14523
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17598 14485 17730 14490
rect 12222 13567 12223 13593
rect 12249 13567 12250 13593
rect 11158 13482 11186 13487
rect 11158 13481 11242 13482
rect 11158 13455 11159 13481
rect 11185 13455 11242 13481
rect 11158 13454 11242 13455
rect 11158 13449 11186 13454
rect 11102 13201 11130 13207
rect 11102 13175 11103 13201
rect 11129 13175 11130 13201
rect 11102 12698 11130 13175
rect 11158 13034 11186 13039
rect 11158 12987 11186 13006
rect 11214 12809 11242 13454
rect 11718 13426 11746 13431
rect 11718 13201 11746 13398
rect 12222 13426 12250 13567
rect 12390 13873 12418 13879
rect 12390 13847 12391 13873
rect 12417 13847 12418 13873
rect 12390 13538 12418 13847
rect 17598 13734 17730 13739
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17598 13701 17730 13706
rect 13846 13593 13874 13599
rect 13846 13567 13847 13593
rect 13873 13567 13874 13593
rect 12390 13491 12418 13510
rect 12670 13538 12698 13543
rect 12222 13393 12250 13398
rect 12278 13482 12306 13487
rect 12278 13257 12306 13454
rect 12278 13231 12279 13257
rect 12305 13231 12306 13257
rect 12278 13225 12306 13231
rect 12670 13426 12698 13510
rect 12782 13482 12810 13487
rect 12782 13435 12810 13454
rect 11718 13175 11719 13201
rect 11745 13175 11746 13201
rect 11718 13169 11746 13175
rect 12166 13201 12194 13207
rect 12166 13175 12167 13201
rect 12193 13175 12194 13201
rect 11942 13145 11970 13151
rect 11942 13119 11943 13145
rect 11969 13119 11970 13145
rect 11662 13033 11690 13039
rect 11662 13007 11663 13033
rect 11689 13007 11690 13033
rect 11662 12865 11690 13007
rect 11662 12839 11663 12865
rect 11689 12839 11690 12865
rect 11662 12833 11690 12839
rect 11214 12783 11215 12809
rect 11241 12783 11242 12809
rect 11214 12777 11242 12783
rect 11438 12810 11466 12815
rect 11102 12665 11130 12670
rect 11158 12753 11186 12759
rect 11158 12727 11159 12753
rect 11185 12727 11186 12753
rect 11102 12306 11130 12311
rect 11046 12305 11130 12306
rect 11046 12279 11103 12305
rect 11129 12279 11130 12305
rect 11046 12278 11130 12279
rect 11046 11969 11074 12278
rect 11102 12273 11130 12278
rect 11046 11943 11047 11969
rect 11073 11943 11074 11969
rect 11046 11937 11074 11943
rect 10822 11913 10850 11919
rect 10822 11887 10823 11913
rect 10849 11887 10850 11913
rect 10654 11858 10682 11863
rect 10654 11811 10682 11830
rect 10766 11857 10794 11863
rect 10766 11831 10767 11857
rect 10793 11831 10794 11857
rect 10430 11713 10458 11718
rect 10710 11746 10738 11751
rect 10710 11129 10738 11718
rect 10710 11103 10711 11129
rect 10737 11103 10738 11129
rect 10710 11097 10738 11103
rect 9814 11047 9815 11073
rect 9841 11047 9842 11073
rect 9814 11041 9842 11047
rect 10542 11074 10570 11079
rect 9918 10990 10050 10995
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 9918 10957 10050 10962
rect 10542 10962 10570 11046
rect 10766 10962 10794 11831
rect 10822 11746 10850 11887
rect 10822 11713 10850 11718
rect 11158 11914 11186 12727
rect 11326 12698 11354 12703
rect 11326 12651 11354 12670
rect 11438 12697 11466 12782
rect 11942 12810 11970 13119
rect 11942 12777 11970 12782
rect 11606 12754 11634 12759
rect 12166 12754 12194 13175
rect 12222 13202 12250 13207
rect 12222 13155 12250 13174
rect 12334 13146 12362 13151
rect 12670 13146 12698 13398
rect 13846 13370 13874 13567
rect 20006 13593 20034 13599
rect 20006 13567 20007 13593
rect 20033 13567 20034 13593
rect 18942 13537 18970 13543
rect 18942 13511 18943 13537
rect 18969 13511 18970 13537
rect 14070 13481 14098 13487
rect 14070 13455 14071 13481
rect 14097 13455 14098 13481
rect 14070 13426 14098 13455
rect 14098 13398 14322 13426
rect 14070 13393 14098 13398
rect 13734 13342 13846 13370
rect 12334 13145 12474 13146
rect 12334 13119 12335 13145
rect 12361 13119 12474 13145
rect 12334 13118 12474 13119
rect 12334 13113 12362 13118
rect 12334 13034 12362 13039
rect 12334 12865 12362 13006
rect 12334 12839 12335 12865
rect 12361 12839 12362 12865
rect 12334 12833 12362 12839
rect 12390 12754 12418 12759
rect 11606 12753 11690 12754
rect 11606 12727 11607 12753
rect 11633 12727 11690 12753
rect 11606 12726 11690 12727
rect 12166 12753 12418 12754
rect 12166 12727 12391 12753
rect 12417 12727 12418 12753
rect 12166 12726 12418 12727
rect 11606 12721 11634 12726
rect 11438 12671 11439 12697
rect 11465 12671 11466 12697
rect 11438 12665 11466 12671
rect 11662 12698 11690 12726
rect 11326 12362 11354 12367
rect 11326 12315 11354 12334
rect 10878 11074 10906 11079
rect 10878 11027 10906 11046
rect 11046 11074 11074 11079
rect 11158 11074 11186 11886
rect 11438 11186 11466 11191
rect 11438 11185 11522 11186
rect 11438 11159 11439 11185
rect 11465 11159 11522 11185
rect 11438 11158 11522 11159
rect 11438 11153 11466 11158
rect 11046 11073 11186 11074
rect 11046 11047 11047 11073
rect 11073 11047 11186 11073
rect 11046 11046 11186 11047
rect 11214 11074 11242 11079
rect 10542 10934 10794 10962
rect 10542 10905 10570 10934
rect 10542 10879 10543 10905
rect 10569 10879 10570 10905
rect 10542 10873 10570 10879
rect 9758 10817 9786 10822
rect 9814 10793 9842 10799
rect 9814 10767 9815 10793
rect 9841 10767 9842 10793
rect 9702 10710 9786 10738
rect 9758 10457 9786 10710
rect 9758 10431 9759 10457
rect 9785 10431 9786 10457
rect 9758 10425 9786 10431
rect 9646 9193 9674 9198
rect 9702 10402 9730 10407
rect 9702 8946 9730 10374
rect 9758 9505 9786 9511
rect 9758 9479 9759 9505
rect 9785 9479 9786 9505
rect 9758 9450 9786 9479
rect 9758 9417 9786 9422
rect 9814 9282 9842 10767
rect 10710 10794 10738 10799
rect 10710 10747 10738 10766
rect 10374 10738 10402 10743
rect 10374 10402 10402 10710
rect 10654 10402 10682 10407
rect 10374 10401 10682 10402
rect 10374 10375 10655 10401
rect 10681 10375 10682 10401
rect 10374 10374 10682 10375
rect 10654 10369 10682 10374
rect 10430 10290 10458 10295
rect 9918 10206 10050 10211
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 9918 10173 10050 10178
rect 10206 9898 10234 9903
rect 10234 9870 10290 9898
rect 10206 9865 10234 9870
rect 9870 9730 9898 9735
rect 9870 9617 9898 9702
rect 9870 9591 9871 9617
rect 9897 9591 9898 9617
rect 9870 9585 9898 9591
rect 10094 9506 10122 9511
rect 9918 9422 10050 9427
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 9918 9389 10050 9394
rect 10094 9338 10122 9478
rect 9926 9310 10122 9338
rect 10150 9505 10178 9511
rect 10150 9479 10151 9505
rect 10177 9479 10178 9505
rect 9870 9282 9898 9287
rect 9814 9254 9870 9282
rect 9870 9225 9898 9254
rect 9870 9199 9871 9225
rect 9897 9199 9898 9225
rect 9870 9193 9898 9199
rect 9702 8918 9786 8946
rect 9702 8834 9730 8839
rect 9534 8833 9730 8834
rect 9534 8807 9703 8833
rect 9729 8807 9730 8833
rect 9534 8806 9730 8807
rect 9702 8801 9730 8806
rect 9198 8582 9394 8610
rect 9478 8722 9506 8727
rect 9086 8471 9087 8497
rect 9113 8471 9114 8497
rect 9086 8386 9114 8471
rect 9142 8498 9170 8503
rect 9142 8451 9170 8470
rect 9086 8353 9114 8358
rect 9198 8274 9226 8582
rect 9254 8498 9282 8503
rect 9422 8498 9450 8503
rect 9254 8497 9450 8498
rect 9254 8471 9255 8497
rect 9281 8471 9423 8497
rect 9449 8471 9450 8497
rect 9254 8470 9450 8471
rect 9254 8465 9282 8470
rect 9422 8465 9450 8470
rect 9478 8497 9506 8694
rect 9478 8471 9479 8497
rect 9505 8471 9506 8497
rect 9478 8465 9506 8471
rect 9758 8498 9786 8918
rect 9926 8777 9954 9310
rect 9982 9226 10010 9231
rect 10010 9198 10066 9226
rect 9982 9193 10010 9198
rect 10038 8833 10066 9198
rect 10150 9170 10178 9479
rect 10150 9137 10178 9142
rect 10206 9505 10234 9511
rect 10206 9479 10207 9505
rect 10233 9479 10234 9505
rect 10206 9058 10234 9479
rect 10038 8807 10039 8833
rect 10065 8807 10066 8833
rect 10038 8801 10066 8807
rect 10094 9030 10206 9058
rect 9926 8751 9927 8777
rect 9953 8751 9954 8777
rect 9926 8745 9954 8751
rect 9918 8638 10050 8643
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 9918 8605 10050 8610
rect 9758 8465 9786 8470
rect 9814 8497 9842 8503
rect 9814 8471 9815 8497
rect 9841 8471 9842 8497
rect 9814 8386 9842 8471
rect 9926 8498 9954 8503
rect 9926 8441 9954 8470
rect 10094 8442 10122 9030
rect 10206 9025 10234 9030
rect 10262 8834 10290 9870
rect 10430 9617 10458 10262
rect 11046 10290 11074 11046
rect 11158 10794 11186 10799
rect 11214 10794 11242 11046
rect 11494 10906 11522 11158
rect 11550 11130 11578 11135
rect 11550 11129 11634 11130
rect 11550 11103 11551 11129
rect 11577 11103 11634 11129
rect 11550 11102 11634 11103
rect 11550 11097 11578 11102
rect 11606 10906 11634 11102
rect 11494 10878 11578 10906
rect 11494 10794 11522 10799
rect 11214 10793 11522 10794
rect 11214 10767 11495 10793
rect 11521 10767 11522 10793
rect 11214 10766 11522 10767
rect 11046 10257 11074 10262
rect 11102 10737 11130 10743
rect 11102 10711 11103 10737
rect 11129 10711 11130 10737
rect 10430 9591 10431 9617
rect 10457 9591 10458 9617
rect 10374 9562 10402 9567
rect 10374 9282 10402 9534
rect 10430 9282 10458 9591
rect 10598 9954 10626 9959
rect 10430 9254 10570 9282
rect 9926 8415 9927 8441
rect 9953 8415 9954 8441
rect 9926 8409 9954 8415
rect 10038 8414 10122 8442
rect 10150 8806 10290 8834
rect 10318 9225 10346 9231
rect 10318 9199 10319 9225
rect 10345 9199 10346 9225
rect 10318 9114 10346 9199
rect 10318 8834 10346 9086
rect 10374 9058 10402 9254
rect 10374 9025 10402 9030
rect 10430 9169 10458 9175
rect 10430 9143 10431 9169
rect 10457 9143 10458 9169
rect 10430 8890 10458 9143
rect 10430 8857 10458 8862
rect 10486 9113 10514 9119
rect 10486 9087 10487 9113
rect 10513 9087 10514 9113
rect 10374 8834 10402 8839
rect 10318 8806 10374 8834
rect 9814 8353 9842 8358
rect 9422 8330 9450 8335
rect 10038 8330 10066 8414
rect 9422 8329 9506 8330
rect 9422 8303 9423 8329
rect 9449 8303 9506 8329
rect 9422 8302 9506 8303
rect 9422 8297 9450 8302
rect 8806 8161 8862 8162
rect 8806 8135 8807 8161
rect 8833 8135 8862 8161
rect 8806 8134 8862 8135
rect 8806 8129 8834 8134
rect 8862 8115 8890 8134
rect 9030 8246 9226 8274
rect 9366 8274 9394 8279
rect 8974 8049 9002 8055
rect 8974 8023 8975 8049
rect 9001 8023 9002 8049
rect 8862 7937 8890 7943
rect 8862 7911 8863 7937
rect 8889 7911 8890 7937
rect 8806 7714 8834 7719
rect 8806 7574 8834 7686
rect 8862 7657 8890 7911
rect 8862 7631 8863 7657
rect 8889 7631 8890 7657
rect 8862 7625 8890 7631
rect 8918 7714 8946 7719
rect 8918 7657 8946 7686
rect 8918 7631 8919 7657
rect 8945 7631 8946 7657
rect 8918 7625 8946 7631
rect 8806 7546 8946 7574
rect 8750 7233 8778 7238
rect 7854 6986 7882 6991
rect 7854 6537 7882 6958
rect 7854 6511 7855 6537
rect 7881 6511 7882 6537
rect 7854 6505 7882 6511
rect 8918 6537 8946 7546
rect 8918 6511 8919 6537
rect 8945 6511 8946 6537
rect 7518 6455 7519 6481
rect 7545 6455 7546 6481
rect 7518 6449 7546 6455
rect 2238 5894 2370 5899
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2238 5861 2370 5866
rect 2238 5110 2370 5115
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2238 5077 2370 5082
rect 2238 4326 2370 4331
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2238 4293 2370 4298
rect 2238 3542 2370 3547
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2238 3509 2370 3514
rect 2238 2758 2370 2763
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2238 2725 2370 2730
rect 8918 2169 8946 6511
rect 8918 2143 8919 2169
rect 8945 2143 8946 2169
rect 8918 2137 8946 2143
rect 8974 7321 9002 8023
rect 9030 7657 9058 8246
rect 9030 7631 9031 7657
rect 9057 7631 9058 7657
rect 9030 7625 9058 7631
rect 9198 7658 9226 7663
rect 9198 7611 9226 7630
rect 9366 7658 9394 8246
rect 9366 7611 9394 7630
rect 9478 7714 9506 8302
rect 9926 8302 10066 8330
rect 9758 8162 9786 8167
rect 9758 8049 9786 8134
rect 9870 8106 9898 8111
rect 9926 8106 9954 8302
rect 9870 8105 9954 8106
rect 9870 8079 9871 8105
rect 9897 8079 9954 8105
rect 9870 8078 9954 8079
rect 9870 8073 9898 8078
rect 9758 8023 9759 8049
rect 9785 8023 9786 8049
rect 9758 8017 9786 8023
rect 9982 8050 10010 8055
rect 9982 8003 10010 8022
rect 10094 8050 10122 8055
rect 10150 8050 10178 8806
rect 10374 8801 10402 8806
rect 10486 8554 10514 9087
rect 10486 8521 10514 8526
rect 10542 8330 10570 9254
rect 10598 9225 10626 9926
rect 11102 9954 11130 10711
rect 11102 9921 11130 9926
rect 10990 9674 11018 9679
rect 10990 9627 11018 9646
rect 10822 9618 10850 9623
rect 10654 9562 10682 9567
rect 10654 9515 10682 9534
rect 10822 9562 10850 9590
rect 11158 9618 11186 10766
rect 11494 10094 11522 10766
rect 11382 10066 11522 10094
rect 11326 10010 11354 10015
rect 11326 9963 11354 9982
rect 11158 9571 11186 9590
rect 11382 9617 11410 10066
rect 11550 9674 11578 10878
rect 11606 10873 11634 10878
rect 11662 11074 11690 12670
rect 12334 11298 12362 11303
rect 12334 11185 12362 11270
rect 12334 11159 12335 11185
rect 12361 11159 12362 11185
rect 12334 11153 12362 11159
rect 11606 10738 11634 10743
rect 11662 10738 11690 11046
rect 11606 10737 11690 10738
rect 11606 10711 11607 10737
rect 11633 10711 11690 10737
rect 11606 10710 11690 10711
rect 11718 11129 11746 11135
rect 11718 11103 11719 11129
rect 11745 11103 11746 11129
rect 11606 10705 11634 10710
rect 11718 10094 11746 11103
rect 11998 11130 12026 11135
rect 11998 11083 12026 11102
rect 12390 11129 12418 12726
rect 12446 12698 12474 13118
rect 12614 13145 12698 13146
rect 12614 13119 12671 13145
rect 12697 13119 12698 13145
rect 12614 13118 12698 13119
rect 12446 12665 12474 12670
rect 12502 12810 12530 12815
rect 12502 12697 12530 12782
rect 12502 12671 12503 12697
rect 12529 12671 12530 12697
rect 12502 12665 12530 12671
rect 12614 11577 12642 13118
rect 12670 13113 12698 13118
rect 13678 13202 13706 13207
rect 13006 13090 13034 13095
rect 12838 13089 13034 13090
rect 12838 13063 13007 13089
rect 13033 13063 13034 13089
rect 12838 13062 13034 13063
rect 12838 12809 12866 13062
rect 13006 13057 13034 13062
rect 13510 13090 13538 13095
rect 12838 12783 12839 12809
rect 12865 12783 12866 12809
rect 12838 12777 12866 12783
rect 13510 12809 13538 13062
rect 13678 12865 13706 13174
rect 13678 12839 13679 12865
rect 13705 12839 13706 12865
rect 13678 12833 13706 12839
rect 13510 12783 13511 12809
rect 13537 12783 13538 12809
rect 13510 12777 13538 12783
rect 13734 12809 13762 13342
rect 13846 13337 13874 13342
rect 14294 13257 14322 13398
rect 14294 13231 14295 13257
rect 14321 13231 14322 13257
rect 14070 13090 14098 13095
rect 14070 13043 14098 13062
rect 13734 12783 13735 12809
rect 13761 12783 13762 12809
rect 13734 12777 13762 12783
rect 12782 12754 12810 12759
rect 12782 12707 12810 12726
rect 13454 12754 13482 12759
rect 13454 12707 13482 12726
rect 12670 12698 12698 12703
rect 12670 12651 12698 12670
rect 12726 11970 12754 11975
rect 12670 11914 12698 11919
rect 12670 11867 12698 11886
rect 12726 11913 12754 11942
rect 13062 11969 13090 11975
rect 13062 11943 13063 11969
rect 13089 11943 13090 11969
rect 12726 11887 12727 11913
rect 12753 11887 12754 11913
rect 12726 11881 12754 11887
rect 12838 11914 12866 11919
rect 12950 11914 12978 11919
rect 12838 11913 12978 11914
rect 12838 11887 12839 11913
rect 12865 11887 12951 11913
rect 12977 11887 12978 11913
rect 12838 11886 12978 11887
rect 12838 11881 12866 11886
rect 12950 11881 12978 11886
rect 13006 11857 13034 11863
rect 13006 11831 13007 11857
rect 13033 11831 13034 11857
rect 13006 11633 13034 11831
rect 13006 11607 13007 11633
rect 13033 11607 13034 11633
rect 13006 11601 13034 11607
rect 12614 11551 12615 11577
rect 12641 11551 12642 11577
rect 12614 11545 12642 11551
rect 13062 11298 13090 11943
rect 14070 11970 14098 11975
rect 13062 11265 13090 11270
rect 13230 11913 13258 11919
rect 13230 11887 13231 11913
rect 13257 11887 13258 11913
rect 12390 11103 12391 11129
rect 12417 11103 12418 11129
rect 12390 11097 12418 11103
rect 12614 11185 12642 11191
rect 12614 11159 12615 11185
rect 12641 11159 12642 11185
rect 12614 11074 12642 11159
rect 13062 11185 13090 11191
rect 13062 11159 13063 11185
rect 13089 11159 13090 11185
rect 12614 11041 12642 11046
rect 13006 11129 13034 11135
rect 13006 11103 13007 11129
rect 13033 11103 13034 11129
rect 11886 10906 11914 10911
rect 11550 9641 11578 9646
rect 11606 10066 11746 10094
rect 11830 10682 11858 10687
rect 11382 9591 11383 9617
rect 11409 9591 11410 9617
rect 10822 9561 10906 9562
rect 10822 9535 10823 9561
rect 10849 9535 10906 9561
rect 10822 9534 10906 9535
rect 10822 9529 10850 9534
rect 10878 9337 10906 9534
rect 10878 9311 10879 9337
rect 10905 9311 10906 9337
rect 10878 9305 10906 9311
rect 11214 9450 11242 9455
rect 10598 9199 10599 9225
rect 10625 9199 10626 9225
rect 10598 9193 10626 9199
rect 10766 9226 10794 9231
rect 10766 9179 10794 9198
rect 10710 9170 10738 9175
rect 10710 8946 10738 9142
rect 11046 9170 11074 9175
rect 11046 9123 11074 9142
rect 10934 9114 10962 9119
rect 10934 9113 11018 9114
rect 10934 9087 10935 9113
rect 10961 9087 11018 9113
rect 10934 9086 11018 9087
rect 10934 9081 10962 9086
rect 10654 8918 10738 8946
rect 10654 8498 10682 8918
rect 10654 8451 10682 8470
rect 10710 8833 10738 8839
rect 10710 8807 10711 8833
rect 10737 8807 10738 8833
rect 10710 8442 10738 8807
rect 10710 8409 10738 8414
rect 10766 8834 10794 8839
rect 10766 8441 10794 8806
rect 10990 8778 11018 9086
rect 11046 8890 11074 8895
rect 11046 8843 11074 8862
rect 11158 8778 11186 8783
rect 10990 8750 11158 8778
rect 11046 8554 11074 8559
rect 11046 8507 11074 8526
rect 11158 8553 11186 8750
rect 11158 8527 11159 8553
rect 11185 8527 11186 8553
rect 11158 8521 11186 8527
rect 11214 8722 11242 9422
rect 11326 9226 11354 9231
rect 11326 9179 11354 9198
rect 11214 8497 11242 8694
rect 11382 8554 11410 9591
rect 11606 9617 11634 10066
rect 11606 9591 11607 9617
rect 11633 9591 11634 9617
rect 11606 9338 11634 9591
rect 11606 9305 11634 9310
rect 11830 9338 11858 10654
rect 11886 9561 11914 10878
rect 11998 10737 12026 10743
rect 11998 10711 11999 10737
rect 12025 10711 12026 10737
rect 11886 9535 11887 9561
rect 11913 9535 11914 9561
rect 11886 9529 11914 9535
rect 11942 10066 11970 10071
rect 11830 9305 11858 9310
rect 11606 8554 11634 8559
rect 11382 8553 11634 8554
rect 11382 8527 11607 8553
rect 11633 8527 11634 8553
rect 11382 8526 11634 8527
rect 11606 8521 11634 8526
rect 11774 8554 11802 8559
rect 11774 8507 11802 8526
rect 11214 8471 11215 8497
rect 11241 8471 11242 8497
rect 11214 8465 11242 8471
rect 11942 8497 11970 10038
rect 11998 9562 12026 10711
rect 11998 9226 12026 9534
rect 12110 10737 12138 10743
rect 12110 10711 12111 10737
rect 12137 10711 12138 10737
rect 12110 9450 12138 10711
rect 12334 10737 12362 10743
rect 12334 10711 12335 10737
rect 12361 10711 12362 10737
rect 12278 10681 12306 10687
rect 12278 10655 12279 10681
rect 12305 10655 12306 10681
rect 12278 10094 12306 10655
rect 12166 10066 12194 10071
rect 12166 10019 12194 10038
rect 12222 10066 12306 10094
rect 12334 10094 12362 10711
rect 12558 10345 12586 10351
rect 12558 10319 12559 10345
rect 12585 10319 12586 10345
rect 12558 10094 12586 10319
rect 12334 10066 12474 10094
rect 12558 10066 12642 10094
rect 12110 9422 12194 9450
rect 12054 9338 12082 9343
rect 12054 9291 12082 9310
rect 12110 9226 12138 9231
rect 11998 9225 12082 9226
rect 11998 9199 11999 9225
rect 12025 9199 12082 9225
rect 11998 9198 12082 9199
rect 11998 9193 12026 9198
rect 11942 8471 11943 8497
rect 11969 8471 11970 8497
rect 10766 8415 10767 8441
rect 10793 8415 10794 8441
rect 10766 8409 10794 8415
rect 10934 8330 10962 8335
rect 10542 8302 10794 8330
rect 10094 8049 10178 8050
rect 10094 8023 10095 8049
rect 10121 8023 10178 8049
rect 10094 8022 10178 8023
rect 10262 8049 10290 8055
rect 10262 8023 10263 8049
rect 10289 8023 10290 8049
rect 10094 8017 10122 8022
rect 10038 7938 10066 7943
rect 10038 7937 10178 7938
rect 10038 7911 10039 7937
rect 10065 7911 10178 7937
rect 10038 7910 10178 7911
rect 10038 7905 10066 7910
rect 9918 7854 10050 7859
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 9918 7821 10050 7826
rect 10150 7770 10178 7910
rect 10262 7882 10290 8023
rect 10262 7849 10290 7854
rect 10150 7742 10290 7770
rect 9478 7657 9506 7686
rect 9478 7631 9479 7657
rect 9505 7631 9506 7657
rect 9478 7625 9506 7631
rect 10038 7714 10066 7719
rect 9086 7602 9114 7607
rect 9086 7555 9114 7574
rect 9310 7601 9338 7607
rect 9310 7575 9311 7601
rect 9337 7575 9338 7601
rect 8974 7295 8975 7321
rect 9001 7295 9002 7321
rect 8750 2058 8778 2063
rect 2238 1974 2370 1979
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2238 1941 2370 1946
rect 8750 400 8778 2030
rect 8974 1777 9002 7295
rect 9198 7266 9226 7271
rect 9142 6538 9170 6543
rect 9198 6538 9226 7238
rect 9310 6986 9338 7575
rect 9310 6953 9338 6958
rect 9590 7266 9618 7271
rect 9590 6986 9618 7238
rect 10038 7265 10066 7686
rect 10038 7239 10039 7265
rect 10065 7239 10066 7265
rect 10038 7233 10066 7239
rect 10150 7658 10178 7663
rect 10150 7265 10178 7630
rect 10150 7239 10151 7265
rect 10177 7239 10178 7265
rect 10150 7233 10178 7239
rect 10206 7154 10234 7159
rect 10094 7153 10234 7154
rect 10094 7127 10207 7153
rect 10233 7127 10234 7153
rect 10094 7126 10234 7127
rect 9918 7070 10050 7075
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 9918 7037 10050 7042
rect 9590 6985 9786 6986
rect 9590 6959 9591 6985
rect 9617 6959 9786 6985
rect 9590 6958 9786 6959
rect 9142 6537 9226 6538
rect 9142 6511 9143 6537
rect 9169 6511 9226 6537
rect 9142 6510 9226 6511
rect 9142 6505 9170 6510
rect 9534 6202 9562 6207
rect 9590 6202 9618 6958
rect 9758 6873 9786 6958
rect 9758 6847 9759 6873
rect 9785 6847 9786 6873
rect 9758 6841 9786 6847
rect 9918 6286 10050 6291
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 9918 6253 10050 6258
rect 9534 6201 9730 6202
rect 9534 6175 9535 6201
rect 9561 6175 9730 6201
rect 9534 6174 9730 6175
rect 9534 6169 9562 6174
rect 9702 6089 9730 6174
rect 10094 6145 10122 7126
rect 10206 7121 10234 7126
rect 10150 6930 10178 6935
rect 10262 6930 10290 7742
rect 10374 7266 10402 7271
rect 10710 7266 10738 7271
rect 10374 7265 10738 7266
rect 10374 7239 10375 7265
rect 10401 7239 10711 7265
rect 10737 7239 10738 7265
rect 10374 7238 10738 7239
rect 10766 7266 10794 8302
rect 10934 8329 11074 8330
rect 10934 8303 10935 8329
rect 10961 8303 11074 8329
rect 10934 8302 11074 8303
rect 10934 8297 10962 8302
rect 10990 8050 11018 8055
rect 10990 7769 11018 8022
rect 10990 7743 10991 7769
rect 11017 7743 11018 7769
rect 10990 7737 11018 7743
rect 11046 7938 11074 8302
rect 11046 7713 11074 7910
rect 11942 7882 11970 8471
rect 12054 8441 12082 9198
rect 12110 9179 12138 9198
rect 12110 9058 12138 9063
rect 12166 9058 12194 9422
rect 12222 9226 12250 10066
rect 12334 10009 12362 10015
rect 12334 9983 12335 10009
rect 12361 9983 12362 10009
rect 12278 9897 12306 9903
rect 12278 9871 12279 9897
rect 12305 9871 12306 9897
rect 12278 9450 12306 9871
rect 12334 9618 12362 9983
rect 12334 9585 12362 9590
rect 12390 9562 12418 9567
rect 12390 9515 12418 9534
rect 12278 9417 12306 9422
rect 12222 9193 12250 9198
rect 12446 9170 12474 10066
rect 12614 10010 12642 10066
rect 12614 9963 12642 9982
rect 13006 9673 13034 11103
rect 13062 11130 13090 11159
rect 13230 11186 13258 11887
rect 13958 11522 13986 11527
rect 13230 11153 13258 11158
rect 13342 11298 13370 11303
rect 13342 11185 13370 11270
rect 13958 11297 13986 11494
rect 14070 11521 14098 11942
rect 14294 11578 14322 13231
rect 18830 13370 18858 13375
rect 18830 13145 18858 13342
rect 18830 13119 18831 13145
rect 18857 13119 18858 13145
rect 18830 13113 18858 13119
rect 18942 13090 18970 13511
rect 18942 13057 18970 13062
rect 19950 13426 19978 13431
rect 19950 13089 19978 13398
rect 20006 13146 20034 13567
rect 20006 13113 20034 13118
rect 19950 13063 19951 13089
rect 19977 13063 19978 13089
rect 19950 13057 19978 13063
rect 17598 12950 17730 12955
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17598 12917 17730 12922
rect 17598 12166 17730 12171
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17598 12133 17730 12138
rect 20006 12025 20034 12031
rect 20006 11999 20007 12025
rect 20033 11999 20034 12025
rect 18830 11970 18858 11975
rect 18830 11923 18858 11942
rect 20006 11802 20034 11999
rect 20006 11769 20034 11774
rect 14070 11495 14071 11521
rect 14097 11495 14098 11521
rect 14070 11489 14098 11495
rect 14182 11577 14322 11578
rect 14182 11551 14295 11577
rect 14321 11551 14322 11577
rect 14182 11550 14322 11551
rect 13958 11271 13959 11297
rect 13985 11271 13986 11297
rect 13958 11265 13986 11271
rect 14182 11242 14210 11550
rect 14294 11545 14322 11550
rect 18942 11577 18970 11583
rect 18942 11551 18943 11577
rect 18969 11551 18970 11577
rect 14630 11522 14658 11527
rect 14630 11475 14658 11494
rect 15694 11522 15722 11527
rect 14070 11241 14210 11242
rect 14070 11215 14183 11241
rect 14209 11215 14210 11241
rect 14070 11214 14210 11215
rect 13342 11159 13343 11185
rect 13369 11159 13370 11185
rect 13342 11153 13370 11159
rect 13902 11186 13930 11191
rect 13062 11097 13090 11102
rect 13286 11130 13314 11135
rect 13286 11083 13314 11102
rect 13398 11129 13426 11135
rect 13398 11103 13399 11129
rect 13425 11103 13426 11129
rect 13398 10905 13426 11103
rect 13622 11130 13650 11135
rect 13790 11130 13818 11135
rect 13622 11129 13818 11130
rect 13622 11103 13623 11129
rect 13649 11103 13791 11129
rect 13817 11103 13818 11129
rect 13622 11102 13818 11103
rect 13622 11097 13650 11102
rect 13790 11097 13818 11102
rect 13902 11129 13930 11158
rect 13902 11103 13903 11129
rect 13929 11103 13930 11129
rect 13398 10879 13399 10905
rect 13425 10879 13426 10905
rect 13398 10873 13426 10879
rect 13510 11074 13538 11079
rect 13510 10905 13538 11046
rect 13510 10879 13511 10905
rect 13537 10879 13538 10905
rect 13510 10873 13538 10879
rect 13566 10793 13594 10799
rect 13566 10767 13567 10793
rect 13593 10767 13594 10793
rect 13566 10094 13594 10767
rect 13902 10094 13930 11103
rect 14070 10794 14098 11214
rect 14182 11209 14210 11214
rect 14014 10793 14098 10794
rect 14014 10767 14071 10793
rect 14097 10767 14098 10793
rect 14014 10766 14098 10767
rect 14014 10458 14042 10766
rect 14070 10761 14098 10766
rect 14238 11130 14266 11135
rect 14014 10411 14042 10430
rect 14126 10346 14154 10351
rect 14126 10299 14154 10318
rect 14238 10345 14266 11102
rect 15694 11130 15722 11494
rect 15694 11097 15722 11102
rect 15918 11521 15946 11527
rect 15918 11495 15919 11521
rect 15945 11495 15946 11521
rect 14742 11074 14770 11079
rect 14742 11027 14770 11046
rect 14910 11074 14938 11079
rect 14910 11027 14938 11046
rect 14406 10737 14434 10743
rect 14406 10711 14407 10737
rect 14433 10711 14434 10737
rect 14350 10458 14378 10463
rect 14238 10319 14239 10345
rect 14265 10319 14266 10345
rect 14238 10313 14266 10319
rect 14294 10345 14322 10351
rect 14294 10319 14295 10345
rect 14321 10319 14322 10345
rect 13566 10066 13650 10094
rect 13902 10066 14154 10094
rect 13006 9647 13007 9673
rect 13033 9647 13034 9673
rect 12726 9618 12754 9623
rect 12614 9170 12642 9175
rect 12446 9142 12614 9170
rect 12138 9030 12194 9058
rect 12110 8889 12138 9030
rect 12390 8946 12418 8951
rect 12390 8899 12418 8918
rect 12110 8863 12111 8889
rect 12137 8863 12138 8889
rect 12110 8857 12138 8863
rect 12278 8833 12306 8839
rect 12278 8807 12279 8833
rect 12305 8807 12306 8833
rect 12278 8778 12306 8807
rect 12278 8745 12306 8750
rect 12558 8721 12586 8727
rect 12558 8695 12559 8721
rect 12585 8695 12586 8721
rect 12054 8415 12055 8441
rect 12081 8415 12082 8441
rect 12054 8409 12082 8415
rect 12334 8442 12362 8447
rect 11942 7849 11970 7854
rect 11046 7687 11047 7713
rect 11073 7687 11074 7713
rect 11046 7681 11074 7687
rect 10878 7657 10906 7663
rect 10878 7631 10879 7657
rect 10905 7631 10906 7657
rect 10878 7574 10906 7631
rect 11942 7658 11970 7663
rect 10878 7546 11018 7574
rect 10878 7266 10906 7271
rect 10766 7265 10906 7266
rect 10766 7239 10879 7265
rect 10905 7239 10906 7265
rect 10766 7238 10906 7239
rect 10374 7233 10402 7238
rect 10710 7233 10738 7238
rect 10878 7233 10906 7238
rect 10150 6929 10290 6930
rect 10150 6903 10151 6929
rect 10177 6903 10290 6929
rect 10150 6902 10290 6903
rect 10822 7153 10850 7159
rect 10822 7127 10823 7153
rect 10849 7127 10850 7153
rect 10150 6897 10178 6902
rect 10094 6119 10095 6145
rect 10121 6119 10122 6145
rect 10094 6113 10122 6119
rect 10710 6762 10738 6767
rect 9702 6063 9703 6089
rect 9729 6063 9730 6089
rect 9702 6057 9730 6063
rect 9918 5502 10050 5507
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 9918 5469 10050 5474
rect 9918 4718 10050 4723
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 9918 4685 10050 4690
rect 9918 3934 10050 3939
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 9918 3901 10050 3906
rect 9918 3150 10050 3155
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 9918 3117 10050 3122
rect 9918 2366 10050 2371
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 9918 2333 10050 2338
rect 9366 2058 9394 2063
rect 9366 2011 9394 2030
rect 8974 1751 8975 1777
rect 9001 1751 9002 1777
rect 8974 1745 9002 1751
rect 9310 1833 9338 1839
rect 9310 1807 9311 1833
rect 9337 1807 9338 1833
rect 9310 1694 9338 1807
rect 10710 1777 10738 6734
rect 10822 6034 10850 7127
rect 10990 6762 11018 7546
rect 11942 7265 11970 7630
rect 12334 7658 12362 8414
rect 12558 8050 12586 8695
rect 12614 8554 12642 9142
rect 12726 8889 12754 9590
rect 13006 9506 13034 9647
rect 13622 9673 13650 10066
rect 13622 9647 13623 9673
rect 13649 9647 13650 9673
rect 13230 9618 13258 9623
rect 13230 9571 13258 9590
rect 13454 9617 13482 9623
rect 13454 9591 13455 9617
rect 13481 9591 13482 9617
rect 13006 9473 13034 9478
rect 12726 8863 12727 8889
rect 12753 8863 12754 8889
rect 12726 8857 12754 8863
rect 13062 9282 13090 9287
rect 12838 8833 12866 8839
rect 12838 8807 12839 8833
rect 12865 8807 12866 8833
rect 12838 8778 12866 8807
rect 12838 8745 12866 8750
rect 13006 8778 13034 8783
rect 13006 8721 13034 8750
rect 13006 8695 13007 8721
rect 13033 8695 13034 8721
rect 13006 8689 13034 8695
rect 12614 8521 12642 8526
rect 12726 8050 12754 8055
rect 12558 8049 12754 8050
rect 12558 8023 12727 8049
rect 12753 8023 12754 8049
rect 12558 8022 12754 8023
rect 12726 8017 12754 8022
rect 13062 8049 13090 9254
rect 13398 9170 13426 9175
rect 13454 9170 13482 9591
rect 13622 9618 13650 9647
rect 13622 9585 13650 9590
rect 14126 9617 14154 10066
rect 14294 9674 14322 10319
rect 14294 9641 14322 9646
rect 14350 10065 14378 10430
rect 14406 10094 14434 10711
rect 15470 10737 15498 10743
rect 15470 10711 15471 10737
rect 15497 10711 15498 10737
rect 14574 10458 14602 10463
rect 14574 10401 14602 10430
rect 14574 10375 14575 10401
rect 14601 10375 14602 10401
rect 14574 10369 14602 10375
rect 14910 10402 14938 10407
rect 14406 10066 14546 10094
rect 14350 10039 14351 10065
rect 14377 10039 14378 10065
rect 14126 9591 14127 9617
rect 14153 9591 14154 9617
rect 14126 9585 14154 9591
rect 14294 9561 14322 9567
rect 14294 9535 14295 9561
rect 14321 9535 14322 9561
rect 13846 9505 13874 9511
rect 14014 9506 14042 9511
rect 14238 9506 14266 9511
rect 13846 9479 13847 9505
rect 13873 9479 13874 9505
rect 13846 9338 13874 9479
rect 13734 9310 13846 9338
rect 13426 9142 13482 9170
rect 13678 9169 13706 9175
rect 13678 9143 13679 9169
rect 13705 9143 13706 9169
rect 13398 9137 13426 9142
rect 13174 9114 13202 9119
rect 13174 8833 13202 9086
rect 13174 8807 13175 8833
rect 13201 8807 13202 8833
rect 13174 8801 13202 8807
rect 13342 8946 13370 8951
rect 13342 8833 13370 8918
rect 13678 8946 13706 9143
rect 13678 8913 13706 8918
rect 13342 8807 13343 8833
rect 13369 8807 13370 8833
rect 13342 8801 13370 8807
rect 13678 8834 13706 8839
rect 13734 8834 13762 9310
rect 13846 9305 13874 9310
rect 13902 9505 14042 9506
rect 13902 9479 14015 9505
rect 14041 9479 14042 9505
rect 13902 9478 14042 9479
rect 13902 9282 13930 9478
rect 14014 9473 14042 9478
rect 14070 9505 14266 9506
rect 14070 9479 14239 9505
rect 14265 9479 14266 9505
rect 14070 9478 14266 9479
rect 14070 9338 14098 9478
rect 14238 9473 14266 9478
rect 14294 9450 14322 9535
rect 14294 9417 14322 9422
rect 13902 9249 13930 9254
rect 13958 9310 14098 9338
rect 14294 9338 14322 9343
rect 14350 9338 14378 10039
rect 14518 9617 14546 10066
rect 14686 9674 14714 9679
rect 14714 9646 14826 9674
rect 14686 9641 14714 9646
rect 14518 9591 14519 9617
rect 14545 9591 14546 9617
rect 14518 9585 14546 9591
rect 14798 9617 14826 9646
rect 14798 9591 14799 9617
rect 14825 9591 14826 9617
rect 14798 9585 14826 9591
rect 14686 9562 14714 9567
rect 14686 9515 14714 9534
rect 14910 9561 14938 10374
rect 14966 10346 14994 10351
rect 14966 10299 14994 10318
rect 14910 9535 14911 9561
rect 14937 9535 14938 9561
rect 14910 9529 14938 9535
rect 14966 9562 14994 9567
rect 15134 9562 15162 9567
rect 14966 9561 15162 9562
rect 14966 9535 14967 9561
rect 14993 9535 15135 9561
rect 15161 9535 15162 9561
rect 14966 9534 15162 9535
rect 14630 9506 14658 9511
rect 14630 9459 14658 9478
rect 14294 9337 14378 9338
rect 14294 9311 14295 9337
rect 14321 9311 14378 9337
rect 14294 9310 14378 9311
rect 13678 8833 13762 8834
rect 13678 8807 13679 8833
rect 13705 8807 13762 8833
rect 13678 8806 13762 8807
rect 13678 8801 13706 8806
rect 13230 8778 13258 8783
rect 13230 8731 13258 8750
rect 13958 8778 13986 9310
rect 13734 8442 13762 8447
rect 13062 8023 13063 8049
rect 13089 8023 13090 8049
rect 13062 8017 13090 8023
rect 13622 8414 13734 8442
rect 13510 7993 13538 7999
rect 13510 7967 13511 7993
rect 13537 7967 13538 7993
rect 12334 7625 12362 7630
rect 12614 7938 12642 7943
rect 12614 7574 12642 7910
rect 12838 7938 12866 7943
rect 12838 7891 12866 7910
rect 12894 7937 12922 7943
rect 12894 7911 12895 7937
rect 12921 7911 12922 7937
rect 12726 7882 12754 7887
rect 12670 7658 12698 7663
rect 12670 7611 12698 7630
rect 12726 7574 12754 7854
rect 12894 7770 12922 7911
rect 12950 7938 12978 7943
rect 12950 7891 12978 7910
rect 13454 7938 13482 7943
rect 13454 7891 13482 7910
rect 12894 7742 13034 7770
rect 13006 7713 13034 7742
rect 13006 7687 13007 7713
rect 13033 7687 13034 7713
rect 13006 7681 13034 7687
rect 13510 7714 13538 7967
rect 13510 7681 13538 7686
rect 13622 7658 13650 8414
rect 13734 8395 13762 8414
rect 13958 7994 13986 8750
rect 14070 9226 14098 9231
rect 14294 9226 14322 9310
rect 14070 9225 14322 9226
rect 14070 9199 14071 9225
rect 14097 9199 14322 9225
rect 14070 9198 14322 9199
rect 14686 9282 14714 9287
rect 14014 8722 14042 8727
rect 14014 8050 14042 8694
rect 14070 8442 14098 9198
rect 14630 8834 14658 8839
rect 14630 8777 14658 8806
rect 14686 8833 14714 9254
rect 14966 9282 14994 9534
rect 15134 9529 15162 9534
rect 15302 9562 15330 9567
rect 15302 9515 15330 9534
rect 15190 9506 15218 9511
rect 15190 9459 15218 9478
rect 15470 9506 15498 10711
rect 15694 10738 15722 10743
rect 15918 10738 15946 11495
rect 18830 11466 18858 11471
rect 17598 11382 17730 11387
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17598 11349 17730 11354
rect 18830 11185 18858 11438
rect 18830 11159 18831 11185
rect 18857 11159 18858 11185
rect 18830 11153 18858 11159
rect 18942 11074 18970 11551
rect 20006 11466 20034 11471
rect 20006 11419 20034 11438
rect 20006 11241 20034 11247
rect 20006 11215 20007 11241
rect 20033 11215 20034 11241
rect 20006 11130 20034 11215
rect 20006 11097 20034 11102
rect 18942 11041 18970 11046
rect 15694 10737 15946 10738
rect 15694 10711 15695 10737
rect 15721 10711 15946 10737
rect 15694 10710 15946 10711
rect 15694 10458 15722 10710
rect 17598 10598 17730 10603
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17598 10565 17730 10570
rect 15694 10425 15722 10430
rect 16030 10457 16058 10463
rect 16030 10431 16031 10457
rect 16057 10431 16058 10457
rect 16030 10402 16058 10431
rect 20006 10457 20034 10463
rect 20006 10431 20007 10457
rect 20033 10431 20034 10457
rect 16030 10369 16058 10374
rect 18830 10402 18858 10407
rect 18830 10355 18858 10374
rect 20006 10122 20034 10431
rect 20006 10089 20034 10094
rect 18830 10009 18858 10015
rect 18830 9983 18831 10009
rect 18857 9983 18858 10009
rect 17598 9814 17730 9819
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17598 9781 17730 9786
rect 15470 9473 15498 9478
rect 18830 9506 18858 9983
rect 20006 9897 20034 9903
rect 20006 9871 20007 9897
rect 20033 9871 20034 9897
rect 20006 9786 20034 9871
rect 20006 9753 20034 9758
rect 18830 9473 18858 9478
rect 14966 9249 14994 9254
rect 17598 9030 17730 9035
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17598 8997 17730 9002
rect 20006 8889 20034 8895
rect 20006 8863 20007 8889
rect 20033 8863 20034 8889
rect 14686 8807 14687 8833
rect 14713 8807 14714 8833
rect 14686 8801 14714 8807
rect 15190 8834 15218 8839
rect 14630 8751 14631 8777
rect 14657 8751 14658 8777
rect 14630 8745 14658 8751
rect 14518 8722 14546 8727
rect 14518 8675 14546 8694
rect 14070 8409 14098 8414
rect 14294 8442 14322 8447
rect 14126 8385 14154 8391
rect 14126 8359 14127 8385
rect 14153 8359 14154 8385
rect 14070 8162 14098 8167
rect 14126 8162 14154 8359
rect 14070 8161 14154 8162
rect 14070 8135 14071 8161
rect 14097 8135 14154 8161
rect 14070 8134 14154 8135
rect 14070 8129 14098 8134
rect 14014 8022 14098 8050
rect 13958 7966 14042 7994
rect 14014 7965 14042 7966
rect 14014 7939 14015 7965
rect 14041 7939 14042 7965
rect 14070 7993 14098 8022
rect 14070 7967 14071 7993
rect 14097 7967 14098 7993
rect 14070 7961 14098 7967
rect 14014 7933 14042 7939
rect 14294 7769 14322 8414
rect 15190 8385 15218 8806
rect 18830 8834 18858 8839
rect 18830 8787 18858 8806
rect 15414 8442 15442 8447
rect 15414 8395 15442 8414
rect 20006 8442 20034 8863
rect 20006 8409 20034 8414
rect 15190 8359 15191 8385
rect 15217 8359 15218 8385
rect 15190 8353 15218 8359
rect 17598 8246 17730 8251
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17598 8213 17730 8218
rect 20006 8105 20034 8111
rect 20006 8079 20007 8105
rect 20033 8079 20034 8105
rect 14294 7743 14295 7769
rect 14321 7743 14322 7769
rect 14294 7737 14322 7743
rect 18830 8049 18858 8055
rect 18830 8023 18831 8049
rect 18857 8023 18858 8049
rect 12614 7546 12698 7574
rect 12726 7546 12978 7574
rect 11942 7239 11943 7265
rect 11969 7239 11970 7265
rect 11942 7233 11970 7239
rect 12278 7210 12306 7215
rect 12278 7163 12306 7182
rect 12670 6985 12698 7546
rect 12670 6959 12671 6985
rect 12697 6959 12698 6985
rect 12670 6953 12698 6959
rect 12726 7210 12754 7215
rect 12726 6985 12754 7182
rect 12726 6959 12727 6985
rect 12753 6959 12754 6985
rect 12726 6953 12754 6959
rect 12950 6929 12978 7546
rect 12950 6903 12951 6929
rect 12977 6903 12978 6929
rect 12950 6897 12978 6903
rect 13342 7321 13370 7327
rect 13342 7295 13343 7321
rect 13369 7295 13370 7321
rect 13118 6874 13146 6879
rect 13118 6827 13146 6846
rect 13342 6874 13370 7295
rect 13622 7321 13650 7630
rect 14070 7658 14098 7663
rect 14070 7601 14098 7630
rect 18830 7658 18858 8023
rect 20006 7770 20034 8079
rect 20006 7737 20034 7742
rect 18830 7625 18858 7630
rect 14070 7575 14071 7601
rect 14097 7575 14098 7601
rect 14070 7569 14098 7575
rect 17598 7462 17730 7467
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17598 7429 17730 7434
rect 13622 7295 13623 7321
rect 13649 7295 13650 7321
rect 13622 7289 13650 7295
rect 13342 6841 13370 6846
rect 13678 6874 13706 6879
rect 10990 6729 11018 6734
rect 11214 6817 11242 6823
rect 11214 6791 11215 6817
rect 11241 6791 11242 6817
rect 11214 6762 11242 6791
rect 13006 6817 13034 6823
rect 13006 6791 13007 6817
rect 13033 6791 13034 6817
rect 11214 6729 11242 6734
rect 12782 6762 12810 6767
rect 13006 6762 13034 6791
rect 12782 6761 13034 6762
rect 12782 6735 12783 6761
rect 12809 6735 13034 6761
rect 12782 6734 13034 6735
rect 12782 6729 12810 6734
rect 11158 6034 11186 6039
rect 10822 6033 11186 6034
rect 10822 6007 11159 6033
rect 11185 6007 11186 6033
rect 10822 6006 11186 6007
rect 11102 2169 11130 6006
rect 11158 6001 11186 6006
rect 11102 2143 11103 2169
rect 11129 2143 11130 2169
rect 11102 2137 11130 2143
rect 10710 1751 10711 1777
rect 10737 1751 10738 1777
rect 10710 1745 10738 1751
rect 10766 2058 10794 2063
rect 9086 1666 9338 1694
rect 9086 400 9114 1666
rect 9918 1582 10050 1587
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 9918 1549 10050 1554
rect 10766 400 10794 2030
rect 11382 2058 11410 2063
rect 11382 2011 11410 2030
rect 12782 1833 12810 1839
rect 12782 1807 12783 1833
rect 12809 1807 12810 1833
rect 11214 1666 11242 1671
rect 11102 1665 11242 1666
rect 11102 1639 11215 1665
rect 11241 1639 11242 1665
rect 11102 1638 11242 1639
rect 11102 400 11130 1638
rect 11214 1633 11242 1638
rect 12782 400 12810 1807
rect 13678 1777 13706 6846
rect 17598 6678 17730 6683
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17598 6645 17730 6650
rect 17598 5894 17730 5899
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17598 5861 17730 5866
rect 17598 5110 17730 5115
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17598 5077 17730 5082
rect 17598 4326 17730 4331
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17598 4293 17730 4298
rect 17598 3542 17730 3547
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17598 3509 17730 3514
rect 17598 2758 17730 2763
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17598 2725 17730 2730
rect 17598 1974 17730 1979
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17598 1941 17730 1946
rect 13678 1751 13679 1777
rect 13705 1751 13706 1777
rect 13678 1745 13706 1751
rect 8736 0 8792 400
rect 9072 0 9128 400
rect 10752 0 10808 400
rect 11088 0 11144 400
rect 12768 0 12824 400
<< via2 >>
rect 2238 19221 2266 19222
rect 2238 19195 2239 19221
rect 2239 19195 2265 19221
rect 2265 19195 2266 19221
rect 2238 19194 2266 19195
rect 2290 19221 2318 19222
rect 2290 19195 2291 19221
rect 2291 19195 2317 19221
rect 2317 19195 2318 19221
rect 2290 19194 2318 19195
rect 2342 19221 2370 19222
rect 2342 19195 2343 19221
rect 2343 19195 2369 19221
rect 2369 19195 2370 19221
rect 2342 19194 2370 19195
rect 7686 19137 7714 19138
rect 7686 19111 7687 19137
rect 7687 19111 7713 19137
rect 7713 19111 7714 19137
rect 7686 19110 7714 19111
rect 8078 19110 8106 19138
rect 2238 18437 2266 18438
rect 2238 18411 2239 18437
rect 2239 18411 2265 18437
rect 2265 18411 2266 18437
rect 2238 18410 2266 18411
rect 2290 18437 2318 18438
rect 2290 18411 2291 18437
rect 2291 18411 2317 18437
rect 2317 18411 2318 18437
rect 2290 18410 2318 18411
rect 2342 18437 2370 18438
rect 2342 18411 2343 18437
rect 2343 18411 2369 18437
rect 2369 18411 2370 18437
rect 2342 18410 2370 18411
rect 2238 17653 2266 17654
rect 2238 17627 2239 17653
rect 2239 17627 2265 17653
rect 2265 17627 2266 17653
rect 2238 17626 2266 17627
rect 2290 17653 2318 17654
rect 2290 17627 2291 17653
rect 2291 17627 2317 17653
rect 2317 17627 2318 17653
rect 2290 17626 2318 17627
rect 2342 17653 2370 17654
rect 2342 17627 2343 17653
rect 2343 17627 2369 17653
rect 2369 17627 2370 17653
rect 2342 17626 2370 17627
rect 2238 16869 2266 16870
rect 2238 16843 2239 16869
rect 2239 16843 2265 16869
rect 2265 16843 2266 16869
rect 2238 16842 2266 16843
rect 2290 16869 2318 16870
rect 2290 16843 2291 16869
rect 2291 16843 2317 16869
rect 2317 16843 2318 16869
rect 2290 16842 2318 16843
rect 2342 16869 2370 16870
rect 2342 16843 2343 16869
rect 2343 16843 2369 16869
rect 2369 16843 2370 16869
rect 2342 16842 2370 16843
rect 2238 16085 2266 16086
rect 2238 16059 2239 16085
rect 2239 16059 2265 16085
rect 2265 16059 2266 16085
rect 2238 16058 2266 16059
rect 2290 16085 2318 16086
rect 2290 16059 2291 16085
rect 2291 16059 2317 16085
rect 2317 16059 2318 16085
rect 2290 16058 2318 16059
rect 2342 16085 2370 16086
rect 2342 16059 2343 16085
rect 2343 16059 2369 16085
rect 2369 16059 2370 16085
rect 2342 16058 2370 16059
rect 2238 15301 2266 15302
rect 2238 15275 2239 15301
rect 2239 15275 2265 15301
rect 2265 15275 2266 15301
rect 2238 15274 2266 15275
rect 2290 15301 2318 15302
rect 2290 15275 2291 15301
rect 2291 15275 2317 15301
rect 2317 15275 2318 15301
rect 2290 15274 2318 15275
rect 2342 15301 2370 15302
rect 2342 15275 2343 15301
rect 2343 15275 2369 15301
rect 2369 15275 2370 15301
rect 2342 15274 2370 15275
rect 2238 14517 2266 14518
rect 2238 14491 2239 14517
rect 2239 14491 2265 14517
rect 2265 14491 2266 14517
rect 2238 14490 2266 14491
rect 2290 14517 2318 14518
rect 2290 14491 2291 14517
rect 2291 14491 2317 14517
rect 2317 14491 2318 14517
rect 2290 14490 2318 14491
rect 2342 14517 2370 14518
rect 2342 14491 2343 14517
rect 2343 14491 2369 14517
rect 2369 14491 2370 14517
rect 2342 14490 2370 14491
rect 7350 14014 7378 14042
rect 2238 13733 2266 13734
rect 2238 13707 2239 13733
rect 2239 13707 2265 13733
rect 2265 13707 2266 13733
rect 2238 13706 2266 13707
rect 2290 13733 2318 13734
rect 2290 13707 2291 13733
rect 2291 13707 2317 13733
rect 2317 13707 2318 13733
rect 2290 13706 2318 13707
rect 2342 13733 2370 13734
rect 2342 13707 2343 13733
rect 2343 13707 2369 13733
rect 2369 13707 2370 13733
rect 2342 13706 2370 13707
rect 8750 18718 8778 18746
rect 8414 18326 8442 18354
rect 7966 14014 7994 14042
rect 8694 14041 8722 14042
rect 8694 14015 8695 14041
rect 8695 14015 8721 14041
rect 8721 14015 8722 14041
rect 8694 14014 8722 14015
rect 2086 13454 2114 13482
rect 966 11774 994 11802
rect 966 11465 994 11466
rect 966 11439 967 11465
rect 967 11439 993 11465
rect 993 11439 994 11465
rect 966 11438 994 11439
rect 966 11241 994 11242
rect 966 11215 967 11241
rect 967 11215 993 11241
rect 993 11215 994 11241
rect 966 11214 994 11215
rect 2238 12949 2266 12950
rect 2238 12923 2239 12949
rect 2239 12923 2265 12949
rect 2265 12923 2266 12949
rect 2238 12922 2266 12923
rect 2290 12949 2318 12950
rect 2290 12923 2291 12949
rect 2291 12923 2317 12949
rect 2317 12923 2318 12949
rect 2290 12922 2318 12923
rect 2342 12949 2370 12950
rect 2342 12923 2343 12949
rect 2343 12923 2369 12949
rect 2369 12923 2370 12949
rect 2342 12922 2370 12923
rect 2238 12165 2266 12166
rect 2238 12139 2239 12165
rect 2239 12139 2265 12165
rect 2265 12139 2266 12165
rect 2238 12138 2266 12139
rect 2290 12165 2318 12166
rect 2290 12139 2291 12165
rect 2291 12139 2317 12165
rect 2317 12139 2318 12165
rect 2290 12138 2318 12139
rect 2342 12165 2370 12166
rect 2342 12139 2343 12165
rect 2343 12139 2369 12165
rect 2369 12139 2370 12165
rect 2342 12138 2370 12139
rect 2142 11969 2170 11970
rect 2142 11943 2143 11969
rect 2143 11943 2169 11969
rect 2169 11943 2170 11969
rect 2142 11942 2170 11943
rect 2142 11577 2170 11578
rect 2142 11551 2143 11577
rect 2143 11551 2169 11577
rect 2169 11551 2170 11577
rect 2142 11550 2170 11551
rect 5614 11550 5642 11578
rect 2238 11381 2266 11382
rect 2238 11355 2239 11381
rect 2239 11355 2265 11381
rect 2265 11355 2266 11381
rect 2238 11354 2266 11355
rect 2290 11381 2318 11382
rect 2290 11355 2291 11381
rect 2291 11355 2317 11381
rect 2317 11355 2318 11381
rect 2290 11354 2318 11355
rect 2342 11381 2370 11382
rect 2342 11355 2343 11381
rect 2343 11355 2369 11381
rect 2369 11355 2370 11381
rect 2342 11354 2370 11355
rect 2142 11185 2170 11186
rect 2142 11159 2143 11185
rect 2143 11159 2169 11185
rect 2169 11159 2170 11185
rect 2142 11158 2170 11159
rect 2086 10710 2114 10738
rect 6006 11521 6034 11522
rect 6006 11495 6007 11521
rect 6007 11495 6033 11521
rect 6033 11495 6034 11521
rect 6006 11494 6034 11495
rect 7350 13089 7378 13090
rect 7350 13063 7351 13089
rect 7351 13063 7377 13089
rect 7377 13063 7378 13089
rect 7350 13062 7378 13063
rect 7854 13062 7882 13090
rect 7910 12697 7938 12698
rect 7910 12671 7911 12697
rect 7911 12671 7937 12697
rect 7937 12671 7938 12697
rect 7910 12670 7938 12671
rect 8806 13454 8834 13482
rect 9918 18829 9946 18830
rect 9918 18803 9919 18829
rect 9919 18803 9945 18829
rect 9945 18803 9946 18829
rect 9918 18802 9946 18803
rect 9970 18829 9998 18830
rect 9970 18803 9971 18829
rect 9971 18803 9997 18829
rect 9997 18803 9998 18829
rect 9970 18802 9998 18803
rect 10022 18829 10050 18830
rect 10022 18803 10023 18829
rect 10023 18803 10049 18829
rect 10049 18803 10050 18829
rect 10022 18802 10050 18803
rect 9366 18745 9394 18746
rect 9366 18719 9367 18745
rect 9367 18719 9393 18745
rect 9393 18719 9394 18745
rect 9366 18718 9394 18719
rect 17598 19221 17626 19222
rect 17598 19195 17599 19221
rect 17599 19195 17625 19221
rect 17625 19195 17626 19221
rect 17598 19194 17626 19195
rect 17650 19221 17678 19222
rect 17650 19195 17651 19221
rect 17651 19195 17677 19221
rect 17677 19195 17678 19221
rect 17650 19194 17678 19195
rect 17702 19221 17730 19222
rect 17702 19195 17703 19221
rect 17703 19195 17729 19221
rect 17729 19195 17730 19221
rect 17702 19194 17730 19195
rect 12110 19110 12138 19138
rect 12782 19137 12810 19138
rect 12782 19111 12783 19137
rect 12783 19111 12809 19137
rect 12809 19111 12810 19137
rect 12782 19110 12810 19111
rect 10430 18718 10458 18746
rect 9030 18353 9058 18354
rect 9030 18327 9031 18353
rect 9031 18327 9057 18353
rect 9057 18327 9058 18353
rect 9030 18326 9058 18327
rect 9918 18045 9946 18046
rect 9918 18019 9919 18045
rect 9919 18019 9945 18045
rect 9945 18019 9946 18045
rect 9918 18018 9946 18019
rect 9970 18045 9998 18046
rect 9970 18019 9971 18045
rect 9971 18019 9997 18045
rect 9997 18019 9998 18045
rect 9970 18018 9998 18019
rect 10022 18045 10050 18046
rect 10022 18019 10023 18045
rect 10023 18019 10049 18045
rect 10049 18019 10050 18045
rect 10022 18018 10050 18019
rect 9918 17261 9946 17262
rect 9918 17235 9919 17261
rect 9919 17235 9945 17261
rect 9945 17235 9946 17261
rect 9918 17234 9946 17235
rect 9970 17261 9998 17262
rect 9970 17235 9971 17261
rect 9971 17235 9997 17261
rect 9997 17235 9998 17261
rect 9970 17234 9998 17235
rect 10022 17261 10050 17262
rect 10022 17235 10023 17261
rect 10023 17235 10049 17261
rect 10049 17235 10050 17261
rect 10022 17234 10050 17235
rect 9918 16477 9946 16478
rect 9918 16451 9919 16477
rect 9919 16451 9945 16477
rect 9945 16451 9946 16477
rect 9918 16450 9946 16451
rect 9970 16477 9998 16478
rect 9970 16451 9971 16477
rect 9971 16451 9997 16477
rect 9997 16451 9998 16477
rect 9970 16450 9998 16451
rect 10022 16477 10050 16478
rect 10022 16451 10023 16477
rect 10023 16451 10049 16477
rect 10049 16451 10050 16477
rect 10022 16450 10050 16451
rect 9918 15693 9946 15694
rect 9918 15667 9919 15693
rect 9919 15667 9945 15693
rect 9945 15667 9946 15693
rect 9918 15666 9946 15667
rect 9970 15693 9998 15694
rect 9970 15667 9971 15693
rect 9971 15667 9997 15693
rect 9997 15667 9998 15693
rect 9970 15666 9998 15667
rect 10022 15693 10050 15694
rect 10022 15667 10023 15693
rect 10023 15667 10049 15693
rect 10049 15667 10050 15693
rect 10022 15666 10050 15667
rect 9918 14909 9946 14910
rect 9918 14883 9919 14909
rect 9919 14883 9945 14909
rect 9945 14883 9946 14909
rect 9918 14882 9946 14883
rect 9970 14909 9998 14910
rect 9970 14883 9971 14909
rect 9971 14883 9997 14909
rect 9997 14883 9998 14909
rect 9970 14882 9998 14883
rect 10022 14909 10050 14910
rect 10022 14883 10023 14909
rect 10023 14883 10049 14909
rect 10049 14883 10050 14909
rect 10022 14882 10050 14883
rect 9918 14125 9946 14126
rect 9918 14099 9919 14125
rect 9919 14099 9945 14125
rect 9945 14099 9946 14125
rect 9918 14098 9946 14099
rect 9970 14125 9998 14126
rect 9970 14099 9971 14125
rect 9971 14099 9997 14125
rect 9997 14099 9998 14125
rect 9970 14098 9998 14099
rect 10022 14125 10050 14126
rect 10022 14099 10023 14125
rect 10023 14099 10049 14125
rect 10049 14099 10050 14125
rect 10022 14098 10050 14099
rect 9086 14014 9114 14042
rect 9142 13846 9170 13874
rect 9366 13846 9394 13874
rect 8414 12614 8442 12642
rect 8974 13118 9002 13146
rect 8582 12697 8610 12698
rect 8582 12671 8583 12697
rect 8583 12671 8609 12697
rect 8609 12671 8610 12697
rect 8582 12670 8610 12671
rect 7462 11942 7490 11970
rect 8638 12641 8666 12642
rect 8638 12615 8639 12641
rect 8639 12615 8665 12641
rect 8665 12615 8666 12641
rect 8638 12614 8666 12615
rect 8918 12670 8946 12698
rect 8526 11774 8554 11802
rect 6958 11382 6986 11410
rect 7238 11382 7266 11410
rect 6006 11158 6034 11186
rect 5614 11102 5642 11130
rect 7182 11129 7210 11130
rect 7182 11103 7183 11129
rect 7183 11103 7209 11129
rect 7209 11103 7210 11129
rect 7182 11102 7210 11103
rect 2238 10597 2266 10598
rect 2238 10571 2239 10597
rect 2239 10571 2265 10597
rect 2265 10571 2266 10597
rect 2238 10570 2266 10571
rect 2290 10597 2318 10598
rect 2290 10571 2291 10597
rect 2291 10571 2317 10597
rect 2317 10571 2318 10597
rect 2290 10570 2318 10571
rect 2342 10597 2370 10598
rect 2342 10571 2343 10597
rect 2343 10571 2369 10597
rect 2369 10571 2370 10597
rect 2342 10570 2370 10571
rect 4998 10457 5026 10458
rect 4998 10431 4999 10457
rect 4999 10431 5025 10457
rect 5025 10431 5026 10457
rect 4998 10430 5026 10431
rect 6734 10430 6762 10458
rect 7686 11577 7714 11578
rect 7686 11551 7687 11577
rect 7687 11551 7713 11577
rect 7713 11551 7714 11577
rect 7686 11550 7714 11551
rect 8302 11606 8330 11634
rect 7742 11494 7770 11522
rect 7406 11382 7434 11410
rect 7406 11129 7434 11130
rect 7406 11103 7407 11129
rect 7407 11103 7433 11129
rect 7433 11103 7434 11129
rect 7406 11102 7434 11103
rect 7126 10598 7154 10626
rect 7350 10878 7378 10906
rect 7742 11185 7770 11186
rect 7742 11159 7743 11185
rect 7743 11159 7769 11185
rect 7769 11159 7770 11185
rect 7742 11158 7770 11159
rect 7574 10934 7602 10962
rect 2142 10401 2170 10402
rect 2142 10375 2143 10401
rect 2143 10375 2169 10401
rect 2169 10375 2170 10401
rect 2142 10374 2170 10375
rect 6062 10345 6090 10346
rect 6062 10319 6063 10345
rect 6063 10319 6089 10345
rect 6089 10319 6090 10345
rect 6062 10318 6090 10319
rect 966 10094 994 10122
rect 6678 10345 6706 10346
rect 6678 10319 6679 10345
rect 6679 10319 6705 10345
rect 6705 10319 6706 10345
rect 6678 10318 6706 10319
rect 7406 10486 7434 10514
rect 6566 9953 6594 9954
rect 6566 9927 6567 9953
rect 6567 9927 6593 9953
rect 6593 9927 6594 9953
rect 6566 9926 6594 9927
rect 2238 9813 2266 9814
rect 2238 9787 2239 9813
rect 2239 9787 2265 9813
rect 2265 9787 2266 9813
rect 2238 9786 2266 9787
rect 2290 9813 2318 9814
rect 2290 9787 2291 9813
rect 2291 9787 2317 9813
rect 2317 9787 2318 9813
rect 2290 9786 2318 9787
rect 2342 9813 2370 9814
rect 2342 9787 2343 9813
rect 2343 9787 2369 9813
rect 2369 9787 2370 9813
rect 2342 9786 2370 9787
rect 2238 9029 2266 9030
rect 2238 9003 2239 9029
rect 2239 9003 2265 9029
rect 2265 9003 2266 9029
rect 2238 9002 2266 9003
rect 2290 9029 2318 9030
rect 2290 9003 2291 9029
rect 2291 9003 2317 9029
rect 2317 9003 2318 9029
rect 2290 9002 2318 9003
rect 2342 9029 2370 9030
rect 2342 9003 2343 9029
rect 2343 9003 2369 9029
rect 2369 9003 2370 9029
rect 2342 9002 2370 9003
rect 966 8889 994 8890
rect 966 8863 967 8889
rect 967 8863 993 8889
rect 993 8863 994 8889
rect 966 8862 994 8863
rect 2142 8833 2170 8834
rect 2142 8807 2143 8833
rect 2143 8807 2169 8833
rect 2169 8807 2170 8833
rect 2142 8806 2170 8807
rect 5614 8806 5642 8834
rect 6734 9926 6762 9954
rect 7182 10009 7210 10010
rect 7182 9983 7183 10009
rect 7183 9983 7209 10009
rect 7209 9983 7210 10009
rect 7182 9982 7210 9983
rect 7070 9870 7098 9898
rect 6958 9478 6986 9506
rect 6510 8777 6538 8778
rect 6510 8751 6511 8777
rect 6511 8751 6537 8777
rect 6537 8751 6538 8777
rect 6510 8750 6538 8751
rect 6678 9142 6706 9170
rect 6846 8806 6874 8834
rect 7070 9169 7098 9170
rect 7070 9143 7071 9169
rect 7071 9143 7097 9169
rect 7097 9143 7098 9169
rect 7070 9142 7098 9143
rect 6790 8777 6818 8778
rect 6790 8751 6791 8777
rect 6791 8751 6817 8777
rect 6817 8751 6818 8777
rect 6790 8750 6818 8751
rect 7462 10009 7490 10010
rect 7462 9983 7463 10009
rect 7463 9983 7489 10009
rect 7489 9983 7490 10009
rect 7462 9982 7490 9983
rect 7686 10905 7714 10906
rect 7686 10879 7687 10905
rect 7687 10879 7713 10905
rect 7713 10879 7714 10905
rect 7686 10878 7714 10879
rect 7686 10486 7714 10514
rect 8190 11382 8218 11410
rect 8638 11550 8666 11578
rect 9086 12782 9114 12810
rect 8750 11270 8778 11298
rect 8302 11158 8330 11186
rect 8806 11185 8834 11186
rect 8806 11159 8807 11185
rect 8807 11159 8833 11185
rect 8833 11159 8834 11185
rect 8806 11158 8834 11159
rect 9366 13454 9394 13482
rect 11046 18745 11074 18746
rect 11046 18719 11047 18745
rect 11047 18719 11073 18745
rect 11073 18719 11074 18745
rect 11046 18718 11074 18719
rect 17598 18437 17626 18438
rect 17598 18411 17599 18437
rect 17599 18411 17625 18437
rect 17625 18411 17626 18437
rect 17598 18410 17626 18411
rect 17650 18437 17678 18438
rect 17650 18411 17651 18437
rect 17651 18411 17677 18437
rect 17677 18411 17678 18437
rect 17650 18410 17678 18411
rect 17702 18437 17730 18438
rect 17702 18411 17703 18437
rect 17703 18411 17729 18437
rect 17729 18411 17730 18437
rect 17702 18410 17730 18411
rect 17598 17653 17626 17654
rect 17598 17627 17599 17653
rect 17599 17627 17625 17653
rect 17625 17627 17626 17653
rect 17598 17626 17626 17627
rect 17650 17653 17678 17654
rect 17650 17627 17651 17653
rect 17651 17627 17677 17653
rect 17677 17627 17678 17653
rect 17650 17626 17678 17627
rect 17702 17653 17730 17654
rect 17702 17627 17703 17653
rect 17703 17627 17729 17653
rect 17729 17627 17730 17653
rect 17702 17626 17730 17627
rect 17598 16869 17626 16870
rect 17598 16843 17599 16869
rect 17599 16843 17625 16869
rect 17625 16843 17626 16869
rect 17598 16842 17626 16843
rect 17650 16869 17678 16870
rect 17650 16843 17651 16869
rect 17651 16843 17677 16869
rect 17677 16843 17678 16869
rect 17650 16842 17678 16843
rect 17702 16869 17730 16870
rect 17702 16843 17703 16869
rect 17703 16843 17729 16869
rect 17729 16843 17730 16869
rect 17702 16842 17730 16843
rect 17598 16085 17626 16086
rect 17598 16059 17599 16085
rect 17599 16059 17625 16085
rect 17625 16059 17626 16085
rect 17598 16058 17626 16059
rect 17650 16085 17678 16086
rect 17650 16059 17651 16085
rect 17651 16059 17677 16085
rect 17677 16059 17678 16085
rect 17650 16058 17678 16059
rect 17702 16085 17730 16086
rect 17702 16059 17703 16085
rect 17703 16059 17729 16085
rect 17729 16059 17730 16085
rect 17702 16058 17730 16059
rect 9918 13341 9946 13342
rect 9918 13315 9919 13341
rect 9919 13315 9945 13341
rect 9945 13315 9946 13341
rect 9918 13314 9946 13315
rect 9970 13341 9998 13342
rect 9970 13315 9971 13341
rect 9971 13315 9997 13341
rect 9997 13315 9998 13341
rect 9970 13314 9998 13315
rect 10022 13341 10050 13342
rect 10022 13315 10023 13341
rect 10023 13315 10049 13341
rect 10049 13315 10050 13341
rect 10022 13314 10050 13315
rect 10878 13873 10906 13874
rect 10878 13847 10879 13873
rect 10879 13847 10905 13873
rect 10905 13847 10906 13873
rect 10878 13846 10906 13847
rect 10822 13537 10850 13538
rect 10822 13511 10823 13537
rect 10823 13511 10849 13537
rect 10849 13511 10850 13537
rect 10822 13510 10850 13511
rect 9198 12697 9226 12698
rect 9198 12671 9199 12697
rect 9199 12671 9225 12697
rect 9225 12671 9226 12697
rect 9198 12670 9226 12671
rect 9534 13033 9562 13034
rect 9534 13007 9535 13033
rect 9535 13007 9561 13033
rect 9561 13007 9562 13033
rect 9534 13006 9562 13007
rect 10038 13006 10066 13034
rect 9422 12670 9450 12698
rect 9982 12726 10010 12754
rect 10206 12670 10234 12698
rect 9254 12334 9282 12362
rect 9646 12361 9674 12362
rect 9646 12335 9647 12361
rect 9647 12335 9673 12361
rect 9673 12335 9674 12361
rect 9646 12334 9674 12335
rect 9142 11633 9170 11634
rect 9142 11607 9143 11633
rect 9143 11607 9169 11633
rect 9169 11607 9170 11633
rect 9142 11606 9170 11607
rect 8470 10990 8498 11018
rect 8750 11046 8778 11074
rect 7910 10934 7938 10962
rect 7630 9534 7658 9562
rect 8078 10598 8106 10626
rect 8526 10486 8554 10514
rect 8582 10401 8610 10402
rect 8582 10375 8583 10401
rect 8583 10375 8609 10401
rect 8609 10375 8610 10401
rect 8582 10374 8610 10375
rect 8470 10345 8498 10346
rect 8470 10319 8471 10345
rect 8471 10319 8497 10345
rect 8497 10319 8498 10345
rect 8470 10318 8498 10319
rect 8918 11185 8946 11186
rect 8918 11159 8919 11185
rect 8919 11159 8945 11185
rect 8945 11159 8946 11185
rect 8918 11158 8946 11159
rect 8806 10262 8834 10290
rect 8862 10934 8890 10962
rect 8414 10065 8442 10066
rect 8414 10039 8415 10065
rect 8415 10039 8441 10065
rect 8441 10039 8442 10065
rect 8414 10038 8442 10039
rect 8022 9870 8050 9898
rect 7966 9646 7994 9674
rect 7854 9422 7882 9450
rect 8414 9505 8442 9506
rect 8414 9479 8415 9505
rect 8415 9479 8441 9505
rect 8441 9479 8442 9505
rect 8414 9478 8442 9479
rect 8414 9142 8442 9170
rect 7462 9030 7490 9058
rect 7126 8694 7154 8722
rect 8302 8470 8330 8498
rect 8806 9953 8834 9954
rect 8806 9927 8807 9953
rect 8807 9927 8833 9953
rect 8833 9927 8834 9953
rect 8806 9926 8834 9927
rect 8582 9561 8610 9562
rect 8582 9535 8583 9561
rect 8583 9535 8609 9561
rect 8609 9535 8610 9561
rect 8582 9534 8610 9535
rect 8918 10905 8946 10906
rect 8918 10879 8919 10905
rect 8919 10879 8945 10905
rect 8945 10879 8946 10905
rect 8918 10878 8946 10879
rect 9366 11774 9394 11802
rect 9254 11382 9282 11410
rect 9142 10990 9170 11018
rect 9310 10905 9338 10906
rect 9310 10879 9311 10905
rect 9311 10879 9337 10905
rect 9337 10879 9338 10905
rect 9310 10878 9338 10879
rect 8974 10486 9002 10514
rect 8974 10262 9002 10290
rect 8918 9702 8946 9730
rect 8638 9478 8666 9506
rect 8526 9198 8554 9226
rect 8526 8470 8554 8498
rect 2238 8245 2266 8246
rect 2238 8219 2239 8245
rect 2239 8219 2265 8245
rect 2265 8219 2266 8245
rect 2238 8218 2266 8219
rect 2290 8245 2318 8246
rect 2290 8219 2291 8245
rect 2291 8219 2317 8245
rect 2317 8219 2318 8245
rect 2290 8218 2318 8219
rect 2342 8245 2370 8246
rect 2342 8219 2343 8245
rect 2343 8219 2369 8245
rect 2369 8219 2370 8245
rect 2342 8218 2370 8219
rect 8694 9422 8722 9450
rect 8918 9422 8946 9450
rect 8750 9030 8778 9058
rect 8582 8246 8610 8274
rect 8358 7713 8386 7714
rect 8358 7687 8359 7713
rect 8359 7687 8385 7713
rect 8385 7687 8386 7713
rect 8358 7686 8386 7687
rect 8470 7657 8498 7658
rect 8470 7631 8471 7657
rect 8471 7631 8497 7657
rect 8497 7631 8498 7657
rect 8470 7630 8498 7631
rect 7910 7574 7938 7602
rect 2238 7461 2266 7462
rect 2238 7435 2239 7461
rect 2239 7435 2265 7461
rect 2265 7435 2266 7461
rect 2238 7434 2266 7435
rect 2290 7461 2318 7462
rect 2290 7435 2291 7461
rect 2291 7435 2317 7461
rect 2317 7435 2318 7461
rect 2290 7434 2318 7435
rect 2342 7461 2370 7462
rect 2342 7435 2343 7461
rect 2343 7435 2369 7461
rect 2369 7435 2370 7461
rect 2342 7434 2370 7435
rect 7574 7265 7602 7266
rect 7574 7239 7575 7265
rect 7575 7239 7601 7265
rect 7601 7239 7602 7265
rect 7574 7238 7602 7239
rect 2238 6677 2266 6678
rect 2238 6651 2239 6677
rect 2239 6651 2265 6677
rect 2265 6651 2266 6677
rect 2238 6650 2266 6651
rect 2290 6677 2318 6678
rect 2290 6651 2291 6677
rect 2291 6651 2317 6677
rect 2317 6651 2318 6677
rect 2290 6650 2318 6651
rect 2342 6677 2370 6678
rect 2342 6651 2343 6677
rect 2343 6651 2369 6677
rect 2369 6651 2370 6677
rect 2342 6650 2370 6651
rect 9254 10654 9282 10682
rect 9198 10038 9226 10066
rect 9086 9758 9114 9786
rect 9142 9702 9170 9730
rect 9086 9225 9114 9226
rect 9086 9199 9087 9225
rect 9087 9199 9113 9225
rect 9113 9199 9114 9225
rect 9086 9198 9114 9199
rect 9198 9422 9226 9450
rect 9086 8918 9114 8946
rect 8862 8750 8890 8778
rect 9646 11774 9674 11802
rect 9758 11830 9786 11858
rect 9478 11185 9506 11186
rect 9478 11159 9479 11185
rect 9479 11159 9505 11185
rect 9505 11159 9506 11185
rect 9478 11158 9506 11159
rect 9646 10990 9674 11018
rect 9702 11270 9730 11298
rect 9590 10934 9618 10962
rect 9646 10878 9674 10906
rect 9590 10822 9618 10850
rect 9590 10401 9618 10402
rect 9590 10375 9591 10401
rect 9591 10375 9617 10401
rect 9617 10375 9618 10401
rect 9590 10374 9618 10375
rect 9534 10345 9562 10346
rect 9534 10319 9535 10345
rect 9535 10319 9561 10345
rect 9561 10319 9562 10345
rect 9534 10318 9562 10319
rect 9366 9926 9394 9954
rect 9422 10038 9450 10066
rect 9478 9758 9506 9786
rect 9534 9646 9562 9674
rect 9478 9310 9506 9338
rect 9310 9142 9338 9170
rect 9366 9086 9394 9114
rect 9254 8750 9282 8778
rect 9534 9198 9562 9226
rect 10150 12614 10178 12642
rect 9918 12557 9946 12558
rect 9918 12531 9919 12557
rect 9919 12531 9945 12557
rect 9945 12531 9946 12557
rect 9918 12530 9946 12531
rect 9970 12557 9998 12558
rect 9970 12531 9971 12557
rect 9971 12531 9997 12557
rect 9997 12531 9998 12557
rect 9970 12530 9998 12531
rect 10022 12557 10050 12558
rect 10022 12531 10023 12557
rect 10023 12531 10049 12557
rect 10049 12531 10050 12557
rect 10022 12530 10050 12531
rect 10206 11830 10234 11858
rect 9918 11773 9946 11774
rect 9918 11747 9919 11773
rect 9919 11747 9945 11773
rect 9945 11747 9946 11773
rect 9918 11746 9946 11747
rect 9970 11773 9998 11774
rect 9970 11747 9971 11773
rect 9971 11747 9997 11773
rect 9997 11747 9998 11773
rect 9970 11746 9998 11747
rect 10022 11773 10050 11774
rect 10022 11747 10023 11773
rect 10023 11747 10049 11773
rect 10049 11747 10050 11773
rect 10022 11746 10050 11747
rect 10766 13118 10794 13146
rect 10654 13006 10682 13034
rect 10654 12753 10682 12754
rect 10654 12727 10655 12753
rect 10655 12727 10681 12753
rect 10681 12727 10682 12753
rect 10654 12726 10682 12727
rect 10990 13033 11018 13034
rect 10990 13007 10991 13033
rect 10991 13007 11017 13033
rect 11017 13007 11018 13033
rect 10990 13006 11018 13007
rect 10990 12782 11018 12810
rect 10598 12641 10626 12642
rect 10598 12615 10599 12641
rect 10599 12615 10625 12641
rect 10625 12615 10626 12641
rect 10598 12614 10626 12615
rect 17598 15301 17626 15302
rect 17598 15275 17599 15301
rect 17599 15275 17625 15301
rect 17625 15275 17626 15301
rect 17598 15274 17626 15275
rect 17650 15301 17678 15302
rect 17650 15275 17651 15301
rect 17651 15275 17677 15301
rect 17677 15275 17678 15301
rect 17650 15274 17678 15275
rect 17702 15301 17730 15302
rect 17702 15275 17703 15301
rect 17703 15275 17729 15301
rect 17729 15275 17730 15301
rect 17702 15274 17730 15275
rect 17598 14517 17626 14518
rect 17598 14491 17599 14517
rect 17599 14491 17625 14517
rect 17625 14491 17626 14517
rect 17598 14490 17626 14491
rect 17650 14517 17678 14518
rect 17650 14491 17651 14517
rect 17651 14491 17677 14517
rect 17677 14491 17678 14517
rect 17650 14490 17678 14491
rect 17702 14517 17730 14518
rect 17702 14491 17703 14517
rect 17703 14491 17729 14517
rect 17729 14491 17730 14517
rect 17702 14490 17730 14491
rect 11158 13033 11186 13034
rect 11158 13007 11159 13033
rect 11159 13007 11185 13033
rect 11185 13007 11186 13033
rect 11158 13006 11186 13007
rect 11718 13398 11746 13426
rect 17598 13733 17626 13734
rect 17598 13707 17599 13733
rect 17599 13707 17625 13733
rect 17625 13707 17626 13733
rect 17598 13706 17626 13707
rect 17650 13733 17678 13734
rect 17650 13707 17651 13733
rect 17651 13707 17677 13733
rect 17677 13707 17678 13733
rect 17650 13706 17678 13707
rect 17702 13733 17730 13734
rect 17702 13707 17703 13733
rect 17703 13707 17729 13733
rect 17729 13707 17730 13733
rect 17702 13706 17730 13707
rect 12390 13537 12418 13538
rect 12390 13511 12391 13537
rect 12391 13511 12417 13537
rect 12417 13511 12418 13537
rect 12390 13510 12418 13511
rect 12670 13510 12698 13538
rect 12222 13398 12250 13426
rect 12278 13454 12306 13482
rect 12782 13481 12810 13482
rect 12782 13455 12783 13481
rect 12783 13455 12809 13481
rect 12809 13455 12810 13481
rect 12782 13454 12810 13455
rect 12670 13398 12698 13426
rect 11438 12782 11466 12810
rect 11102 12670 11130 12698
rect 10654 11857 10682 11858
rect 10654 11831 10655 11857
rect 10655 11831 10681 11857
rect 10681 11831 10682 11857
rect 10654 11830 10682 11831
rect 10430 11718 10458 11746
rect 10710 11718 10738 11746
rect 10542 11046 10570 11074
rect 9918 10989 9946 10990
rect 9918 10963 9919 10989
rect 9919 10963 9945 10989
rect 9945 10963 9946 10989
rect 9918 10962 9946 10963
rect 9970 10989 9998 10990
rect 9970 10963 9971 10989
rect 9971 10963 9997 10989
rect 9997 10963 9998 10989
rect 9970 10962 9998 10963
rect 10022 10989 10050 10990
rect 10022 10963 10023 10989
rect 10023 10963 10049 10989
rect 10049 10963 10050 10989
rect 10022 10962 10050 10963
rect 10822 11718 10850 11746
rect 11326 12697 11354 12698
rect 11326 12671 11327 12697
rect 11327 12671 11353 12697
rect 11353 12671 11354 12697
rect 11326 12670 11354 12671
rect 11942 12782 11970 12810
rect 12222 13201 12250 13202
rect 12222 13175 12223 13201
rect 12223 13175 12249 13201
rect 12249 13175 12250 13201
rect 12222 13174 12250 13175
rect 14070 13398 14098 13426
rect 13846 13342 13874 13370
rect 12334 13006 12362 13034
rect 11662 12670 11690 12698
rect 11326 12361 11354 12362
rect 11326 12335 11327 12361
rect 11327 12335 11353 12361
rect 11353 12335 11354 12361
rect 11326 12334 11354 12335
rect 11158 11886 11186 11914
rect 10878 11073 10906 11074
rect 10878 11047 10879 11073
rect 10879 11047 10905 11073
rect 10905 11047 10906 11073
rect 10878 11046 10906 11047
rect 11214 11073 11242 11074
rect 11214 11047 11215 11073
rect 11215 11047 11241 11073
rect 11241 11047 11242 11073
rect 11214 11046 11242 11047
rect 9758 10822 9786 10850
rect 9646 9198 9674 9226
rect 9702 10374 9730 10402
rect 9758 9422 9786 9450
rect 10710 10793 10738 10794
rect 10710 10767 10711 10793
rect 10711 10767 10737 10793
rect 10737 10767 10738 10793
rect 10710 10766 10738 10767
rect 10374 10737 10402 10738
rect 10374 10711 10375 10737
rect 10375 10711 10401 10737
rect 10401 10711 10402 10737
rect 10374 10710 10402 10711
rect 10430 10262 10458 10290
rect 9918 10205 9946 10206
rect 9918 10179 9919 10205
rect 9919 10179 9945 10205
rect 9945 10179 9946 10205
rect 9918 10178 9946 10179
rect 9970 10205 9998 10206
rect 9970 10179 9971 10205
rect 9971 10179 9997 10205
rect 9997 10179 9998 10205
rect 9970 10178 9998 10179
rect 10022 10205 10050 10206
rect 10022 10179 10023 10205
rect 10023 10179 10049 10205
rect 10049 10179 10050 10205
rect 10022 10178 10050 10179
rect 10206 9870 10234 9898
rect 9870 9702 9898 9730
rect 10094 9505 10122 9506
rect 10094 9479 10095 9505
rect 10095 9479 10121 9505
rect 10121 9479 10122 9505
rect 10094 9478 10122 9479
rect 9918 9421 9946 9422
rect 9918 9395 9919 9421
rect 9919 9395 9945 9421
rect 9945 9395 9946 9421
rect 9918 9394 9946 9395
rect 9970 9421 9998 9422
rect 9970 9395 9971 9421
rect 9971 9395 9997 9421
rect 9997 9395 9998 9421
rect 9970 9394 9998 9395
rect 10022 9421 10050 9422
rect 10022 9395 10023 9421
rect 10023 9395 10049 9421
rect 10049 9395 10050 9421
rect 10022 9394 10050 9395
rect 9870 9254 9898 9282
rect 9478 8694 9506 8722
rect 9142 8497 9170 8498
rect 9142 8471 9143 8497
rect 9143 8471 9169 8497
rect 9169 8471 9170 8497
rect 9142 8470 9170 8471
rect 9086 8358 9114 8386
rect 9982 9198 10010 9226
rect 10150 9142 10178 9170
rect 10206 9030 10234 9058
rect 9918 8637 9946 8638
rect 9918 8611 9919 8637
rect 9919 8611 9945 8637
rect 9945 8611 9946 8637
rect 9918 8610 9946 8611
rect 9970 8637 9998 8638
rect 9970 8611 9971 8637
rect 9971 8611 9997 8637
rect 9997 8611 9998 8637
rect 9970 8610 9998 8611
rect 10022 8637 10050 8638
rect 10022 8611 10023 8637
rect 10023 8611 10049 8637
rect 10049 8611 10050 8637
rect 10022 8610 10050 8611
rect 9758 8470 9786 8498
rect 9926 8470 9954 8498
rect 11158 10793 11186 10794
rect 11158 10767 11159 10793
rect 11159 10767 11185 10793
rect 11185 10767 11186 10793
rect 11158 10766 11186 10767
rect 11046 10262 11074 10290
rect 10374 9534 10402 9562
rect 10374 9254 10402 9282
rect 10598 9926 10626 9954
rect 10318 9086 10346 9114
rect 10374 9030 10402 9058
rect 10430 8862 10458 8890
rect 10374 8806 10402 8834
rect 9814 8358 9842 8386
rect 8862 8134 8890 8162
rect 9366 8246 9394 8274
rect 8806 7686 8834 7714
rect 8918 7686 8946 7714
rect 8750 7238 8778 7266
rect 7854 6958 7882 6986
rect 2238 5893 2266 5894
rect 2238 5867 2239 5893
rect 2239 5867 2265 5893
rect 2265 5867 2266 5893
rect 2238 5866 2266 5867
rect 2290 5893 2318 5894
rect 2290 5867 2291 5893
rect 2291 5867 2317 5893
rect 2317 5867 2318 5893
rect 2290 5866 2318 5867
rect 2342 5893 2370 5894
rect 2342 5867 2343 5893
rect 2343 5867 2369 5893
rect 2369 5867 2370 5893
rect 2342 5866 2370 5867
rect 2238 5109 2266 5110
rect 2238 5083 2239 5109
rect 2239 5083 2265 5109
rect 2265 5083 2266 5109
rect 2238 5082 2266 5083
rect 2290 5109 2318 5110
rect 2290 5083 2291 5109
rect 2291 5083 2317 5109
rect 2317 5083 2318 5109
rect 2290 5082 2318 5083
rect 2342 5109 2370 5110
rect 2342 5083 2343 5109
rect 2343 5083 2369 5109
rect 2369 5083 2370 5109
rect 2342 5082 2370 5083
rect 2238 4325 2266 4326
rect 2238 4299 2239 4325
rect 2239 4299 2265 4325
rect 2265 4299 2266 4325
rect 2238 4298 2266 4299
rect 2290 4325 2318 4326
rect 2290 4299 2291 4325
rect 2291 4299 2317 4325
rect 2317 4299 2318 4325
rect 2290 4298 2318 4299
rect 2342 4325 2370 4326
rect 2342 4299 2343 4325
rect 2343 4299 2369 4325
rect 2369 4299 2370 4325
rect 2342 4298 2370 4299
rect 2238 3541 2266 3542
rect 2238 3515 2239 3541
rect 2239 3515 2265 3541
rect 2265 3515 2266 3541
rect 2238 3514 2266 3515
rect 2290 3541 2318 3542
rect 2290 3515 2291 3541
rect 2291 3515 2317 3541
rect 2317 3515 2318 3541
rect 2290 3514 2318 3515
rect 2342 3541 2370 3542
rect 2342 3515 2343 3541
rect 2343 3515 2369 3541
rect 2369 3515 2370 3541
rect 2342 3514 2370 3515
rect 2238 2757 2266 2758
rect 2238 2731 2239 2757
rect 2239 2731 2265 2757
rect 2265 2731 2266 2757
rect 2238 2730 2266 2731
rect 2290 2757 2318 2758
rect 2290 2731 2291 2757
rect 2291 2731 2317 2757
rect 2317 2731 2318 2757
rect 2290 2730 2318 2731
rect 2342 2757 2370 2758
rect 2342 2731 2343 2757
rect 2343 2731 2369 2757
rect 2369 2731 2370 2757
rect 2342 2730 2370 2731
rect 9198 7657 9226 7658
rect 9198 7631 9199 7657
rect 9199 7631 9225 7657
rect 9225 7631 9226 7657
rect 9198 7630 9226 7631
rect 9366 7657 9394 7658
rect 9366 7631 9367 7657
rect 9367 7631 9393 7657
rect 9393 7631 9394 7657
rect 9366 7630 9394 7631
rect 9758 8134 9786 8162
rect 9982 8049 10010 8050
rect 9982 8023 9983 8049
rect 9983 8023 10009 8049
rect 10009 8023 10010 8049
rect 9982 8022 10010 8023
rect 10486 8526 10514 8554
rect 11102 9926 11130 9954
rect 10990 9673 11018 9674
rect 10990 9647 10991 9673
rect 10991 9647 11017 9673
rect 11017 9647 11018 9673
rect 10990 9646 11018 9647
rect 10822 9590 10850 9618
rect 10654 9561 10682 9562
rect 10654 9535 10655 9561
rect 10655 9535 10681 9561
rect 10681 9535 10682 9561
rect 10654 9534 10682 9535
rect 11326 10009 11354 10010
rect 11326 9983 11327 10009
rect 11327 9983 11353 10009
rect 11353 9983 11354 10009
rect 11326 9982 11354 9983
rect 11158 9617 11186 9618
rect 11158 9591 11159 9617
rect 11159 9591 11185 9617
rect 11185 9591 11186 9617
rect 11158 9590 11186 9591
rect 11606 10878 11634 10906
rect 12334 11270 12362 11298
rect 11662 11046 11690 11074
rect 11998 11129 12026 11130
rect 11998 11103 11999 11129
rect 11999 11103 12025 11129
rect 12025 11103 12026 11129
rect 11998 11102 12026 11103
rect 12446 12670 12474 12698
rect 12502 12782 12530 12810
rect 13678 13174 13706 13202
rect 13510 13062 13538 13090
rect 14070 13089 14098 13090
rect 14070 13063 14071 13089
rect 14071 13063 14097 13089
rect 14097 13063 14098 13089
rect 14070 13062 14098 13063
rect 12782 12753 12810 12754
rect 12782 12727 12783 12753
rect 12783 12727 12809 12753
rect 12809 12727 12810 12753
rect 12782 12726 12810 12727
rect 13454 12753 13482 12754
rect 13454 12727 13455 12753
rect 13455 12727 13481 12753
rect 13481 12727 13482 12753
rect 13454 12726 13482 12727
rect 12670 12697 12698 12698
rect 12670 12671 12671 12697
rect 12671 12671 12697 12697
rect 12697 12671 12698 12697
rect 12670 12670 12698 12671
rect 12726 11942 12754 11970
rect 12670 11913 12698 11914
rect 12670 11887 12671 11913
rect 12671 11887 12697 11913
rect 12697 11887 12698 11913
rect 12670 11886 12698 11887
rect 14070 11942 14098 11970
rect 13062 11270 13090 11298
rect 12614 11046 12642 11074
rect 11886 10878 11914 10906
rect 11550 9646 11578 9674
rect 11830 10654 11858 10682
rect 11214 9422 11242 9450
rect 10766 9225 10794 9226
rect 10766 9199 10767 9225
rect 10767 9199 10793 9225
rect 10793 9199 10794 9225
rect 10766 9198 10794 9199
rect 10710 9142 10738 9170
rect 11046 9169 11074 9170
rect 11046 9143 11047 9169
rect 11047 9143 11073 9169
rect 11073 9143 11074 9169
rect 11046 9142 11074 9143
rect 10654 8497 10682 8498
rect 10654 8471 10655 8497
rect 10655 8471 10681 8497
rect 10681 8471 10682 8497
rect 10654 8470 10682 8471
rect 10710 8414 10738 8442
rect 10766 8806 10794 8834
rect 11046 8889 11074 8890
rect 11046 8863 11047 8889
rect 11047 8863 11073 8889
rect 11073 8863 11074 8889
rect 11046 8862 11074 8863
rect 11158 8750 11186 8778
rect 11046 8553 11074 8554
rect 11046 8527 11047 8553
rect 11047 8527 11073 8553
rect 11073 8527 11074 8553
rect 11046 8526 11074 8527
rect 11326 9225 11354 9226
rect 11326 9199 11327 9225
rect 11327 9199 11353 9225
rect 11353 9199 11354 9225
rect 11326 9198 11354 9199
rect 11214 8694 11242 8722
rect 11606 9310 11634 9338
rect 11942 10038 11970 10066
rect 11830 9310 11858 9338
rect 11774 8553 11802 8554
rect 11774 8527 11775 8553
rect 11775 8527 11801 8553
rect 11801 8527 11802 8553
rect 11774 8526 11802 8527
rect 11998 9534 12026 9562
rect 12166 10065 12194 10066
rect 12166 10039 12167 10065
rect 12167 10039 12193 10065
rect 12193 10039 12194 10065
rect 12166 10038 12194 10039
rect 12054 9337 12082 9338
rect 12054 9311 12055 9337
rect 12055 9311 12081 9337
rect 12081 9311 12082 9337
rect 12054 9310 12082 9311
rect 9918 7853 9946 7854
rect 9918 7827 9919 7853
rect 9919 7827 9945 7853
rect 9945 7827 9946 7853
rect 9918 7826 9946 7827
rect 9970 7853 9998 7854
rect 9970 7827 9971 7853
rect 9971 7827 9997 7853
rect 9997 7827 9998 7853
rect 9970 7826 9998 7827
rect 10022 7853 10050 7854
rect 10022 7827 10023 7853
rect 10023 7827 10049 7853
rect 10049 7827 10050 7853
rect 10022 7826 10050 7827
rect 10262 7854 10290 7882
rect 9478 7686 9506 7714
rect 10038 7686 10066 7714
rect 9086 7601 9114 7602
rect 9086 7575 9087 7601
rect 9087 7575 9113 7601
rect 9113 7575 9114 7601
rect 9086 7574 9114 7575
rect 8750 2030 8778 2058
rect 2238 1973 2266 1974
rect 2238 1947 2239 1973
rect 2239 1947 2265 1973
rect 2265 1947 2266 1973
rect 2238 1946 2266 1947
rect 2290 1973 2318 1974
rect 2290 1947 2291 1973
rect 2291 1947 2317 1973
rect 2317 1947 2318 1973
rect 2290 1946 2318 1947
rect 2342 1973 2370 1974
rect 2342 1947 2343 1973
rect 2343 1947 2369 1973
rect 2369 1947 2370 1973
rect 2342 1946 2370 1947
rect 9198 7265 9226 7266
rect 9198 7239 9199 7265
rect 9199 7239 9225 7265
rect 9225 7239 9226 7265
rect 9198 7238 9226 7239
rect 9310 6958 9338 6986
rect 9590 7238 9618 7266
rect 10150 7630 10178 7658
rect 9918 7069 9946 7070
rect 9918 7043 9919 7069
rect 9919 7043 9945 7069
rect 9945 7043 9946 7069
rect 9918 7042 9946 7043
rect 9970 7069 9998 7070
rect 9970 7043 9971 7069
rect 9971 7043 9997 7069
rect 9997 7043 9998 7069
rect 9970 7042 9998 7043
rect 10022 7069 10050 7070
rect 10022 7043 10023 7069
rect 10023 7043 10049 7069
rect 10049 7043 10050 7069
rect 10022 7042 10050 7043
rect 9918 6285 9946 6286
rect 9918 6259 9919 6285
rect 9919 6259 9945 6285
rect 9945 6259 9946 6285
rect 9918 6258 9946 6259
rect 9970 6285 9998 6286
rect 9970 6259 9971 6285
rect 9971 6259 9997 6285
rect 9997 6259 9998 6285
rect 9970 6258 9998 6259
rect 10022 6285 10050 6286
rect 10022 6259 10023 6285
rect 10023 6259 10049 6285
rect 10049 6259 10050 6285
rect 10022 6258 10050 6259
rect 10990 8022 11018 8050
rect 11046 7910 11074 7938
rect 12110 9225 12138 9226
rect 12110 9199 12111 9225
rect 12111 9199 12137 9225
rect 12137 9199 12138 9225
rect 12110 9198 12138 9199
rect 12334 9590 12362 9618
rect 12390 9561 12418 9562
rect 12390 9535 12391 9561
rect 12391 9535 12417 9561
rect 12417 9535 12418 9561
rect 12390 9534 12418 9535
rect 12278 9422 12306 9450
rect 12222 9198 12250 9226
rect 12614 10009 12642 10010
rect 12614 9983 12615 10009
rect 12615 9983 12641 10009
rect 12641 9983 12642 10009
rect 12614 9982 12642 9983
rect 13958 11494 13986 11522
rect 13230 11158 13258 11186
rect 13342 11270 13370 11298
rect 18830 13342 18858 13370
rect 18942 13062 18970 13090
rect 19950 13398 19978 13426
rect 20006 13118 20034 13146
rect 17598 12949 17626 12950
rect 17598 12923 17599 12949
rect 17599 12923 17625 12949
rect 17625 12923 17626 12949
rect 17598 12922 17626 12923
rect 17650 12949 17678 12950
rect 17650 12923 17651 12949
rect 17651 12923 17677 12949
rect 17677 12923 17678 12949
rect 17650 12922 17678 12923
rect 17702 12949 17730 12950
rect 17702 12923 17703 12949
rect 17703 12923 17729 12949
rect 17729 12923 17730 12949
rect 17702 12922 17730 12923
rect 17598 12165 17626 12166
rect 17598 12139 17599 12165
rect 17599 12139 17625 12165
rect 17625 12139 17626 12165
rect 17598 12138 17626 12139
rect 17650 12165 17678 12166
rect 17650 12139 17651 12165
rect 17651 12139 17677 12165
rect 17677 12139 17678 12165
rect 17650 12138 17678 12139
rect 17702 12165 17730 12166
rect 17702 12139 17703 12165
rect 17703 12139 17729 12165
rect 17729 12139 17730 12165
rect 17702 12138 17730 12139
rect 18830 11969 18858 11970
rect 18830 11943 18831 11969
rect 18831 11943 18857 11969
rect 18857 11943 18858 11969
rect 18830 11942 18858 11943
rect 20006 11774 20034 11802
rect 14630 11521 14658 11522
rect 14630 11495 14631 11521
rect 14631 11495 14657 11521
rect 14657 11495 14658 11521
rect 14630 11494 14658 11495
rect 15694 11521 15722 11522
rect 15694 11495 15695 11521
rect 15695 11495 15721 11521
rect 15721 11495 15722 11521
rect 15694 11494 15722 11495
rect 13902 11158 13930 11186
rect 13062 11102 13090 11130
rect 13286 11129 13314 11130
rect 13286 11103 13287 11129
rect 13287 11103 13313 11129
rect 13313 11103 13314 11129
rect 13286 11102 13314 11103
rect 13510 11046 13538 11074
rect 14238 11102 14266 11130
rect 14014 10457 14042 10458
rect 14014 10431 14015 10457
rect 14015 10431 14041 10457
rect 14041 10431 14042 10457
rect 14014 10430 14042 10431
rect 14126 10345 14154 10346
rect 14126 10319 14127 10345
rect 14127 10319 14153 10345
rect 14153 10319 14154 10345
rect 14126 10318 14154 10319
rect 15694 11102 15722 11130
rect 14742 11073 14770 11074
rect 14742 11047 14743 11073
rect 14743 11047 14769 11073
rect 14769 11047 14770 11073
rect 14742 11046 14770 11047
rect 14910 11073 14938 11074
rect 14910 11047 14911 11073
rect 14911 11047 14937 11073
rect 14937 11047 14938 11073
rect 14910 11046 14938 11047
rect 14350 10430 14378 10458
rect 12726 9590 12754 9618
rect 12614 9169 12642 9170
rect 12614 9143 12615 9169
rect 12615 9143 12641 9169
rect 12641 9143 12642 9169
rect 12614 9142 12642 9143
rect 12110 9030 12138 9058
rect 12390 8945 12418 8946
rect 12390 8919 12391 8945
rect 12391 8919 12417 8945
rect 12417 8919 12418 8945
rect 12390 8918 12418 8919
rect 12278 8750 12306 8778
rect 12334 8441 12362 8442
rect 12334 8415 12335 8441
rect 12335 8415 12361 8441
rect 12361 8415 12362 8441
rect 12334 8414 12362 8415
rect 11942 7854 11970 7882
rect 11942 7630 11970 7658
rect 10710 6734 10738 6762
rect 9918 5501 9946 5502
rect 9918 5475 9919 5501
rect 9919 5475 9945 5501
rect 9945 5475 9946 5501
rect 9918 5474 9946 5475
rect 9970 5501 9998 5502
rect 9970 5475 9971 5501
rect 9971 5475 9997 5501
rect 9997 5475 9998 5501
rect 9970 5474 9998 5475
rect 10022 5501 10050 5502
rect 10022 5475 10023 5501
rect 10023 5475 10049 5501
rect 10049 5475 10050 5501
rect 10022 5474 10050 5475
rect 9918 4717 9946 4718
rect 9918 4691 9919 4717
rect 9919 4691 9945 4717
rect 9945 4691 9946 4717
rect 9918 4690 9946 4691
rect 9970 4717 9998 4718
rect 9970 4691 9971 4717
rect 9971 4691 9997 4717
rect 9997 4691 9998 4717
rect 9970 4690 9998 4691
rect 10022 4717 10050 4718
rect 10022 4691 10023 4717
rect 10023 4691 10049 4717
rect 10049 4691 10050 4717
rect 10022 4690 10050 4691
rect 9918 3933 9946 3934
rect 9918 3907 9919 3933
rect 9919 3907 9945 3933
rect 9945 3907 9946 3933
rect 9918 3906 9946 3907
rect 9970 3933 9998 3934
rect 9970 3907 9971 3933
rect 9971 3907 9997 3933
rect 9997 3907 9998 3933
rect 9970 3906 9998 3907
rect 10022 3933 10050 3934
rect 10022 3907 10023 3933
rect 10023 3907 10049 3933
rect 10049 3907 10050 3933
rect 10022 3906 10050 3907
rect 9918 3149 9946 3150
rect 9918 3123 9919 3149
rect 9919 3123 9945 3149
rect 9945 3123 9946 3149
rect 9918 3122 9946 3123
rect 9970 3149 9998 3150
rect 9970 3123 9971 3149
rect 9971 3123 9997 3149
rect 9997 3123 9998 3149
rect 9970 3122 9998 3123
rect 10022 3149 10050 3150
rect 10022 3123 10023 3149
rect 10023 3123 10049 3149
rect 10049 3123 10050 3149
rect 10022 3122 10050 3123
rect 9918 2365 9946 2366
rect 9918 2339 9919 2365
rect 9919 2339 9945 2365
rect 9945 2339 9946 2365
rect 9918 2338 9946 2339
rect 9970 2365 9998 2366
rect 9970 2339 9971 2365
rect 9971 2339 9997 2365
rect 9997 2339 9998 2365
rect 9970 2338 9998 2339
rect 10022 2365 10050 2366
rect 10022 2339 10023 2365
rect 10023 2339 10049 2365
rect 10049 2339 10050 2365
rect 10022 2338 10050 2339
rect 9366 2057 9394 2058
rect 9366 2031 9367 2057
rect 9367 2031 9393 2057
rect 9393 2031 9394 2057
rect 9366 2030 9394 2031
rect 13230 9617 13258 9618
rect 13230 9591 13231 9617
rect 13231 9591 13257 9617
rect 13257 9591 13258 9617
rect 13230 9590 13258 9591
rect 13006 9478 13034 9506
rect 13062 9254 13090 9282
rect 12838 8750 12866 8778
rect 13006 8750 13034 8778
rect 12614 8526 12642 8554
rect 13622 9590 13650 9618
rect 14294 9646 14322 9674
rect 14574 10430 14602 10458
rect 14910 10374 14938 10402
rect 13846 9310 13874 9338
rect 13398 9142 13426 9170
rect 13174 9086 13202 9114
rect 13342 8918 13370 8946
rect 13678 8918 13706 8946
rect 14294 9422 14322 9450
rect 13902 9254 13930 9282
rect 14686 9646 14714 9674
rect 14686 9561 14714 9562
rect 14686 9535 14687 9561
rect 14687 9535 14713 9561
rect 14713 9535 14714 9561
rect 14686 9534 14714 9535
rect 14966 10345 14994 10346
rect 14966 10319 14967 10345
rect 14967 10319 14993 10345
rect 14993 10319 14994 10345
rect 14966 10318 14994 10319
rect 14630 9505 14658 9506
rect 14630 9479 14631 9505
rect 14631 9479 14657 9505
rect 14657 9479 14658 9505
rect 14630 9478 14658 9479
rect 13230 8777 13258 8778
rect 13230 8751 13231 8777
rect 13231 8751 13257 8777
rect 13257 8751 13258 8777
rect 13230 8750 13258 8751
rect 13958 8750 13986 8778
rect 13734 8441 13762 8442
rect 13734 8415 13735 8441
rect 13735 8415 13761 8441
rect 13761 8415 13762 8441
rect 13734 8414 13762 8415
rect 12334 7630 12362 7658
rect 12614 7910 12642 7938
rect 12838 7937 12866 7938
rect 12838 7911 12839 7937
rect 12839 7911 12865 7937
rect 12865 7911 12866 7937
rect 12838 7910 12866 7911
rect 12726 7854 12754 7882
rect 12670 7657 12698 7658
rect 12670 7631 12671 7657
rect 12671 7631 12697 7657
rect 12697 7631 12698 7657
rect 12670 7630 12698 7631
rect 12950 7937 12978 7938
rect 12950 7911 12951 7937
rect 12951 7911 12977 7937
rect 12977 7911 12978 7937
rect 12950 7910 12978 7911
rect 13454 7937 13482 7938
rect 13454 7911 13455 7937
rect 13455 7911 13481 7937
rect 13481 7911 13482 7937
rect 13454 7910 13482 7911
rect 13510 7686 13538 7714
rect 14686 9254 14714 9282
rect 14014 8694 14042 8722
rect 14630 8806 14658 8834
rect 15302 9561 15330 9562
rect 15302 9535 15303 9561
rect 15303 9535 15329 9561
rect 15329 9535 15330 9561
rect 15302 9534 15330 9535
rect 15190 9505 15218 9506
rect 15190 9479 15191 9505
rect 15191 9479 15217 9505
rect 15217 9479 15218 9505
rect 15190 9478 15218 9479
rect 18830 11438 18858 11466
rect 17598 11381 17626 11382
rect 17598 11355 17599 11381
rect 17599 11355 17625 11381
rect 17625 11355 17626 11381
rect 17598 11354 17626 11355
rect 17650 11381 17678 11382
rect 17650 11355 17651 11381
rect 17651 11355 17677 11381
rect 17677 11355 17678 11381
rect 17650 11354 17678 11355
rect 17702 11381 17730 11382
rect 17702 11355 17703 11381
rect 17703 11355 17729 11381
rect 17729 11355 17730 11381
rect 17702 11354 17730 11355
rect 20006 11465 20034 11466
rect 20006 11439 20007 11465
rect 20007 11439 20033 11465
rect 20033 11439 20034 11465
rect 20006 11438 20034 11439
rect 20006 11102 20034 11130
rect 18942 11046 18970 11074
rect 17598 10597 17626 10598
rect 17598 10571 17599 10597
rect 17599 10571 17625 10597
rect 17625 10571 17626 10597
rect 17598 10570 17626 10571
rect 17650 10597 17678 10598
rect 17650 10571 17651 10597
rect 17651 10571 17677 10597
rect 17677 10571 17678 10597
rect 17650 10570 17678 10571
rect 17702 10597 17730 10598
rect 17702 10571 17703 10597
rect 17703 10571 17729 10597
rect 17729 10571 17730 10597
rect 17702 10570 17730 10571
rect 15694 10430 15722 10458
rect 16030 10374 16058 10402
rect 18830 10401 18858 10402
rect 18830 10375 18831 10401
rect 18831 10375 18857 10401
rect 18857 10375 18858 10401
rect 18830 10374 18858 10375
rect 20006 10094 20034 10122
rect 17598 9813 17626 9814
rect 17598 9787 17599 9813
rect 17599 9787 17625 9813
rect 17625 9787 17626 9813
rect 17598 9786 17626 9787
rect 17650 9813 17678 9814
rect 17650 9787 17651 9813
rect 17651 9787 17677 9813
rect 17677 9787 17678 9813
rect 17650 9786 17678 9787
rect 17702 9813 17730 9814
rect 17702 9787 17703 9813
rect 17703 9787 17729 9813
rect 17729 9787 17730 9813
rect 17702 9786 17730 9787
rect 15470 9478 15498 9506
rect 20006 9758 20034 9786
rect 18830 9478 18858 9506
rect 14966 9254 14994 9282
rect 17598 9029 17626 9030
rect 17598 9003 17599 9029
rect 17599 9003 17625 9029
rect 17625 9003 17626 9029
rect 17598 9002 17626 9003
rect 17650 9029 17678 9030
rect 17650 9003 17651 9029
rect 17651 9003 17677 9029
rect 17677 9003 17678 9029
rect 17650 9002 17678 9003
rect 17702 9029 17730 9030
rect 17702 9003 17703 9029
rect 17703 9003 17729 9029
rect 17729 9003 17730 9029
rect 17702 9002 17730 9003
rect 15190 8806 15218 8834
rect 14518 8721 14546 8722
rect 14518 8695 14519 8721
rect 14519 8695 14545 8721
rect 14545 8695 14546 8721
rect 14518 8694 14546 8695
rect 14070 8414 14098 8442
rect 14294 8414 14322 8442
rect 18830 8833 18858 8834
rect 18830 8807 18831 8833
rect 18831 8807 18857 8833
rect 18857 8807 18858 8833
rect 18830 8806 18858 8807
rect 15414 8441 15442 8442
rect 15414 8415 15415 8441
rect 15415 8415 15441 8441
rect 15441 8415 15442 8441
rect 15414 8414 15442 8415
rect 20006 8414 20034 8442
rect 17598 8245 17626 8246
rect 17598 8219 17599 8245
rect 17599 8219 17625 8245
rect 17625 8219 17626 8245
rect 17598 8218 17626 8219
rect 17650 8245 17678 8246
rect 17650 8219 17651 8245
rect 17651 8219 17677 8245
rect 17677 8219 17678 8245
rect 17650 8218 17678 8219
rect 17702 8245 17730 8246
rect 17702 8219 17703 8245
rect 17703 8219 17729 8245
rect 17729 8219 17730 8245
rect 17702 8218 17730 8219
rect 13622 7630 13650 7658
rect 12278 7209 12306 7210
rect 12278 7183 12279 7209
rect 12279 7183 12305 7209
rect 12305 7183 12306 7209
rect 12278 7182 12306 7183
rect 12726 7182 12754 7210
rect 13118 6873 13146 6874
rect 13118 6847 13119 6873
rect 13119 6847 13145 6873
rect 13145 6847 13146 6873
rect 13118 6846 13146 6847
rect 14070 7630 14098 7658
rect 20006 7742 20034 7770
rect 18830 7630 18858 7658
rect 17598 7461 17626 7462
rect 17598 7435 17599 7461
rect 17599 7435 17625 7461
rect 17625 7435 17626 7461
rect 17598 7434 17626 7435
rect 17650 7461 17678 7462
rect 17650 7435 17651 7461
rect 17651 7435 17677 7461
rect 17677 7435 17678 7461
rect 17650 7434 17678 7435
rect 17702 7461 17730 7462
rect 17702 7435 17703 7461
rect 17703 7435 17729 7461
rect 17729 7435 17730 7461
rect 17702 7434 17730 7435
rect 13342 6846 13370 6874
rect 13678 6846 13706 6874
rect 10990 6734 11018 6762
rect 11214 6734 11242 6762
rect 10766 2030 10794 2058
rect 9918 1581 9946 1582
rect 9918 1555 9919 1581
rect 9919 1555 9945 1581
rect 9945 1555 9946 1581
rect 9918 1554 9946 1555
rect 9970 1581 9998 1582
rect 9970 1555 9971 1581
rect 9971 1555 9997 1581
rect 9997 1555 9998 1581
rect 9970 1554 9998 1555
rect 10022 1581 10050 1582
rect 10022 1555 10023 1581
rect 10023 1555 10049 1581
rect 10049 1555 10050 1581
rect 10022 1554 10050 1555
rect 11382 2057 11410 2058
rect 11382 2031 11383 2057
rect 11383 2031 11409 2057
rect 11409 2031 11410 2057
rect 11382 2030 11410 2031
rect 17598 6677 17626 6678
rect 17598 6651 17599 6677
rect 17599 6651 17625 6677
rect 17625 6651 17626 6677
rect 17598 6650 17626 6651
rect 17650 6677 17678 6678
rect 17650 6651 17651 6677
rect 17651 6651 17677 6677
rect 17677 6651 17678 6677
rect 17650 6650 17678 6651
rect 17702 6677 17730 6678
rect 17702 6651 17703 6677
rect 17703 6651 17729 6677
rect 17729 6651 17730 6677
rect 17702 6650 17730 6651
rect 17598 5893 17626 5894
rect 17598 5867 17599 5893
rect 17599 5867 17625 5893
rect 17625 5867 17626 5893
rect 17598 5866 17626 5867
rect 17650 5893 17678 5894
rect 17650 5867 17651 5893
rect 17651 5867 17677 5893
rect 17677 5867 17678 5893
rect 17650 5866 17678 5867
rect 17702 5893 17730 5894
rect 17702 5867 17703 5893
rect 17703 5867 17729 5893
rect 17729 5867 17730 5893
rect 17702 5866 17730 5867
rect 17598 5109 17626 5110
rect 17598 5083 17599 5109
rect 17599 5083 17625 5109
rect 17625 5083 17626 5109
rect 17598 5082 17626 5083
rect 17650 5109 17678 5110
rect 17650 5083 17651 5109
rect 17651 5083 17677 5109
rect 17677 5083 17678 5109
rect 17650 5082 17678 5083
rect 17702 5109 17730 5110
rect 17702 5083 17703 5109
rect 17703 5083 17729 5109
rect 17729 5083 17730 5109
rect 17702 5082 17730 5083
rect 17598 4325 17626 4326
rect 17598 4299 17599 4325
rect 17599 4299 17625 4325
rect 17625 4299 17626 4325
rect 17598 4298 17626 4299
rect 17650 4325 17678 4326
rect 17650 4299 17651 4325
rect 17651 4299 17677 4325
rect 17677 4299 17678 4325
rect 17650 4298 17678 4299
rect 17702 4325 17730 4326
rect 17702 4299 17703 4325
rect 17703 4299 17729 4325
rect 17729 4299 17730 4325
rect 17702 4298 17730 4299
rect 17598 3541 17626 3542
rect 17598 3515 17599 3541
rect 17599 3515 17625 3541
rect 17625 3515 17626 3541
rect 17598 3514 17626 3515
rect 17650 3541 17678 3542
rect 17650 3515 17651 3541
rect 17651 3515 17677 3541
rect 17677 3515 17678 3541
rect 17650 3514 17678 3515
rect 17702 3541 17730 3542
rect 17702 3515 17703 3541
rect 17703 3515 17729 3541
rect 17729 3515 17730 3541
rect 17702 3514 17730 3515
rect 17598 2757 17626 2758
rect 17598 2731 17599 2757
rect 17599 2731 17625 2757
rect 17625 2731 17626 2757
rect 17598 2730 17626 2731
rect 17650 2757 17678 2758
rect 17650 2731 17651 2757
rect 17651 2731 17677 2757
rect 17677 2731 17678 2757
rect 17650 2730 17678 2731
rect 17702 2757 17730 2758
rect 17702 2731 17703 2757
rect 17703 2731 17729 2757
rect 17729 2731 17730 2757
rect 17702 2730 17730 2731
rect 17598 1973 17626 1974
rect 17598 1947 17599 1973
rect 17599 1947 17625 1973
rect 17625 1947 17626 1973
rect 17598 1946 17626 1947
rect 17650 1973 17678 1974
rect 17650 1947 17651 1973
rect 17651 1947 17677 1973
rect 17677 1947 17678 1973
rect 17650 1946 17678 1947
rect 17702 1973 17730 1974
rect 17702 1947 17703 1973
rect 17703 1947 17729 1973
rect 17729 1947 17730 1973
rect 17702 1946 17730 1947
<< metal3 >>
rect 2233 19194 2238 19222
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2370 19194 2375 19222
rect 17593 19194 17598 19222
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17730 19194 17735 19222
rect 7681 19110 7686 19138
rect 7714 19110 8078 19138
rect 8106 19110 8111 19138
rect 12105 19110 12110 19138
rect 12138 19110 12782 19138
rect 12810 19110 12815 19138
rect 9913 18802 9918 18830
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 10050 18802 10055 18830
rect 8745 18718 8750 18746
rect 8778 18718 9366 18746
rect 9394 18718 9399 18746
rect 10425 18718 10430 18746
rect 10458 18718 11046 18746
rect 11074 18718 11079 18746
rect 2233 18410 2238 18438
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2370 18410 2375 18438
rect 17593 18410 17598 18438
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17730 18410 17735 18438
rect 8409 18326 8414 18354
rect 8442 18326 9030 18354
rect 9058 18326 9063 18354
rect 9913 18018 9918 18046
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 10050 18018 10055 18046
rect 2233 17626 2238 17654
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2370 17626 2375 17654
rect 17593 17626 17598 17654
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17730 17626 17735 17654
rect 9913 17234 9918 17262
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 10050 17234 10055 17262
rect 2233 16842 2238 16870
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2370 16842 2375 16870
rect 17593 16842 17598 16870
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17730 16842 17735 16870
rect 9913 16450 9918 16478
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 10050 16450 10055 16478
rect 2233 16058 2238 16086
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2370 16058 2375 16086
rect 17593 16058 17598 16086
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17730 16058 17735 16086
rect 9913 15666 9918 15694
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 10050 15666 10055 15694
rect 2233 15274 2238 15302
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2370 15274 2375 15302
rect 17593 15274 17598 15302
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17730 15274 17735 15302
rect 9913 14882 9918 14910
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 10050 14882 10055 14910
rect 2233 14490 2238 14518
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2370 14490 2375 14518
rect 17593 14490 17598 14518
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17730 14490 17735 14518
rect 9913 14098 9918 14126
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 10050 14098 10055 14126
rect 7345 14014 7350 14042
rect 7378 14014 7966 14042
rect 7994 14014 8694 14042
rect 8722 14014 9086 14042
rect 9114 14014 9119 14042
rect 9137 13846 9142 13874
rect 9170 13846 9366 13874
rect 9394 13846 10878 13874
rect 10906 13846 10911 13874
rect 2233 13706 2238 13734
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2370 13706 2375 13734
rect 17593 13706 17598 13734
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17730 13706 17735 13734
rect 10817 13510 10822 13538
rect 10850 13510 12390 13538
rect 12418 13510 12670 13538
rect 12698 13510 12703 13538
rect 0 13482 400 13496
rect 20600 13482 21000 13496
rect 0 13454 2086 13482
rect 2114 13454 2119 13482
rect 8801 13454 8806 13482
rect 8834 13454 9366 13482
rect 9394 13454 9399 13482
rect 12273 13454 12278 13482
rect 12306 13454 12782 13482
rect 12810 13454 12815 13482
rect 19950 13454 21000 13482
rect 0 13440 400 13454
rect 19950 13426 19978 13454
rect 20600 13440 21000 13454
rect 11713 13398 11718 13426
rect 11746 13398 12222 13426
rect 12250 13398 12255 13426
rect 12665 13398 12670 13426
rect 12698 13398 14070 13426
rect 14098 13398 14103 13426
rect 19945 13398 19950 13426
rect 19978 13398 19983 13426
rect 13841 13342 13846 13370
rect 13874 13342 18830 13370
rect 18858 13342 18863 13370
rect 9913 13314 9918 13342
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 10050 13314 10055 13342
rect 12217 13174 12222 13202
rect 12250 13174 13678 13202
rect 13706 13174 13711 13202
rect 20600 13146 21000 13160
rect 8969 13118 8974 13146
rect 9002 13118 10766 13146
rect 10794 13118 10799 13146
rect 20001 13118 20006 13146
rect 20034 13118 21000 13146
rect 20600 13104 21000 13118
rect 7345 13062 7350 13090
rect 7378 13062 7854 13090
rect 7882 13062 7887 13090
rect 13505 13062 13510 13090
rect 13538 13062 14070 13090
rect 14098 13062 18942 13090
rect 18970 13062 18975 13090
rect 9529 13006 9534 13034
rect 9562 13006 10038 13034
rect 10066 13006 10071 13034
rect 10649 13006 10654 13034
rect 10682 13006 10990 13034
rect 11018 13006 11023 13034
rect 11153 13006 11158 13034
rect 11186 13006 12334 13034
rect 12362 13006 12367 13034
rect 2233 12922 2238 12950
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2370 12922 2375 12950
rect 17593 12922 17598 12950
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17730 12922 17735 12950
rect 9081 12782 9086 12810
rect 9114 12782 10990 12810
rect 11018 12782 11438 12810
rect 11466 12782 11942 12810
rect 11970 12782 12502 12810
rect 12530 12782 12535 12810
rect 9977 12726 9982 12754
rect 10010 12726 10654 12754
rect 10682 12726 10687 12754
rect 12777 12726 12782 12754
rect 12810 12726 13454 12754
rect 13482 12726 13487 12754
rect 7905 12670 7910 12698
rect 7938 12670 8582 12698
rect 8610 12670 8615 12698
rect 8913 12670 8918 12698
rect 8946 12670 9198 12698
rect 9226 12670 9422 12698
rect 9450 12670 9455 12698
rect 10201 12670 10206 12698
rect 10234 12670 11102 12698
rect 11130 12670 11326 12698
rect 11354 12670 11359 12698
rect 11657 12670 11662 12698
rect 11690 12670 12446 12698
rect 12474 12670 12670 12698
rect 12698 12670 12703 12698
rect 8409 12614 8414 12642
rect 8442 12614 8638 12642
rect 8666 12614 8671 12642
rect 10145 12614 10150 12642
rect 10178 12614 10598 12642
rect 10626 12614 10631 12642
rect 9913 12530 9918 12558
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 10050 12530 10055 12558
rect 9249 12334 9254 12362
rect 9282 12334 9646 12362
rect 9674 12334 11326 12362
rect 11354 12334 11359 12362
rect 2233 12138 2238 12166
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2370 12138 2375 12166
rect 17593 12138 17598 12166
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17730 12138 17735 12166
rect 2137 11942 2142 11970
rect 2170 11942 7462 11970
rect 7490 11942 7495 11970
rect 12721 11942 12726 11970
rect 12754 11942 14070 11970
rect 14098 11942 18830 11970
rect 18858 11942 18863 11970
rect 11153 11886 11158 11914
rect 11186 11886 12670 11914
rect 12698 11886 12703 11914
rect 9753 11830 9758 11858
rect 9786 11830 10206 11858
rect 10234 11830 10654 11858
rect 10682 11830 10687 11858
rect 0 11802 400 11816
rect 20600 11802 21000 11816
rect 0 11774 966 11802
rect 994 11774 999 11802
rect 8521 11774 8526 11802
rect 8554 11774 9254 11802
rect 9282 11774 9287 11802
rect 9361 11774 9366 11802
rect 9394 11774 9646 11802
rect 9674 11774 9679 11802
rect 20001 11774 20006 11802
rect 20034 11774 21000 11802
rect 0 11760 400 11774
rect 9913 11746 9918 11774
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 10050 11746 10055 11774
rect 20600 11760 21000 11774
rect 10425 11718 10430 11746
rect 10458 11718 10710 11746
rect 10738 11718 10822 11746
rect 10850 11718 10855 11746
rect 8297 11606 8302 11634
rect 8330 11606 9142 11634
rect 9170 11606 9175 11634
rect 10430 11578 10458 11718
rect 2137 11550 2142 11578
rect 2170 11550 5614 11578
rect 5642 11550 5647 11578
rect 7681 11550 7686 11578
rect 7714 11550 8638 11578
rect 8666 11550 10458 11578
rect 6001 11494 6006 11522
rect 6034 11494 7742 11522
rect 7770 11494 7775 11522
rect 13953 11494 13958 11522
rect 13986 11494 14630 11522
rect 14658 11494 14663 11522
rect 15689 11494 15694 11522
rect 15722 11494 15974 11522
rect 0 11466 400 11480
rect 15946 11466 15974 11494
rect 20600 11466 21000 11480
rect 0 11438 966 11466
rect 994 11438 999 11466
rect 15946 11438 18830 11466
rect 18858 11438 18863 11466
rect 20001 11438 20006 11466
rect 20034 11438 21000 11466
rect 0 11424 400 11438
rect 20600 11424 21000 11438
rect 6953 11382 6958 11410
rect 6986 11382 7238 11410
rect 7266 11382 7406 11410
rect 7434 11382 8190 11410
rect 8218 11382 9254 11410
rect 9282 11382 9287 11410
rect 2233 11354 2238 11382
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2370 11354 2375 11382
rect 17593 11354 17598 11382
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17730 11354 17735 11382
rect 8745 11270 8750 11298
rect 8778 11270 9702 11298
rect 9730 11270 12334 11298
rect 12362 11270 13062 11298
rect 13090 11270 13342 11298
rect 13370 11270 13375 11298
rect 961 11214 966 11242
rect 994 11214 999 11242
rect 0 11130 400 11144
rect 966 11130 994 11214
rect 2137 11158 2142 11186
rect 2170 11158 6006 11186
rect 6034 11158 6039 11186
rect 7737 11158 7742 11186
rect 7770 11158 8302 11186
rect 8330 11158 8335 11186
rect 8801 11158 8806 11186
rect 8834 11158 8839 11186
rect 8913 11158 8918 11186
rect 8946 11158 9478 11186
rect 9506 11158 9511 11186
rect 13225 11158 13230 11186
rect 13258 11158 13902 11186
rect 13930 11158 13935 11186
rect 8806 11130 8834 11158
rect 20600 11130 21000 11144
rect 0 11102 994 11130
rect 5609 11102 5614 11130
rect 5642 11102 7182 11130
rect 7210 11102 7215 11130
rect 7401 11102 7406 11130
rect 7434 11102 8834 11130
rect 11993 11102 11998 11130
rect 12026 11102 13062 11130
rect 13090 11102 13286 11130
rect 13314 11102 14238 11130
rect 14266 11102 14271 11130
rect 14742 11102 15694 11130
rect 15722 11102 15727 11130
rect 20001 11102 20006 11130
rect 20034 11102 21000 11130
rect 0 11088 400 11102
rect 14742 11074 14770 11102
rect 20600 11088 21000 11102
rect 8745 11046 8750 11074
rect 8778 11046 10542 11074
rect 10570 11046 10575 11074
rect 10873 11046 10878 11074
rect 10906 11046 11214 11074
rect 11242 11046 11247 11074
rect 11657 11046 11662 11074
rect 11690 11046 12614 11074
rect 12642 11046 12647 11074
rect 13505 11046 13510 11074
rect 13538 11046 14742 11074
rect 14770 11046 14775 11074
rect 14905 11046 14910 11074
rect 14938 11046 18942 11074
rect 18970 11046 18975 11074
rect 8465 10990 8470 11018
rect 8498 10990 9142 11018
rect 9170 10990 9646 11018
rect 9674 10990 9679 11018
rect 9913 10962 9918 10990
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 10050 10962 10055 10990
rect 7569 10934 7574 10962
rect 7602 10934 7910 10962
rect 7938 10934 7943 10962
rect 8857 10934 8862 10962
rect 8890 10934 9590 10962
rect 9618 10934 9623 10962
rect 7910 10906 7938 10934
rect 7345 10878 7350 10906
rect 7378 10878 7686 10906
rect 7714 10878 7719 10906
rect 7910 10878 8918 10906
rect 8946 10878 8951 10906
rect 9305 10878 9310 10906
rect 9338 10878 9646 10906
rect 9674 10878 11606 10906
rect 11634 10878 11886 10906
rect 11914 10878 11919 10906
rect 9585 10822 9590 10850
rect 9618 10822 9758 10850
rect 9786 10822 9791 10850
rect 10705 10766 10710 10794
rect 10738 10766 11158 10794
rect 11186 10766 11191 10794
rect 2081 10710 2086 10738
rect 2114 10710 10374 10738
rect 10402 10710 10407 10738
rect 9235 10654 9254 10682
rect 9282 10654 9287 10682
rect 10066 10654 11830 10682
rect 11858 10654 11863 10682
rect 10066 10626 10094 10654
rect 7121 10598 7126 10626
rect 7154 10598 8078 10626
rect 8106 10598 10094 10626
rect 2233 10570 2238 10598
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2370 10570 2375 10598
rect 4186 10430 4998 10458
rect 5026 10430 6734 10458
rect 6762 10430 6767 10458
rect 4186 10402 4214 10430
rect 2137 10374 2142 10402
rect 2170 10374 4214 10402
rect 6057 10318 6062 10346
rect 6090 10318 6678 10346
rect 6706 10318 6711 10346
rect 0 10122 400 10136
rect 7126 10122 7154 10598
rect 17593 10570 17598 10598
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17730 10570 17735 10598
rect 7401 10486 7406 10514
rect 7434 10486 7686 10514
rect 7714 10486 8526 10514
rect 8554 10486 8974 10514
rect 9002 10486 9007 10514
rect 14009 10430 14014 10458
rect 14042 10430 14350 10458
rect 14378 10430 14574 10458
rect 14602 10430 15694 10458
rect 15722 10430 15727 10458
rect 8577 10374 8582 10402
rect 8610 10374 9590 10402
rect 9618 10374 9702 10402
rect 9730 10374 9735 10402
rect 14905 10374 14910 10402
rect 14938 10374 16030 10402
rect 16058 10374 18830 10402
rect 18858 10374 18863 10402
rect 8465 10318 8470 10346
rect 8498 10318 9534 10346
rect 9562 10318 9567 10346
rect 14121 10318 14126 10346
rect 14154 10318 14966 10346
rect 14994 10318 14999 10346
rect 8801 10262 8806 10290
rect 8834 10262 8974 10290
rect 9002 10262 9007 10290
rect 10425 10262 10430 10290
rect 10458 10262 11046 10290
rect 11074 10262 11079 10290
rect 9913 10178 9918 10206
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 10050 10178 10055 10206
rect 20600 10122 21000 10136
rect 0 10094 966 10122
rect 994 10094 999 10122
rect 6734 10094 7154 10122
rect 20001 10094 20006 10122
rect 20034 10094 21000 10122
rect 0 10080 400 10094
rect 6734 9954 6762 10094
rect 20600 10080 21000 10094
rect 8409 10038 8414 10066
rect 8442 10038 9198 10066
rect 9226 10038 9422 10066
rect 9450 10038 10094 10066
rect 11937 10038 11942 10066
rect 11970 10038 12166 10066
rect 12194 10038 12199 10066
rect 7177 9982 7182 10010
rect 7210 9982 7462 10010
rect 7490 9982 7495 10010
rect 10066 9954 10094 10038
rect 11321 9982 11326 10010
rect 11354 9982 12614 10010
rect 12642 9982 12647 10010
rect 6561 9926 6566 9954
rect 6594 9926 6734 9954
rect 6762 9926 6767 9954
rect 8801 9926 8806 9954
rect 8834 9926 9366 9954
rect 9394 9926 9399 9954
rect 10066 9926 10598 9954
rect 10626 9926 11102 9954
rect 11130 9926 11135 9954
rect 7065 9870 7070 9898
rect 7098 9870 8022 9898
rect 8050 9870 10206 9898
rect 10234 9870 10239 9898
rect 2233 9786 2238 9814
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2370 9786 2375 9814
rect 17593 9786 17598 9814
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17730 9786 17735 9814
rect 20600 9786 21000 9800
rect 9081 9758 9086 9786
rect 9114 9758 9478 9786
rect 9506 9758 9511 9786
rect 20001 9758 20006 9786
rect 20034 9758 21000 9786
rect 20600 9744 21000 9758
rect 8913 9702 8918 9730
rect 8946 9702 9142 9730
rect 9170 9702 9870 9730
rect 9898 9702 9903 9730
rect 7961 9646 7966 9674
rect 7994 9646 9534 9674
rect 9562 9646 10990 9674
rect 11018 9646 11550 9674
rect 11578 9646 11583 9674
rect 14289 9646 14294 9674
rect 14322 9646 14686 9674
rect 14714 9646 14719 9674
rect 10817 9590 10822 9618
rect 10850 9590 11158 9618
rect 11186 9590 11191 9618
rect 12329 9590 12334 9618
rect 12362 9590 12726 9618
rect 12754 9590 13230 9618
rect 13258 9590 13622 9618
rect 13650 9590 13655 9618
rect 7625 9534 7630 9562
rect 7658 9534 8582 9562
rect 8610 9534 10094 9562
rect 10369 9534 10374 9562
rect 10402 9534 10654 9562
rect 10682 9534 10687 9562
rect 11993 9534 11998 9562
rect 12026 9534 12390 9562
rect 12418 9534 12423 9562
rect 14681 9534 14686 9562
rect 14714 9534 15302 9562
rect 15330 9534 15335 9562
rect 6953 9478 6958 9506
rect 6986 9478 8414 9506
rect 8442 9478 8638 9506
rect 8666 9478 8671 9506
rect 10066 9478 10094 9534
rect 10122 9478 10127 9506
rect 13001 9478 13006 9506
rect 13034 9478 14630 9506
rect 14658 9478 14663 9506
rect 15185 9478 15190 9506
rect 15218 9478 15470 9506
rect 15498 9478 18830 9506
rect 18858 9478 18863 9506
rect 7849 9422 7854 9450
rect 7882 9422 8694 9450
rect 8722 9422 8918 9450
rect 8946 9422 9198 9450
rect 9226 9422 9758 9450
rect 9786 9422 9791 9450
rect 11209 9422 11214 9450
rect 11242 9422 12278 9450
rect 12306 9422 14294 9450
rect 14322 9422 14327 9450
rect 9913 9394 9918 9422
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 10050 9394 10055 9422
rect 9473 9310 9478 9338
rect 9506 9310 11606 9338
rect 11634 9310 11639 9338
rect 11825 9310 11830 9338
rect 11858 9310 12054 9338
rect 12082 9310 13846 9338
rect 13874 9310 13879 9338
rect 9865 9254 9870 9282
rect 9898 9254 10374 9282
rect 10402 9254 10407 9282
rect 10766 9226 10794 9310
rect 13057 9254 13062 9282
rect 13090 9254 13902 9282
rect 13930 9254 14686 9282
rect 14714 9254 14966 9282
rect 14994 9254 14999 9282
rect 8521 9198 8526 9226
rect 8554 9198 9086 9226
rect 9114 9198 9534 9226
rect 9562 9198 9567 9226
rect 9641 9198 9646 9226
rect 9674 9198 9982 9226
rect 10010 9198 10015 9226
rect 10761 9198 10766 9226
rect 10794 9198 10799 9226
rect 11321 9198 11326 9226
rect 11354 9198 12110 9226
rect 12138 9198 12222 9226
rect 12250 9198 12255 9226
rect 6673 9142 6678 9170
rect 6706 9142 7070 9170
rect 7098 9142 7103 9170
rect 8409 9142 8414 9170
rect 8442 9142 9310 9170
rect 9338 9142 9343 9170
rect 10145 9142 10150 9170
rect 10178 9142 10626 9170
rect 10705 9142 10710 9170
rect 10738 9142 11046 9170
rect 11074 9142 11079 9170
rect 12609 9142 12614 9170
rect 12642 9142 13398 9170
rect 13426 9142 13431 9170
rect 10598 9114 10626 9142
rect 9361 9086 9366 9114
rect 9394 9086 10318 9114
rect 10346 9086 10351 9114
rect 10598 9086 13174 9114
rect 13202 9086 13207 9114
rect 7457 9030 7462 9058
rect 7490 9030 8750 9058
rect 8778 9030 10206 9058
rect 10234 9030 10239 9058
rect 10369 9030 10374 9058
rect 10402 9030 12110 9058
rect 12138 9030 12143 9058
rect 2233 9002 2238 9030
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2370 9002 2375 9030
rect 17593 9002 17598 9030
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17730 9002 17735 9030
rect 9081 8918 9086 8946
rect 9114 8918 12390 8946
rect 12418 8918 12423 8946
rect 13337 8918 13342 8946
rect 13370 8918 13678 8946
rect 13706 8918 13711 8946
rect 961 8862 966 8890
rect 994 8862 999 8890
rect 10425 8862 10430 8890
rect 10458 8862 11046 8890
rect 11074 8862 11079 8890
rect 0 8778 400 8792
rect 966 8778 994 8862
rect 2137 8806 2142 8834
rect 2170 8806 5614 8834
rect 5642 8806 6846 8834
rect 6874 8806 6879 8834
rect 10369 8806 10374 8834
rect 10402 8806 10766 8834
rect 10794 8806 10799 8834
rect 14625 8806 14630 8834
rect 14658 8806 15190 8834
rect 15218 8806 18830 8834
rect 18858 8806 18863 8834
rect 0 8750 994 8778
rect 6505 8750 6510 8778
rect 6538 8750 6790 8778
rect 6818 8750 6823 8778
rect 8857 8750 8862 8778
rect 8890 8750 9254 8778
rect 9282 8750 9287 8778
rect 11153 8750 11158 8778
rect 11186 8750 12278 8778
rect 12306 8750 12838 8778
rect 12866 8750 12871 8778
rect 13001 8750 13006 8778
rect 13034 8750 13230 8778
rect 13258 8750 13958 8778
rect 13986 8750 13991 8778
rect 0 8736 400 8750
rect 7121 8694 7126 8722
rect 7154 8694 9478 8722
rect 9506 8694 11214 8722
rect 11242 8694 11247 8722
rect 14009 8694 14014 8722
rect 14042 8694 14518 8722
rect 14546 8694 14551 8722
rect 9913 8610 9918 8638
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 10050 8610 10055 8638
rect 10481 8526 10486 8554
rect 10514 8526 11046 8554
rect 11074 8526 11079 8554
rect 11769 8526 11774 8554
rect 11802 8526 12614 8554
rect 12642 8526 12647 8554
rect 8297 8470 8302 8498
rect 8330 8470 8526 8498
rect 8554 8470 9142 8498
rect 9170 8470 9175 8498
rect 9753 8470 9758 8498
rect 9786 8470 9926 8498
rect 9954 8470 10654 8498
rect 10682 8470 10687 8498
rect 20600 8442 21000 8456
rect 10705 8414 10710 8442
rect 10738 8414 12334 8442
rect 12362 8414 12367 8442
rect 13729 8414 13734 8442
rect 13762 8414 14070 8442
rect 14098 8414 14294 8442
rect 14322 8414 15414 8442
rect 15442 8414 15447 8442
rect 20001 8414 20006 8442
rect 20034 8414 21000 8442
rect 20600 8400 21000 8414
rect 9081 8358 9086 8386
rect 9114 8358 9814 8386
rect 9842 8358 9847 8386
rect 8577 8246 8582 8274
rect 8610 8246 9366 8274
rect 9394 8246 9399 8274
rect 2233 8218 2238 8246
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2370 8218 2375 8246
rect 17593 8218 17598 8246
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17730 8218 17735 8246
rect 8857 8134 8862 8162
rect 8890 8134 9758 8162
rect 9786 8134 9791 8162
rect 9977 8022 9982 8050
rect 10010 8022 10990 8050
rect 11018 8022 11023 8050
rect 11041 7910 11046 7938
rect 11074 7910 12614 7938
rect 12642 7910 12838 7938
rect 12866 7910 12871 7938
rect 12945 7910 12950 7938
rect 12978 7910 13454 7938
rect 13482 7910 13487 7938
rect 10257 7854 10262 7882
rect 10290 7854 11942 7882
rect 11970 7854 12726 7882
rect 12754 7854 12759 7882
rect 9913 7826 9918 7854
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 10050 7826 10055 7854
rect 10262 7714 10290 7854
rect 20600 7770 21000 7784
rect 20001 7742 20006 7770
rect 20034 7742 21000 7770
rect 20600 7728 21000 7742
rect 8353 7686 8358 7714
rect 8386 7686 8806 7714
rect 8834 7686 8839 7714
rect 8913 7686 8918 7714
rect 8946 7686 9478 7714
rect 9506 7686 9511 7714
rect 10033 7686 10038 7714
rect 10066 7686 10290 7714
rect 13505 7686 13510 7714
rect 13538 7686 14098 7714
rect 14070 7658 14098 7686
rect 8465 7630 8470 7658
rect 8498 7630 9198 7658
rect 9226 7630 9231 7658
rect 9361 7630 9366 7658
rect 9394 7630 10150 7658
rect 10178 7630 10183 7658
rect 11937 7630 11942 7658
rect 11970 7630 12334 7658
rect 12362 7630 12670 7658
rect 12698 7630 13622 7658
rect 13650 7630 13655 7658
rect 14065 7630 14070 7658
rect 14098 7630 18830 7658
rect 18858 7630 18863 7658
rect 7905 7574 7910 7602
rect 7938 7574 9086 7602
rect 9114 7574 9119 7602
rect 2233 7434 2238 7462
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2370 7434 2375 7462
rect 17593 7434 17598 7462
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17730 7434 17735 7462
rect 7569 7238 7574 7266
rect 7602 7238 8750 7266
rect 8778 7238 9198 7266
rect 9226 7238 9590 7266
rect 9618 7238 9623 7266
rect 12273 7182 12278 7210
rect 12306 7182 12726 7210
rect 12754 7182 12759 7210
rect 9913 7042 9918 7070
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 10050 7042 10055 7070
rect 7849 6958 7854 6986
rect 7882 6958 9310 6986
rect 9338 6958 9343 6986
rect 13113 6846 13118 6874
rect 13146 6846 13342 6874
rect 13370 6846 13678 6874
rect 13706 6846 13711 6874
rect 10705 6734 10710 6762
rect 10738 6734 10990 6762
rect 11018 6734 11214 6762
rect 11242 6734 11247 6762
rect 2233 6650 2238 6678
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2370 6650 2375 6678
rect 17593 6650 17598 6678
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17730 6650 17735 6678
rect 9913 6258 9918 6286
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 10050 6258 10055 6286
rect 2233 5866 2238 5894
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2370 5866 2375 5894
rect 17593 5866 17598 5894
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17730 5866 17735 5894
rect 9913 5474 9918 5502
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 10050 5474 10055 5502
rect 2233 5082 2238 5110
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2370 5082 2375 5110
rect 17593 5082 17598 5110
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17730 5082 17735 5110
rect 9913 4690 9918 4718
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 10050 4690 10055 4718
rect 2233 4298 2238 4326
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2370 4298 2375 4326
rect 17593 4298 17598 4326
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17730 4298 17735 4326
rect 9913 3906 9918 3934
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 10050 3906 10055 3934
rect 2233 3514 2238 3542
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2370 3514 2375 3542
rect 17593 3514 17598 3542
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17730 3514 17735 3542
rect 9913 3122 9918 3150
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 10050 3122 10055 3150
rect 2233 2730 2238 2758
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2370 2730 2375 2758
rect 17593 2730 17598 2758
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17730 2730 17735 2758
rect 9913 2338 9918 2366
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 10050 2338 10055 2366
rect 8745 2030 8750 2058
rect 8778 2030 9366 2058
rect 9394 2030 9399 2058
rect 10761 2030 10766 2058
rect 10794 2030 11382 2058
rect 11410 2030 11415 2058
rect 2233 1946 2238 1974
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2370 1946 2375 1974
rect 17593 1946 17598 1974
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17730 1946 17735 1974
rect 9913 1554 9918 1582
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 10050 1554 10055 1582
<< via3 >>
rect 2238 19194 2266 19222
rect 2290 19194 2318 19222
rect 2342 19194 2370 19222
rect 17598 19194 17626 19222
rect 17650 19194 17678 19222
rect 17702 19194 17730 19222
rect 9918 18802 9946 18830
rect 9970 18802 9998 18830
rect 10022 18802 10050 18830
rect 2238 18410 2266 18438
rect 2290 18410 2318 18438
rect 2342 18410 2370 18438
rect 17598 18410 17626 18438
rect 17650 18410 17678 18438
rect 17702 18410 17730 18438
rect 9918 18018 9946 18046
rect 9970 18018 9998 18046
rect 10022 18018 10050 18046
rect 2238 17626 2266 17654
rect 2290 17626 2318 17654
rect 2342 17626 2370 17654
rect 17598 17626 17626 17654
rect 17650 17626 17678 17654
rect 17702 17626 17730 17654
rect 9918 17234 9946 17262
rect 9970 17234 9998 17262
rect 10022 17234 10050 17262
rect 2238 16842 2266 16870
rect 2290 16842 2318 16870
rect 2342 16842 2370 16870
rect 17598 16842 17626 16870
rect 17650 16842 17678 16870
rect 17702 16842 17730 16870
rect 9918 16450 9946 16478
rect 9970 16450 9998 16478
rect 10022 16450 10050 16478
rect 2238 16058 2266 16086
rect 2290 16058 2318 16086
rect 2342 16058 2370 16086
rect 17598 16058 17626 16086
rect 17650 16058 17678 16086
rect 17702 16058 17730 16086
rect 9918 15666 9946 15694
rect 9970 15666 9998 15694
rect 10022 15666 10050 15694
rect 2238 15274 2266 15302
rect 2290 15274 2318 15302
rect 2342 15274 2370 15302
rect 17598 15274 17626 15302
rect 17650 15274 17678 15302
rect 17702 15274 17730 15302
rect 9918 14882 9946 14910
rect 9970 14882 9998 14910
rect 10022 14882 10050 14910
rect 2238 14490 2266 14518
rect 2290 14490 2318 14518
rect 2342 14490 2370 14518
rect 17598 14490 17626 14518
rect 17650 14490 17678 14518
rect 17702 14490 17730 14518
rect 9918 14098 9946 14126
rect 9970 14098 9998 14126
rect 10022 14098 10050 14126
rect 2238 13706 2266 13734
rect 2290 13706 2318 13734
rect 2342 13706 2370 13734
rect 17598 13706 17626 13734
rect 17650 13706 17678 13734
rect 17702 13706 17730 13734
rect 9918 13314 9946 13342
rect 9970 13314 9998 13342
rect 10022 13314 10050 13342
rect 2238 12922 2266 12950
rect 2290 12922 2318 12950
rect 2342 12922 2370 12950
rect 17598 12922 17626 12950
rect 17650 12922 17678 12950
rect 17702 12922 17730 12950
rect 9918 12530 9946 12558
rect 9970 12530 9998 12558
rect 10022 12530 10050 12558
rect 2238 12138 2266 12166
rect 2290 12138 2318 12166
rect 2342 12138 2370 12166
rect 17598 12138 17626 12166
rect 17650 12138 17678 12166
rect 17702 12138 17730 12166
rect 9254 11774 9282 11802
rect 9918 11746 9946 11774
rect 9970 11746 9998 11774
rect 10022 11746 10050 11774
rect 2238 11354 2266 11382
rect 2290 11354 2318 11382
rect 2342 11354 2370 11382
rect 17598 11354 17626 11382
rect 17650 11354 17678 11382
rect 17702 11354 17730 11382
rect 9918 10962 9946 10990
rect 9970 10962 9998 10990
rect 10022 10962 10050 10990
rect 9254 10654 9282 10682
rect 2238 10570 2266 10598
rect 2290 10570 2318 10598
rect 2342 10570 2370 10598
rect 17598 10570 17626 10598
rect 17650 10570 17678 10598
rect 17702 10570 17730 10598
rect 9918 10178 9946 10206
rect 9970 10178 9998 10206
rect 10022 10178 10050 10206
rect 2238 9786 2266 9814
rect 2290 9786 2318 9814
rect 2342 9786 2370 9814
rect 17598 9786 17626 9814
rect 17650 9786 17678 9814
rect 17702 9786 17730 9814
rect 9918 9394 9946 9422
rect 9970 9394 9998 9422
rect 10022 9394 10050 9422
rect 2238 9002 2266 9030
rect 2290 9002 2318 9030
rect 2342 9002 2370 9030
rect 17598 9002 17626 9030
rect 17650 9002 17678 9030
rect 17702 9002 17730 9030
rect 9918 8610 9946 8638
rect 9970 8610 9998 8638
rect 10022 8610 10050 8638
rect 2238 8218 2266 8246
rect 2290 8218 2318 8246
rect 2342 8218 2370 8246
rect 17598 8218 17626 8246
rect 17650 8218 17678 8246
rect 17702 8218 17730 8246
rect 9918 7826 9946 7854
rect 9970 7826 9998 7854
rect 10022 7826 10050 7854
rect 2238 7434 2266 7462
rect 2290 7434 2318 7462
rect 2342 7434 2370 7462
rect 17598 7434 17626 7462
rect 17650 7434 17678 7462
rect 17702 7434 17730 7462
rect 9918 7042 9946 7070
rect 9970 7042 9998 7070
rect 10022 7042 10050 7070
rect 2238 6650 2266 6678
rect 2290 6650 2318 6678
rect 2342 6650 2370 6678
rect 17598 6650 17626 6678
rect 17650 6650 17678 6678
rect 17702 6650 17730 6678
rect 9918 6258 9946 6286
rect 9970 6258 9998 6286
rect 10022 6258 10050 6286
rect 2238 5866 2266 5894
rect 2290 5866 2318 5894
rect 2342 5866 2370 5894
rect 17598 5866 17626 5894
rect 17650 5866 17678 5894
rect 17702 5866 17730 5894
rect 9918 5474 9946 5502
rect 9970 5474 9998 5502
rect 10022 5474 10050 5502
rect 2238 5082 2266 5110
rect 2290 5082 2318 5110
rect 2342 5082 2370 5110
rect 17598 5082 17626 5110
rect 17650 5082 17678 5110
rect 17702 5082 17730 5110
rect 9918 4690 9946 4718
rect 9970 4690 9998 4718
rect 10022 4690 10050 4718
rect 2238 4298 2266 4326
rect 2290 4298 2318 4326
rect 2342 4298 2370 4326
rect 17598 4298 17626 4326
rect 17650 4298 17678 4326
rect 17702 4298 17730 4326
rect 9918 3906 9946 3934
rect 9970 3906 9998 3934
rect 10022 3906 10050 3934
rect 2238 3514 2266 3542
rect 2290 3514 2318 3542
rect 2342 3514 2370 3542
rect 17598 3514 17626 3542
rect 17650 3514 17678 3542
rect 17702 3514 17730 3542
rect 9918 3122 9946 3150
rect 9970 3122 9998 3150
rect 10022 3122 10050 3150
rect 2238 2730 2266 2758
rect 2290 2730 2318 2758
rect 2342 2730 2370 2758
rect 17598 2730 17626 2758
rect 17650 2730 17678 2758
rect 17702 2730 17730 2758
rect 9918 2338 9946 2366
rect 9970 2338 9998 2366
rect 10022 2338 10050 2366
rect 2238 1946 2266 1974
rect 2290 1946 2318 1974
rect 2342 1946 2370 1974
rect 17598 1946 17626 1974
rect 17650 1946 17678 1974
rect 17702 1946 17730 1974
rect 9918 1554 9946 1582
rect 9970 1554 9998 1582
rect 10022 1554 10050 1582
<< metal4 >>
rect 2224 19222 2384 19238
rect 2224 19194 2238 19222
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2370 19194 2384 19222
rect 2224 18438 2384 19194
rect 2224 18410 2238 18438
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2370 18410 2384 18438
rect 2224 17654 2384 18410
rect 2224 17626 2238 17654
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2370 17626 2384 17654
rect 2224 16870 2384 17626
rect 2224 16842 2238 16870
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2370 16842 2384 16870
rect 2224 16086 2384 16842
rect 2224 16058 2238 16086
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2370 16058 2384 16086
rect 2224 15302 2384 16058
rect 2224 15274 2238 15302
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2370 15274 2384 15302
rect 2224 14518 2384 15274
rect 2224 14490 2238 14518
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2370 14490 2384 14518
rect 2224 13734 2384 14490
rect 2224 13706 2238 13734
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2370 13706 2384 13734
rect 2224 12950 2384 13706
rect 2224 12922 2238 12950
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2370 12922 2384 12950
rect 2224 12166 2384 12922
rect 2224 12138 2238 12166
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2370 12138 2384 12166
rect 2224 11382 2384 12138
rect 9904 18830 10064 19238
rect 9904 18802 9918 18830
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 10050 18802 10064 18830
rect 9904 18046 10064 18802
rect 9904 18018 9918 18046
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 10050 18018 10064 18046
rect 9904 17262 10064 18018
rect 9904 17234 9918 17262
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 10050 17234 10064 17262
rect 9904 16478 10064 17234
rect 9904 16450 9918 16478
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 10050 16450 10064 16478
rect 9904 15694 10064 16450
rect 9904 15666 9918 15694
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 10050 15666 10064 15694
rect 9904 14910 10064 15666
rect 9904 14882 9918 14910
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 10050 14882 10064 14910
rect 9904 14126 10064 14882
rect 9904 14098 9918 14126
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 10050 14098 10064 14126
rect 9904 13342 10064 14098
rect 9904 13314 9918 13342
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 10050 13314 10064 13342
rect 9904 12558 10064 13314
rect 9904 12530 9918 12558
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 10050 12530 10064 12558
rect 2224 11354 2238 11382
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2370 11354 2384 11382
rect 2224 10598 2384 11354
rect 9254 11802 9282 11807
rect 9254 10682 9282 11774
rect 9254 10649 9282 10654
rect 9904 11774 10064 12530
rect 9904 11746 9918 11774
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 10050 11746 10064 11774
rect 9904 10990 10064 11746
rect 9904 10962 9918 10990
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 10050 10962 10064 10990
rect 2224 10570 2238 10598
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2370 10570 2384 10598
rect 2224 9814 2384 10570
rect 2224 9786 2238 9814
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2370 9786 2384 9814
rect 2224 9030 2384 9786
rect 2224 9002 2238 9030
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2370 9002 2384 9030
rect 2224 8246 2384 9002
rect 2224 8218 2238 8246
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2370 8218 2384 8246
rect 2224 7462 2384 8218
rect 2224 7434 2238 7462
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2370 7434 2384 7462
rect 2224 6678 2384 7434
rect 2224 6650 2238 6678
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2370 6650 2384 6678
rect 2224 5894 2384 6650
rect 2224 5866 2238 5894
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2370 5866 2384 5894
rect 2224 5110 2384 5866
rect 2224 5082 2238 5110
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2370 5082 2384 5110
rect 2224 4326 2384 5082
rect 2224 4298 2238 4326
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2370 4298 2384 4326
rect 2224 3542 2384 4298
rect 2224 3514 2238 3542
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2370 3514 2384 3542
rect 2224 2758 2384 3514
rect 2224 2730 2238 2758
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2370 2730 2384 2758
rect 2224 1974 2384 2730
rect 2224 1946 2238 1974
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2370 1946 2384 1974
rect 2224 1538 2384 1946
rect 9904 10206 10064 10962
rect 9904 10178 9918 10206
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 10050 10178 10064 10206
rect 9904 9422 10064 10178
rect 9904 9394 9918 9422
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 10050 9394 10064 9422
rect 9904 8638 10064 9394
rect 9904 8610 9918 8638
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 10050 8610 10064 8638
rect 9904 7854 10064 8610
rect 9904 7826 9918 7854
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 10050 7826 10064 7854
rect 9904 7070 10064 7826
rect 9904 7042 9918 7070
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 10050 7042 10064 7070
rect 9904 6286 10064 7042
rect 9904 6258 9918 6286
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 10050 6258 10064 6286
rect 9904 5502 10064 6258
rect 9904 5474 9918 5502
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 10050 5474 10064 5502
rect 9904 4718 10064 5474
rect 9904 4690 9918 4718
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 10050 4690 10064 4718
rect 9904 3934 10064 4690
rect 9904 3906 9918 3934
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 10050 3906 10064 3934
rect 9904 3150 10064 3906
rect 9904 3122 9918 3150
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 10050 3122 10064 3150
rect 9904 2366 10064 3122
rect 9904 2338 9918 2366
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 10050 2338 10064 2366
rect 9904 1582 10064 2338
rect 9904 1554 9918 1582
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 10050 1554 10064 1582
rect 9904 1538 10064 1554
rect 17584 19222 17744 19238
rect 17584 19194 17598 19222
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17730 19194 17744 19222
rect 17584 18438 17744 19194
rect 17584 18410 17598 18438
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17730 18410 17744 18438
rect 17584 17654 17744 18410
rect 17584 17626 17598 17654
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17730 17626 17744 17654
rect 17584 16870 17744 17626
rect 17584 16842 17598 16870
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17730 16842 17744 16870
rect 17584 16086 17744 16842
rect 17584 16058 17598 16086
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17730 16058 17744 16086
rect 17584 15302 17744 16058
rect 17584 15274 17598 15302
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17730 15274 17744 15302
rect 17584 14518 17744 15274
rect 17584 14490 17598 14518
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17730 14490 17744 14518
rect 17584 13734 17744 14490
rect 17584 13706 17598 13734
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17730 13706 17744 13734
rect 17584 12950 17744 13706
rect 17584 12922 17598 12950
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17730 12922 17744 12950
rect 17584 12166 17744 12922
rect 17584 12138 17598 12166
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17730 12138 17744 12166
rect 17584 11382 17744 12138
rect 17584 11354 17598 11382
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17730 11354 17744 11382
rect 17584 10598 17744 11354
rect 17584 10570 17598 10598
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17730 10570 17744 10598
rect 17584 9814 17744 10570
rect 17584 9786 17598 9814
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17730 9786 17744 9814
rect 17584 9030 17744 9786
rect 17584 9002 17598 9030
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17730 9002 17744 9030
rect 17584 8246 17744 9002
rect 17584 8218 17598 8246
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17730 8218 17744 8246
rect 17584 7462 17744 8218
rect 17584 7434 17598 7462
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17730 7434 17744 7462
rect 17584 6678 17744 7434
rect 17584 6650 17598 6678
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17730 6650 17744 6678
rect 17584 5894 17744 6650
rect 17584 5866 17598 5894
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17730 5866 17744 5894
rect 17584 5110 17744 5866
rect 17584 5082 17598 5110
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17730 5082 17744 5110
rect 17584 4326 17744 5082
rect 17584 4298 17598 4326
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17730 4298 17744 4326
rect 17584 3542 17744 4298
rect 17584 3514 17598 3542
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17730 3514 17744 3542
rect 17584 2758 17744 3514
rect 17584 2730 17598 2758
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17730 2730 17744 2758
rect 17584 1974 17744 2730
rect 17584 1946 17598 1974
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17730 1946 17744 1974
rect 17584 1538 17744 1946
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _106_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 12208 0 -1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _107_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 12432 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _108_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 12208 0 -1 9408
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _109_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 13776 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _110_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 14784 0 1 8624
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _111_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 13328 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _112_
timestamp 1698175906
transform 1 0 10584 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _113_
timestamp 1698175906
transform -1 0 9856 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _114_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8064 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _115_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10584 0 -1 9408
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _116_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 12656 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _117_
timestamp 1698175906
transform 1 0 13944 0 1 7840
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _118_
timestamp 1698175906
transform -1 0 9968 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _119_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 9408 0 1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _120_
timestamp 1698175906
transform 1 0 8176 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _121_
timestamp 1698175906
transform 1 0 9520 0 -1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _122_
timestamp 1698175906
transform -1 0 11424 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _123_
timestamp 1698175906
transform -1 0 10080 0 -1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _124_
timestamp 1698175906
transform -1 0 9184 0 -1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _125_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 10080 0 1 10976
box -43 -43 771 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _126_
timestamp 1698175906
transform -1 0 11872 0 -1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _127_
timestamp 1698175906
transform -1 0 10976 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _128_
timestamp 1698175906
transform -1 0 10528 0 -1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _129_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9912 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _130_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9352 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _131_
timestamp 1698175906
transform -1 0 9800 0 1 13328
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _132_
timestamp 1698175906
transform 1 0 9072 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _133_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9016 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _134_
timestamp 1698175906
transform -1 0 10024 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _135_
timestamp 1698175906
transform -1 0 11480 0 1 9408
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _136_
timestamp 1698175906
transform 1 0 8904 0 1 9408
box -43 -43 771 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _137_
timestamp 1698175906
transform -1 0 9296 0 1 12544
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _138_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 9128 0 -1 13328
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _139_
timestamp 1698175906
transform -1 0 9016 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _140_
timestamp 1698175906
transform -1 0 8568 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _141_
timestamp 1698175906
transform 1 0 7784 0 -1 10192
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _142_
timestamp 1698175906
transform 1 0 9184 0 -1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _143_
timestamp 1698175906
transform -1 0 10192 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _144_
timestamp 1698175906
transform -1 0 7728 0 -1 10192
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _145_
timestamp 1698175906
transform -1 0 7280 0 -1 10192
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _146_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 9968 0 -1 9408
box -43 -43 771 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _147_
timestamp 1698175906
transform -1 0 12208 0 -1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _148_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 12432 0 -1 10192
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _149_
timestamp 1698175906
transform -1 0 11312 0 -1 8624
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _150_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 10584 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _151_
timestamp 1698175906
transform -1 0 11312 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _152_
timestamp 1698175906
transform 1 0 10024 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _153_
timestamp 1698175906
transform 1 0 13104 0 1 8624
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _154_
timestamp 1698175906
transform -1 0 10808 0 -1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _155_
timestamp 1698175906
transform 1 0 9016 0 -1 8624
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _156_
timestamp 1698175906
transform -1 0 9576 0 -1 8624
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _157_
timestamp 1698175906
transform 1 0 8736 0 1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _158_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8736 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _159_
timestamp 1698175906
transform 1 0 6664 0 -1 10192
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _160_
timestamp 1698175906
transform -1 0 8680 0 1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _161_
timestamp 1698175906
transform -1 0 7728 0 1 10192
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _162_
timestamp 1698175906
transform -1 0 6944 0 1 10192
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _163_
timestamp 1698175906
transform -1 0 12040 0 1 10976
box -43 -43 771 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _164_
timestamp 1698175906
transform -1 0 15064 0 1 9408
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _165_
timestamp 1698175906
transform -1 0 14392 0 1 10192
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _166_
timestamp 1698175906
transform 1 0 8512 0 1 9408
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _167_
timestamp 1698175906
transform 1 0 8232 0 -1 7840
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _168_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9184 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _169_
timestamp 1698175906
transform -1 0 13832 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _170_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 11760 0 -1 10976
box -43 -43 883 435
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _171_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 11536 0 1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _172_
timestamp 1698175906
transform 1 0 8680 0 1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _173_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 13160 0 1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _174_
timestamp 1698175906
transform 1 0 9016 0 -1 11760
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _175_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 12432 0 -1 13328
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _176_
timestamp 1698175906
transform -1 0 13608 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _177_
timestamp 1698175906
transform 1 0 10920 0 -1 13328
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _178_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 12264 0 1 12544
box -43 -43 715 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _179_
timestamp 1698175906
transform -1 0 11816 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _180_
timestamp 1698175906
transform -1 0 11760 0 1 12544
box -43 -43 715 435
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _181_
timestamp 1698175906
transform 1 0 10584 0 1 11760
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _182_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 11088 0 1 12544
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _183_
timestamp 1698175906
transform 1 0 7672 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _184_
timestamp 1698175906
transform -1 0 8064 0 -1 11760
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _185_
timestamp 1698175906
transform -1 0 7616 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _186_
timestamp 1698175906
transform 1 0 8456 0 1 12544
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _187_
timestamp 1698175906
transform -1 0 8008 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _188_
timestamp 1698175906
transform -1 0 14392 0 1 9408
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _189_
timestamp 1698175906
transform -1 0 13664 0 -1 10976
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _190_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 13160 0 1 10976
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _191_
timestamp 1698175906
transform 1 0 13720 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _192_
timestamp 1698175906
transform -1 0 10976 0 1 7056
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _193_
timestamp 1698175906
transform -1 0 10416 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _194_
timestamp 1698175906
transform 1 0 6720 0 1 8624
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _195_
timestamp 1698175906
transform -1 0 7224 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _196_
timestamp 1698175906
transform 1 0 10584 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _197_
timestamp 1698175906
transform 1 0 12880 0 -1 7056
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _198_
timestamp 1698175906
transform -1 0 12880 0 -1 7056
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _199_
timestamp 1698175906
transform -1 0 11144 0 -1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _200_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 10304 0 1 7840
box -43 -43 659 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _201_
timestamp 1698175906
transform -1 0 13608 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _202_
timestamp 1698175906
transform 1 0 12208 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _203_
timestamp 1698175906
transform 1 0 12656 0 1 7840
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _204_
timestamp 1698175906
transform -1 0 7952 0 -1 10976
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _205_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8568 0 1 10976
box -43 -43 659 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _206_
timestamp 1698175906
transform -1 0 7504 0 1 10976
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _207_
timestamp 1698175906
transform -1 0 6888 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _208_
timestamp 1698175906
transform 1 0 12600 0 1 11760
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _209_
timestamp 1698175906
transform 1 0 12880 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _210_
timestamp 1698175906
transform 1 0 15064 0 1 9408
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _211_
timestamp 1698175906
transform -1 0 14784 0 1 9408
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _212_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 13664 0 -1 8624
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _213_
timestamp 1698175906
transform 1 0 9072 0 -1 14112
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _214_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 8904 0 1 13328
box -43 -43 1779 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _215_
timestamp 1698175906
transform 1 0 7000 0 1 8624
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _216_
timestamp 1698175906
transform 1 0 6664 0 1 9408
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _217_
timestamp 1698175906
transform 1 0 10584 0 1 8624
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _218_
timestamp 1698175906
transform -1 0 14168 0 -1 9408
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _219_
timestamp 1698175906
transform 1 0 7448 0 1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _220_
timestamp 1698175906
transform -1 0 6552 0 1 10192
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _221_
timestamp 1698175906
transform 1 0 14504 0 1 10192
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _222_
timestamp 1698175906
transform 1 0 7392 0 1 6272
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _223_
timestamp 1698175906
transform 1 0 12320 0 1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _224_
timestamp 1698175906
transform 1 0 12544 0 -1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _225_
timestamp 1698175906
transform 1 0 10696 0 1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _226_
timestamp 1698175906
transform 1 0 9576 0 -1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _227_
timestamp 1698175906
transform -1 0 7560 0 -1 11760
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _228_
timestamp 1698175906
transform 1 0 6888 0 -1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _229_
timestamp 1698175906
transform 1 0 14168 0 -1 11760
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _230_
timestamp 1698175906
transform 1 0 9632 0 -1 6272
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _231_
timestamp 1698175906
transform -1 0 7168 0 -1 8624
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _232_
timestamp 1698175906
transform 1 0 11816 0 1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _233_
timestamp 1698175906
transform 1 0 9688 0 -1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _234_
timestamp 1698175906
transform 1 0 12544 0 -1 7840
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _235_
timestamp 1698175906
transform -1 0 7168 0 -1 10976
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _236_
timestamp 1698175906
transform 1 0 12544 0 -1 11760
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _237_
timestamp 1698175906
transform 1 0 13944 0 -1 10976
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _238_
timestamp 1698175906
transform -1 0 7728 0 1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _239_
timestamp 1698175906
transform 1 0 14672 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _240_
timestamp 1698175906
transform 1 0 8624 0 -1 14112
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _241_
timestamp 1698175906
transform -1 0 9240 0 1 13328
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__109__I dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 13664 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__159__A2
timestamp 1698175906
transform 1 0 6552 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__194__A2
timestamp 1698175906
transform -1 0 6552 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__206__A2
timestamp 1698175906
transform 1 0 8064 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__212__CLK
timestamp 1698175906
transform 1 0 15400 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__213__CLK
timestamp 1698175906
transform -1 0 10920 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__214__CLK
timestamp 1698175906
transform 1 0 9352 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__215__CLK
timestamp 1698175906
transform 1 0 8736 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__216__CLK
timestamp 1698175906
transform 1 0 8400 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__217__CLK
timestamp 1698175906
transform 1 0 12320 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__218__CLK
timestamp 1698175906
transform 1 0 14280 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__219__CLK
timestamp 1698175906
transform 1 0 9184 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__220__CLK
timestamp 1698175906
transform 1 0 6328 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__221__CLK
timestamp 1698175906
transform 1 0 14000 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__222__CLK
timestamp 1698175906
transform 1 0 9128 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__223__CLK
timestamp 1698175906
transform 1 0 14056 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__224__CLK
timestamp 1698175906
transform 1 0 14280 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__225__CLK
timestamp 1698175906
transform -1 0 12432 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__226__CLK
timestamp 1698175906
transform 1 0 11312 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__227__CLK
timestamp 1698175906
transform 1 0 8176 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__228__CLK
timestamp 1698175906
transform 1 0 9240 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__229__CLK
timestamp 1698175906
transform 1 0 15904 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__230__CLK
timestamp 1698175906
transform 1 0 9520 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__231__CLK
timestamp 1698175906
transform 1 0 7280 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__232__CLK
timestamp 1698175906
transform -1 0 13664 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__233__CLK
timestamp 1698175906
transform 1 0 9576 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__234__CLK
timestamp 1698175906
transform 1 0 14280 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__235__CLK
timestamp 1698175906
transform 1 0 7168 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__236__CLK
timestamp 1698175906
transform 1 0 14168 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__237__CLK
timestamp 1698175906
transform 1 0 15680 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1698175906
transform 1 0 10360 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10584 0 1 10192
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1698175906
transform -1 0 11424 0 -1 10192
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1698175906
transform 1 0 12544 0 -1 10192
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 784 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698175906
transform 1 0 2688 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698175906
transform 1 0 4592 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698175906
transform 1 0 6496 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_138 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8400 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_142 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8624 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_172
timestamp 1698175906
transform 1 0 10304 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_176
timestamp 1698175906
transform 1 0 10528 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_206
timestamp 1698175906
transform 1 0 12208 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_210
timestamp 1698175906
transform 1 0 12432 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_240
timestamp 1698175906
transform 1 0 14112 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_274
timestamp 1698175906
transform 1 0 16016 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_308
timestamp 1698175906
transform 1 0 17920 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_342
timestamp 1698175906
transform 1 0 19824 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_346
timestamp 1698175906
transform 1 0 20048 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_348 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 20160 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 784 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698175906
transform 1 0 4368 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698175906
transform 1 0 4704 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698175906
transform 1 0 8288 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_142
timestamp 1698175906
transform 1 0 8624 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_144
timestamp 1698175906
transform 1 0 8736 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_171 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10248 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_179
timestamp 1698175906
transform 1 0 10696 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_207
timestamp 1698175906
transform 1 0 12264 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_209
timestamp 1698175906
transform 1 0 12376 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_212
timestamp 1698175906
transform 1 0 12544 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_276
timestamp 1698175906
transform 1 0 16128 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_282
timestamp 1698175906
transform 1 0 16464 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_346
timestamp 1698175906
transform 1 0 20048 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_348
timestamp 1698175906
transform 1 0 20160 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698175906
transform 1 0 784 0 1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698175906
transform 1 0 2576 0 1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698175906
transform 1 0 2744 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698175906
transform 1 0 6328 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_107
timestamp 1698175906
transform 1 0 6664 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_171
timestamp 1698175906
transform 1 0 10248 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_177
timestamp 1698175906
transform 1 0 10584 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_241
timestamp 1698175906
transform 1 0 14168 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698175906
transform 1 0 14504 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698175906
transform 1 0 18088 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_317
timestamp 1698175906
transform 1 0 18424 0 1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698175906
transform 1 0 784 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698175906
transform 1 0 4368 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698175906
transform 1 0 4704 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698175906
transform 1 0 8288 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_142
timestamp 1698175906
transform 1 0 8624 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_206
timestamp 1698175906
transform 1 0 12208 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_212
timestamp 1698175906
transform 1 0 12544 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_276
timestamp 1698175906
transform 1 0 16128 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_282
timestamp 1698175906
transform 1 0 16464 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_346
timestamp 1698175906
transform 1 0 20048 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_348
timestamp 1698175906
transform 1 0 20160 0 -1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698175906
transform 1 0 784 0 1 3136
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698175906
transform 1 0 2576 0 1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698175906
transform 1 0 2744 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698175906
transform 1 0 6328 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_107
timestamp 1698175906
transform 1 0 6664 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698175906
transform 1 0 10248 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_177
timestamp 1698175906
transform 1 0 10584 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_241
timestamp 1698175906
transform 1 0 14168 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698175906
transform 1 0 14504 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698175906
transform 1 0 18088 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_317
timestamp 1698175906
transform 1 0 18424 0 1 3136
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698175906
transform 1 0 784 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698175906
transform 1 0 4368 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698175906
transform 1 0 4704 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698175906
transform 1 0 8288 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_142
timestamp 1698175906
transform 1 0 8624 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_206
timestamp 1698175906
transform 1 0 12208 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_212
timestamp 1698175906
transform 1 0 12544 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698175906
transform 1 0 16128 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_282
timestamp 1698175906
transform 1 0 16464 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_346
timestamp 1698175906
transform 1 0 20048 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_348
timestamp 1698175906
transform 1 0 20160 0 -1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698175906
transform 1 0 784 0 1 3920
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698175906
transform 1 0 2576 0 1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698175906
transform 1 0 2744 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698175906
transform 1 0 6328 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_107
timestamp 1698175906
transform 1 0 6664 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_171
timestamp 1698175906
transform 1 0 10248 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_177
timestamp 1698175906
transform 1 0 10584 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_241
timestamp 1698175906
transform 1 0 14168 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_247
timestamp 1698175906
transform 1 0 14504 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_311
timestamp 1698175906
transform 1 0 18088 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_317
timestamp 1698175906
transform 1 0 18424 0 1 3920
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698175906
transform 1 0 784 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698175906
transform 1 0 4368 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_72
timestamp 1698175906
transform 1 0 4704 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698175906
transform 1 0 8288 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_142
timestamp 1698175906
transform 1 0 8624 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_206
timestamp 1698175906
transform 1 0 12208 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_212
timestamp 1698175906
transform 1 0 12544 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_276
timestamp 1698175906
transform 1 0 16128 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_282
timestamp 1698175906
transform 1 0 16464 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_346
timestamp 1698175906
transform 1 0 20048 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_348
timestamp 1698175906
transform 1 0 20160 0 -1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698175906
transform 1 0 784 0 1 4704
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698175906
transform 1 0 2576 0 1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_37
timestamp 1698175906
transform 1 0 2744 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_101
timestamp 1698175906
transform 1 0 6328 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_107
timestamp 1698175906
transform 1 0 6664 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_171
timestamp 1698175906
transform 1 0 10248 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_177
timestamp 1698175906
transform 1 0 10584 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_241
timestamp 1698175906
transform 1 0 14168 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_247
timestamp 1698175906
transform 1 0 14504 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_311
timestamp 1698175906
transform 1 0 18088 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_317
timestamp 1698175906
transform 1 0 18424 0 1 4704
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698175906
transform 1 0 784 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698175906
transform 1 0 4368 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_72
timestamp 1698175906
transform 1 0 4704 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_136
timestamp 1698175906
transform 1 0 8288 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_142
timestamp 1698175906
transform 1 0 8624 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_206
timestamp 1698175906
transform 1 0 12208 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_212
timestamp 1698175906
transform 1 0 12544 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_276
timestamp 1698175906
transform 1 0 16128 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_282
timestamp 1698175906
transform 1 0 16464 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_346
timestamp 1698175906
transform 1 0 20048 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_348
timestamp 1698175906
transform 1 0 20160 0 -1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698175906
transform 1 0 784 0 1 5488
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698175906
transform 1 0 2576 0 1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_37
timestamp 1698175906
transform 1 0 2744 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698175906
transform 1 0 6328 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_107
timestamp 1698175906
transform 1 0 6664 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_171
timestamp 1698175906
transform 1 0 10248 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_177
timestamp 1698175906
transform 1 0 10584 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_241
timestamp 1698175906
transform 1 0 14168 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_247
timestamp 1698175906
transform 1 0 14504 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_311
timestamp 1698175906
transform 1 0 18088 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_317
timestamp 1698175906
transform 1 0 18424 0 1 5488
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2
timestamp 1698175906
transform 1 0 784 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698175906
transform 1 0 4368 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_72
timestamp 1698175906
transform 1 0 4704 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698175906
transform 1 0 8288 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_142 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8624 0 -1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_189
timestamp 1698175906
transform 1 0 11256 0 -1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_205
timestamp 1698175906
transform 1 0 12152 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_209
timestamp 1698175906
transform 1 0 12376 0 -1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_212
timestamp 1698175906
transform 1 0 12544 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_276
timestamp 1698175906
transform 1 0 16128 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_282
timestamp 1698175906
transform 1 0 16464 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_346
timestamp 1698175906
transform 1 0 20048 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_348
timestamp 1698175906
transform 1 0 20160 0 -1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698175906
transform 1 0 784 0 1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698175906
transform 1 0 2576 0 1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_37
timestamp 1698175906
transform 1 0 2744 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698175906
transform 1 0 6328 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_107
timestamp 1698175906
transform 1 0 6664 0 1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_115
timestamp 1698175906
transform 1 0 7112 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_119
timestamp 1698175906
transform 1 0 7336 0 1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_149
timestamp 1698175906
transform 1 0 9016 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_153
timestamp 1698175906
transform 1 0 9240 0 1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_169
timestamp 1698175906
transform 1 0 10136 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_173
timestamp 1698175906
transform 1 0 10360 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_177
timestamp 1698175906
transform 1 0 10584 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_241
timestamp 1698175906
transform 1 0 14168 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_247
timestamp 1698175906
transform 1 0 14504 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_311
timestamp 1698175906
transform 1 0 18088 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_317
timestamp 1698175906
transform 1 0 18424 0 1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_2
timestamp 1698175906
transform 1 0 784 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_66
timestamp 1698175906
transform 1 0 4368 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_72
timestamp 1698175906
transform 1 0 4704 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_136
timestamp 1698175906
transform 1 0 8288 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_142
timestamp 1698175906
transform 1 0 8624 0 -1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_158
timestamp 1698175906
transform 1 0 9520 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_190
timestamp 1698175906
transform 1 0 11312 0 -1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_206
timestamp 1698175906
transform 1 0 12208 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_224
timestamp 1698175906
transform 1 0 13216 0 -1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_256
timestamp 1698175906
transform 1 0 15008 0 -1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_272
timestamp 1698175906
transform 1 0 15904 0 -1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_282
timestamp 1698175906
transform 1 0 16464 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_346
timestamp 1698175906
transform 1 0 20048 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_348
timestamp 1698175906
transform 1 0 20160 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698175906
transform 1 0 784 0 1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698175906
transform 1 0 2576 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_37
timestamp 1698175906
transform 1 0 2744 0 1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_101
timestamp 1698175906
transform 1 0 6328 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_107
timestamp 1698175906
transform 1 0 6664 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_115
timestamp 1698175906
transform 1 0 7112 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_119
timestamp 1698175906
transform 1 0 7336 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_150
timestamp 1698175906
transform 1 0 9072 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_154
timestamp 1698175906
transform 1 0 9296 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_162
timestamp 1698175906
transform 1 0 9744 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_174
timestamp 1698175906
transform 1 0 10416 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_177
timestamp 1698175906
transform 1 0 10584 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_184
timestamp 1698175906
transform 1 0 10976 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_192
timestamp 1698175906
transform 1 0 11424 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_196
timestamp 1698175906
transform 1 0 11648 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_198
timestamp 1698175906
transform 1 0 11760 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_228
timestamp 1698175906
transform 1 0 13440 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_232
timestamp 1698175906
transform 1 0 13664 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_240
timestamp 1698175906
transform 1 0 14112 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_244
timestamp 1698175906
transform 1 0 14336 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_247
timestamp 1698175906
transform 1 0 14504 0 1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_311
timestamp 1698175906
transform 1 0 18088 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_317
timestamp 1698175906
transform 1 0 18424 0 1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_2
timestamp 1698175906
transform 1 0 784 0 -1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_66
timestamp 1698175906
transform 1 0 4368 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_72
timestamp 1698175906
transform 1 0 4704 0 -1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_104
timestamp 1698175906
transform 1 0 6496 0 -1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_120
timestamp 1698175906
transform 1 0 7392 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_128
timestamp 1698175906
transform 1 0 7840 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_132
timestamp 1698175906
transform 1 0 8064 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_134
timestamp 1698175906
transform 1 0 8176 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_142
timestamp 1698175906
transform 1 0 8624 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_160
timestamp 1698175906
transform 1 0 9632 0 -1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_176
timestamp 1698175906
transform 1 0 10528 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_180
timestamp 1698175906
transform 1 0 10752 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_187
timestamp 1698175906
transform 1 0 11144 0 -1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_203
timestamp 1698175906
transform 1 0 12040 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_207
timestamp 1698175906
transform 1 0 12264 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_209
timestamp 1698175906
transform 1 0 12376 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_241
timestamp 1698175906
transform 1 0 14168 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_245
timestamp 1698175906
transform 1 0 14392 0 -1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_277
timestamp 1698175906
transform 1 0 16184 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_279
timestamp 1698175906
transform 1 0 16296 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_282
timestamp 1698175906
transform 1 0 16464 0 -1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_346
timestamp 1698175906
transform 1 0 20048 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_348
timestamp 1698175906
transform 1 0 20160 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_2
timestamp 1698175906
transform 1 0 784 0 1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698175906
transform 1 0 2576 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_37
timestamp 1698175906
transform 1 0 2744 0 1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_101
timestamp 1698175906
transform 1 0 6328 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_107
timestamp 1698175906
transform 1 0 6664 0 1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_139
timestamp 1698175906
transform 1 0 8456 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_143
timestamp 1698175906
transform 1 0 8680 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_150
timestamp 1698175906
transform 1 0 9072 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_158
timestamp 1698175906
transform 1 0 9520 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_160
timestamp 1698175906
transform 1 0 9632 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_172
timestamp 1698175906
transform 1 0 10304 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_174
timestamp 1698175906
transform 1 0 10416 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_177
timestamp 1698175906
transform 1 0 10584 0 1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_209
timestamp 1698175906
transform 1 0 12376 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_213
timestamp 1698175906
transform 1 0 12600 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_223
timestamp 1698175906
transform 1 0 13160 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_231
timestamp 1698175906
transform 1 0 13608 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_235
timestamp 1698175906
transform 1 0 13832 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_242
timestamp 1698175906
transform 1 0 14224 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_244
timestamp 1698175906
transform 1 0 14336 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_247
timestamp 1698175906
transform 1 0 14504 0 1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_311
timestamp 1698175906
transform 1 0 18088 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_317
timestamp 1698175906
transform 1 0 18424 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_321
timestamp 1698175906
transform 1 0 18648 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_2
timestamp 1698175906
transform 1 0 784 0 -1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_66
timestamp 1698175906
transform 1 0 4368 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_72
timestamp 1698175906
transform 1 0 4704 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_80
timestamp 1698175906
transform 1 0 5152 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_84
timestamp 1698175906
transform 1 0 5376 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_86
timestamp 1698175906
transform 1 0 5488 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_116
timestamp 1698175906
transform 1 0 7168 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_120
timestamp 1698175906
transform 1 0 7392 0 -1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_136
timestamp 1698175906
transform 1 0 8288 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_142
timestamp 1698175906
transform 1 0 8624 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_146
timestamp 1698175906
transform 1 0 8848 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_148
timestamp 1698175906
transform 1 0 8960 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_159
timestamp 1698175906
transform 1 0 9576 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_161
timestamp 1698175906
transform 1 0 9688 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_168
timestamp 1698175906
transform 1 0 10080 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_176
timestamp 1698175906
transform 1 0 10528 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_190
timestamp 1698175906
transform 1 0 11312 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_206
timestamp 1698175906
transform 1 0 12208 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_212
timestamp 1698175906
transform 1 0 12544 0 -1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_228
timestamp 1698175906
transform 1 0 13440 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_261
timestamp 1698175906
transform 1 0 15288 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_265
timestamp 1698175906
transform 1 0 15512 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_273
timestamp 1698175906
transform 1 0 15960 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_277
timestamp 1698175906
transform 1 0 16184 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_279
timestamp 1698175906
transform 1 0 16296 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_282
timestamp 1698175906
transform 1 0 16464 0 -1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_346
timestamp 1698175906
transform 1 0 20048 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_348
timestamp 1698175906
transform 1 0 20160 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_28
timestamp 1698175906
transform 1 0 2240 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_32
timestamp 1698175906
transform 1 0 2464 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698175906
transform 1 0 2576 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_37
timestamp 1698175906
transform 1 0 2744 0 1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_101
timestamp 1698175906
transform 1 0 6328 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_107
timestamp 1698175906
transform 1 0 6664 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_142
timestamp 1698175906
transform 1 0 8624 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_146
timestamp 1698175906
transform 1 0 8848 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_170
timestamp 1698175906
transform 1 0 10192 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_174
timestamp 1698175906
transform 1 0 10416 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_227
timestamp 1698175906
transform 1 0 13384 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_231
timestamp 1698175906
transform 1 0 13608 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_234
timestamp 1698175906
transform 1 0 13776 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_242
timestamp 1698175906
transform 1 0 14224 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_244
timestamp 1698175906
transform 1 0 14336 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_252
timestamp 1698175906
transform 1 0 14784 0 1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_284
timestamp 1698175906
transform 1 0 16576 0 1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_300
timestamp 1698175906
transform 1 0 17472 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_308
timestamp 1698175906
transform 1 0 17920 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_312
timestamp 1698175906
transform 1 0 18144 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_314
timestamp 1698175906
transform 1 0 18256 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_317
timestamp 1698175906
transform 1 0 18424 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_321
timestamp 1698175906
transform 1 0 18648 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_2
timestamp 1698175906
transform 1 0 784 0 -1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_66
timestamp 1698175906
transform 1 0 4368 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_72
timestamp 1698175906
transform 1 0 4704 0 -1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_104
timestamp 1698175906
transform 1 0 6496 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_108
timestamp 1698175906
transform 1 0 6720 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_117
timestamp 1698175906
transform 1 0 7224 0 -1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_133
timestamp 1698175906
transform 1 0 8120 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_142
timestamp 1698175906
transform 1 0 8624 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_166
timestamp 1698175906
transform 1 0 9968 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_170
timestamp 1698175906
transform 1 0 10192 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_192
timestamp 1698175906
transform 1 0 11424 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_206
timestamp 1698175906
transform 1 0 12208 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_241
timestamp 1698175906
transform 1 0 14168 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_245
timestamp 1698175906
transform 1 0 14392 0 -1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_277
timestamp 1698175906
transform 1 0 16184 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_279
timestamp 1698175906
transform 1 0 16296 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_282
timestamp 1698175906
transform 1 0 16464 0 -1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_346
timestamp 1698175906
transform 1 0 20048 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_348
timestamp 1698175906
transform 1 0 20160 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_2
timestamp 1698175906
transform 1 0 784 0 1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698175906
transform 1 0 2576 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_37
timestamp 1698175906
transform 1 0 2744 0 1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_101
timestamp 1698175906
transform 1 0 6328 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_136
timestamp 1698175906
transform 1 0 8288 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_160
timestamp 1698175906
transform 1 0 9632 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_193
timestamp 1698175906
transform 1 0 11480 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_262
timestamp 1698175906
transform 1 0 15344 0 1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_294
timestamp 1698175906
transform 1 0 17136 0 1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_310
timestamp 1698175906
transform 1 0 18032 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_314
timestamp 1698175906
transform 1 0 18256 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_317
timestamp 1698175906
transform 1 0 18424 0 1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_2
timestamp 1698175906
transform 1 0 784 0 -1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_66
timestamp 1698175906
transform 1 0 4368 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_72
timestamp 1698175906
transform 1 0 4704 0 -1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_88
timestamp 1698175906
transform 1 0 5600 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_96
timestamp 1698175906
transform 1 0 6048 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_100
timestamp 1698175906
transform 1 0 6272 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_103
timestamp 1698175906
transform 1 0 6440 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_112
timestamp 1698175906
transform 1 0 6944 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_118
timestamp 1698175906
transform 1 0 7280 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_120
timestamp 1698175906
transform 1 0 7392 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_126
timestamp 1698175906
transform 1 0 7728 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_192
timestamp 1698175906
transform 1 0 11424 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_200
timestamp 1698175906
transform 1 0 11872 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_262
timestamp 1698175906
transform 1 0 15344 0 -1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_278
timestamp 1698175906
transform 1 0 16240 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_282
timestamp 1698175906
transform 1 0 16464 0 -1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_314
timestamp 1698175906
transform 1 0 18256 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_322
timestamp 1698175906
transform 1 0 18704 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_28
timestamp 1698175906
transform 1 0 2240 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_32
timestamp 1698175906
transform 1 0 2464 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698175906
transform 1 0 2576 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_37
timestamp 1698175906
transform 1 0 2744 0 1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_69
timestamp 1698175906
transform 1 0 4536 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_73
timestamp 1698175906
transform 1 0 4760 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_75
timestamp 1698175906
transform 1 0 4872 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_112
timestamp 1698175906
transform 1 0 6944 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_118
timestamp 1698175906
transform 1 0 7280 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_126
timestamp 1698175906
transform 1 0 7728 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_134
timestamp 1698175906
transform 1 0 8176 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_136
timestamp 1698175906
transform 1 0 8288 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_227
timestamp 1698175906
transform 1 0 13384 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_235
timestamp 1698175906
transform 1 0 13832 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_237
timestamp 1698175906
transform 1 0 13944 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_276
timestamp 1698175906
transform 1 0 16128 0 1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_308
timestamp 1698175906
transform 1 0 17920 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_312
timestamp 1698175906
transform 1 0 18144 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_314
timestamp 1698175906
transform 1 0 18256 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_317
timestamp 1698175906
transform 1 0 18424 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_321
timestamp 1698175906
transform 1 0 18648 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_2
timestamp 1698175906
transform 1 0 784 0 -1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_66
timestamp 1698175906
transform 1 0 4368 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_72
timestamp 1698175906
transform 1 0 4704 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_80
timestamp 1698175906
transform 1 0 5152 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_84
timestamp 1698175906
transform 1 0 5376 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_86
timestamp 1698175906
transform 1 0 5488 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_124
timestamp 1698175906
transform 1 0 7616 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_130
timestamp 1698175906
transform 1 0 7952 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_134
timestamp 1698175906
transform 1 0 8176 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_138
timestamp 1698175906
transform 1 0 8400 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_142
timestamp 1698175906
transform 1 0 8624 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_166
timestamp 1698175906
transform 1 0 9968 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_170
timestamp 1698175906
transform 1 0 10192 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_172
timestamp 1698175906
transform 1 0 10304 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_181
timestamp 1698175906
transform 1 0 10808 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_198
timestamp 1698175906
transform 1 0 11760 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_212
timestamp 1698175906
transform 1 0 12544 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_220
timestamp 1698175906
transform 1 0 12992 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_224
timestamp 1698175906
transform 1 0 13216 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_226
timestamp 1698175906
transform 1 0 13328 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_232
timestamp 1698175906
transform 1 0 13664 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_236
timestamp 1698175906
transform 1 0 13888 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_266
timestamp 1698175906
transform 1 0 15568 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_270
timestamp 1698175906
transform 1 0 15792 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_278
timestamp 1698175906
transform 1 0 16240 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_282
timestamp 1698175906
transform 1 0 16464 0 -1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_346
timestamp 1698175906
transform 1 0 20048 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_348
timestamp 1698175906
transform 1 0 20160 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_28
timestamp 1698175906
transform 1 0 2240 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_32
timestamp 1698175906
transform 1 0 2464 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698175906
transform 1 0 2576 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_37
timestamp 1698175906
transform 1 0 2744 0 1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_101
timestamp 1698175906
transform 1 0 6328 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_111
timestamp 1698175906
transform 1 0 6888 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_122
timestamp 1698175906
transform 1 0 7504 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_124
timestamp 1698175906
transform 1 0 7616 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_133
timestamp 1698175906
transform 1 0 8120 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_152
timestamp 1698175906
transform 1 0 9184 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_154
timestamp 1698175906
transform 1 0 9296 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_168
timestamp 1698175906
transform 1 0 10080 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_172
timestamp 1698175906
transform 1 0 10304 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_174
timestamp 1698175906
transform 1 0 10416 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_177
timestamp 1698175906
transform 1 0 10584 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_203
timestamp 1698175906
transform 1 0 12040 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_239
timestamp 1698175906
transform 1 0 14056 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_243
timestamp 1698175906
transform 1 0 14280 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_247
timestamp 1698175906
transform 1 0 14504 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_249
timestamp 1698175906
transform 1 0 14616 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_256
timestamp 1698175906
transform 1 0 15008 0 1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_288
timestamp 1698175906
transform 1 0 16800 0 1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_304
timestamp 1698175906
transform 1 0 17696 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_312
timestamp 1698175906
transform 1 0 18144 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_314
timestamp 1698175906
transform 1 0 18256 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_317
timestamp 1698175906
transform 1 0 18424 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_321
timestamp 1698175906
transform 1 0 18648 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_28
timestamp 1698175906
transform 1 0 2240 0 -1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_60
timestamp 1698175906
transform 1 0 4032 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_68
timestamp 1698175906
transform 1 0 4480 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_72
timestamp 1698175906
transform 1 0 4704 0 -1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_88
timestamp 1698175906
transform 1 0 5600 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_92
timestamp 1698175906
transform 1 0 5824 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_132
timestamp 1698175906
transform 1 0 8064 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_136
timestamp 1698175906
transform 1 0 8288 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_142
timestamp 1698175906
transform 1 0 8624 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_146
timestamp 1698175906
transform 1 0 8848 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_148
timestamp 1698175906
transform 1 0 8960 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_154
timestamp 1698175906
transform 1 0 9296 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_164
timestamp 1698175906
transform 1 0 9856 0 -1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_196
timestamp 1698175906
transform 1 0 11648 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_204
timestamp 1698175906
transform 1 0 12096 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_208
timestamp 1698175906
transform 1 0 12320 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_270
timestamp 1698175906
transform 1 0 15792 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_274
timestamp 1698175906
transform 1 0 16016 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_278
timestamp 1698175906
transform 1 0 16240 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_282
timestamp 1698175906
transform 1 0 16464 0 -1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_314
timestamp 1698175906
transform 1 0 18256 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_322
timestamp 1698175906
transform 1 0 18704 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_28
timestamp 1698175906
transform 1 0 2240 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_32
timestamp 1698175906
transform 1 0 2464 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698175906
transform 1 0 2576 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_37
timestamp 1698175906
transform 1 0 2744 0 1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_101
timestamp 1698175906
transform 1 0 6328 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_107
timestamp 1698175906
transform 1 0 6664 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_115
timestamp 1698175906
transform 1 0 7112 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_119
timestamp 1698175906
transform 1 0 7336 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_126
timestamp 1698175906
transform 1 0 7728 0 1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_142
timestamp 1698175906
transform 1 0 8624 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_156
timestamp 1698175906
transform 1 0 9408 0 1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_172
timestamp 1698175906
transform 1 0 10304 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_174
timestamp 1698175906
transform 1 0 10416 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_187
timestamp 1698175906
transform 1 0 11144 0 1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_203
timestamp 1698175906
transform 1 0 12040 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_211
timestamp 1698175906
transform 1 0 12488 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_226
timestamp 1698175906
transform 1 0 13328 0 1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_242
timestamp 1698175906
transform 1 0 14224 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_244
timestamp 1698175906
transform 1 0 14336 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_247
timestamp 1698175906
transform 1 0 14504 0 1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_311
timestamp 1698175906
transform 1 0 18088 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_317
timestamp 1698175906
transform 1 0 18424 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_321
timestamp 1698175906
transform 1 0 18648 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_2
timestamp 1698175906
transform 1 0 784 0 -1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_66
timestamp 1698175906
transform 1 0 4368 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_72
timestamp 1698175906
transform 1 0 4704 0 -1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_136
timestamp 1698175906
transform 1 0 8288 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_142
timestamp 1698175906
transform 1 0 8624 0 -1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_158
timestamp 1698175906
transform 1 0 9520 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_188
timestamp 1698175906
transform 1 0 11200 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_192
timestamp 1698175906
transform 1 0 11424 0 -1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_208
timestamp 1698175906
transform 1 0 12320 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_212
timestamp 1698175906
transform 1 0 12544 0 -1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_276
timestamp 1698175906
transform 1 0 16128 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_282
timestamp 1698175906
transform 1 0 16464 0 -1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_346
timestamp 1698175906
transform 1 0 20048 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_348
timestamp 1698175906
transform 1 0 20160 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_2
timestamp 1698175906
transform 1 0 784 0 1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698175906
transform 1 0 2576 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_37
timestamp 1698175906
transform 1 0 2744 0 1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_101
timestamp 1698175906
transform 1 0 6328 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_107
timestamp 1698175906
transform 1 0 6664 0 1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_123
timestamp 1698175906
transform 1 0 7560 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_131
timestamp 1698175906
transform 1 0 8008 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_154
timestamp 1698175906
transform 1 0 9296 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_162
timestamp 1698175906
transform 1 0 9744 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_164
timestamp 1698175906
transform 1 0 9856 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_173
timestamp 1698175906
transform 1 0 10360 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_198
timestamp 1698175906
transform 1 0 11760 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_206
timestamp 1698175906
transform 1 0 12208 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_219
timestamp 1698175906
transform 1 0 12936 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_235
timestamp 1698175906
transform 1 0 13832 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_243
timestamp 1698175906
transform 1 0 14280 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_247
timestamp 1698175906
transform 1 0 14504 0 1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_311
timestamp 1698175906
transform 1 0 18088 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_317
timestamp 1698175906
transform 1 0 18424 0 1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_2
timestamp 1698175906
transform 1 0 784 0 -1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_66
timestamp 1698175906
transform 1 0 4368 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_72
timestamp 1698175906
transform 1 0 4704 0 -1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_104
timestamp 1698175906
transform 1 0 6496 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_108
timestamp 1698175906
transform 1 0 6720 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_110
timestamp 1698175906
transform 1 0 6832 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_151
timestamp 1698175906
transform 1 0 9128 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_163
timestamp 1698175906
transform 1 0 9800 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_176
timestamp 1698175906
transform 1 0 10528 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_180
timestamp 1698175906
transform 1 0 10752 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_182
timestamp 1698175906
transform 1 0 10864 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_189
timestamp 1698175906
transform 1 0 11256 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_193
timestamp 1698175906
transform 1 0 11480 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_199
timestamp 1698175906
transform 1 0 11816 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_241
timestamp 1698175906
transform 1 0 14168 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_245
timestamp 1698175906
transform 1 0 14392 0 -1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_277
timestamp 1698175906
transform 1 0 16184 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_279
timestamp 1698175906
transform 1 0 16296 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_282
timestamp 1698175906
transform 1 0 16464 0 -1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_314
timestamp 1698175906
transform 1 0 18256 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_322
timestamp 1698175906
transform 1 0 18704 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_2
timestamp 1698175906
transform 1 0 784 0 1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698175906
transform 1 0 2576 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_37
timestamp 1698175906
transform 1 0 2744 0 1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_101
timestamp 1698175906
transform 1 0 6328 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_107
timestamp 1698175906
transform 1 0 6664 0 1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_115
timestamp 1698175906
transform 1 0 7112 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_153
timestamp 1698175906
transform 1 0 9240 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_163
timestamp 1698175906
transform 1 0 9800 0 1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_171
timestamp 1698175906
transform 1 0 10248 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_177
timestamp 1698175906
transform 1 0 10584 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_237
timestamp 1698175906
transform 1 0 13944 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_241
timestamp 1698175906
transform 1 0 14168 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_247
timestamp 1698175906
transform 1 0 14504 0 1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_311
timestamp 1698175906
transform 1 0 18088 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_317
timestamp 1698175906
transform 1 0 18424 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_321
timestamp 1698175906
transform 1 0 18648 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_2
timestamp 1698175906
transform 1 0 784 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_66
timestamp 1698175906
transform 1 0 4368 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_72
timestamp 1698175906
transform 1 0 4704 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_136
timestamp 1698175906
transform 1 0 8288 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_148
timestamp 1698175906
transform 1 0 8960 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_179
timestamp 1698175906
transform 1 0 10696 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_183
timestamp 1698175906
transform 1 0 10920 0 -1 14112
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_199
timestamp 1698175906
transform 1 0 11816 0 -1 14112
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_207
timestamp 1698175906
transform 1 0 12264 0 -1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_212
timestamp 1698175906
transform 1 0 12544 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_276
timestamp 1698175906
transform 1 0 16128 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_282
timestamp 1698175906
transform 1 0 16464 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_346
timestamp 1698175906
transform 1 0 20048 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_348
timestamp 1698175906
transform 1 0 20160 0 -1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_2
timestamp 1698175906
transform 1 0 784 0 1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698175906
transform 1 0 2576 0 1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_37
timestamp 1698175906
transform 1 0 2744 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_101
timestamp 1698175906
transform 1 0 6328 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_107
timestamp 1698175906
transform 1 0 6664 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_171
timestamp 1698175906
transform 1 0 10248 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_177
timestamp 1698175906
transform 1 0 10584 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_241
timestamp 1698175906
transform 1 0 14168 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_247
timestamp 1698175906
transform 1 0 14504 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_311
timestamp 1698175906
transform 1 0 18088 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_317
timestamp 1698175906
transform 1 0 18424 0 1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_2
timestamp 1698175906
transform 1 0 784 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_66
timestamp 1698175906
transform 1 0 4368 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_72
timestamp 1698175906
transform 1 0 4704 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_136
timestamp 1698175906
transform 1 0 8288 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_142
timestamp 1698175906
transform 1 0 8624 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_206
timestamp 1698175906
transform 1 0 12208 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_212
timestamp 1698175906
transform 1 0 12544 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_276
timestamp 1698175906
transform 1 0 16128 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_282
timestamp 1698175906
transform 1 0 16464 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_346
timestamp 1698175906
transform 1 0 20048 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_348
timestamp 1698175906
transform 1 0 20160 0 -1 14896
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698175906
transform 1 0 784 0 1 14896
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698175906
transform 1 0 2576 0 1 14896
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_37
timestamp 1698175906
transform 1 0 2744 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_101
timestamp 1698175906
transform 1 0 6328 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_107
timestamp 1698175906
transform 1 0 6664 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_171
timestamp 1698175906
transform 1 0 10248 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_177
timestamp 1698175906
transform 1 0 10584 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_241
timestamp 1698175906
transform 1 0 14168 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_247
timestamp 1698175906
transform 1 0 14504 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_311
timestamp 1698175906
transform 1 0 18088 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_317
timestamp 1698175906
transform 1 0 18424 0 1 14896
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2
timestamp 1698175906
transform 1 0 784 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_66
timestamp 1698175906
transform 1 0 4368 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_72
timestamp 1698175906
transform 1 0 4704 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_136
timestamp 1698175906
transform 1 0 8288 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_142
timestamp 1698175906
transform 1 0 8624 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_206
timestamp 1698175906
transform 1 0 12208 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_212
timestamp 1698175906
transform 1 0 12544 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_276
timestamp 1698175906
transform 1 0 16128 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_282
timestamp 1698175906
transform 1 0 16464 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_346
timestamp 1698175906
transform 1 0 20048 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_348
timestamp 1698175906
transform 1 0 20160 0 -1 15680
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_2
timestamp 1698175906
transform 1 0 784 0 1 15680
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698175906
transform 1 0 2576 0 1 15680
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_37
timestamp 1698175906
transform 1 0 2744 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_101
timestamp 1698175906
transform 1 0 6328 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_107
timestamp 1698175906
transform 1 0 6664 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_171
timestamp 1698175906
transform 1 0 10248 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_177
timestamp 1698175906
transform 1 0 10584 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_241
timestamp 1698175906
transform 1 0 14168 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_247
timestamp 1698175906
transform 1 0 14504 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_311
timestamp 1698175906
transform 1 0 18088 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_317
timestamp 1698175906
transform 1 0 18424 0 1 15680
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2
timestamp 1698175906
transform 1 0 784 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_66
timestamp 1698175906
transform 1 0 4368 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_72
timestamp 1698175906
transform 1 0 4704 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_136
timestamp 1698175906
transform 1 0 8288 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_142
timestamp 1698175906
transform 1 0 8624 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_206
timestamp 1698175906
transform 1 0 12208 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_212
timestamp 1698175906
transform 1 0 12544 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_276
timestamp 1698175906
transform 1 0 16128 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_282
timestamp 1698175906
transform 1 0 16464 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_346
timestamp 1698175906
transform 1 0 20048 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_348
timestamp 1698175906
transform 1 0 20160 0 -1 16464
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698175906
transform 1 0 784 0 1 16464
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698175906
transform 1 0 2576 0 1 16464
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_37
timestamp 1698175906
transform 1 0 2744 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_101
timestamp 1698175906
transform 1 0 6328 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_107
timestamp 1698175906
transform 1 0 6664 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_171
timestamp 1698175906
transform 1 0 10248 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_177
timestamp 1698175906
transform 1 0 10584 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_241
timestamp 1698175906
transform 1 0 14168 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_247
timestamp 1698175906
transform 1 0 14504 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_311
timestamp 1698175906
transform 1 0 18088 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_317
timestamp 1698175906
transform 1 0 18424 0 1 16464
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_2
timestamp 1698175906
transform 1 0 784 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_66
timestamp 1698175906
transform 1 0 4368 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_72
timestamp 1698175906
transform 1 0 4704 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_136
timestamp 1698175906
transform 1 0 8288 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_142
timestamp 1698175906
transform 1 0 8624 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_206
timestamp 1698175906
transform 1 0 12208 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_212
timestamp 1698175906
transform 1 0 12544 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_276
timestamp 1698175906
transform 1 0 16128 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_282
timestamp 1698175906
transform 1 0 16464 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_346
timestamp 1698175906
transform 1 0 20048 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_348
timestamp 1698175906
transform 1 0 20160 0 -1 17248
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698175906
transform 1 0 784 0 1 17248
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698175906
transform 1 0 2576 0 1 17248
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_37
timestamp 1698175906
transform 1 0 2744 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_101
timestamp 1698175906
transform 1 0 6328 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_107
timestamp 1698175906
transform 1 0 6664 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_171
timestamp 1698175906
transform 1 0 10248 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_177
timestamp 1698175906
transform 1 0 10584 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_241
timestamp 1698175906
transform 1 0 14168 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_247
timestamp 1698175906
transform 1 0 14504 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_311
timestamp 1698175906
transform 1 0 18088 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_317
timestamp 1698175906
transform 1 0 18424 0 1 17248
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2
timestamp 1698175906
transform 1 0 784 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1698175906
transform 1 0 4368 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_72
timestamp 1698175906
transform 1 0 4704 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_136
timestamp 1698175906
transform 1 0 8288 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_142
timestamp 1698175906
transform 1 0 8624 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_206
timestamp 1698175906
transform 1 0 12208 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_212
timestamp 1698175906
transform 1 0 12544 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_276
timestamp 1698175906
transform 1 0 16128 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_282
timestamp 1698175906
transform 1 0 16464 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_346
timestamp 1698175906
transform 1 0 20048 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_348
timestamp 1698175906
transform 1 0 20160 0 -1 18032
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_2
timestamp 1698175906
transform 1 0 784 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698175906
transform 1 0 2576 0 1 18032
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_37
timestamp 1698175906
transform 1 0 2744 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_101
timestamp 1698175906
transform 1 0 6328 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_107
timestamp 1698175906
transform 1 0 6664 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_165
timestamp 1698175906
transform 1 0 9912 0 1 18032
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_173
timestamp 1698175906
transform 1 0 10360 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_177
timestamp 1698175906
transform 1 0 10584 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_241
timestamp 1698175906
transform 1 0 14168 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_247
timestamp 1698175906
transform 1 0 14504 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_311
timestamp 1698175906
transform 1 0 18088 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_317
timestamp 1698175906
transform 1 0 18424 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_2
timestamp 1698175906
transform 1 0 784 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_66
timestamp 1698175906
transform 1 0 4368 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_72
timestamp 1698175906
transform 1 0 4704 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_136
timestamp 1698175906
transform 1 0 8288 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_142
timestamp 1698175906
transform 1 0 8624 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_144
timestamp 1698175906
transform 1 0 8736 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_171
timestamp 1698175906
transform 1 0 10248 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_201
timestamp 1698175906
transform 1 0 11928 0 -1 18816
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_209
timestamp 1698175906
transform 1 0 12376 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_212
timestamp 1698175906
transform 1 0 12544 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_276
timestamp 1698175906
transform 1 0 16128 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_282
timestamp 1698175906
transform 1 0 16464 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_346
timestamp 1698175906
transform 1 0 20048 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_348
timestamp 1698175906
transform 1 0 20160 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_2
timestamp 1698175906
transform 1 0 784 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_36
timestamp 1698175906
transform 1 0 2688 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_70
timestamp 1698175906
transform 1 0 4592 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_104
timestamp 1698175906
transform 1 0 6496 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_108
timestamp 1698175906
transform 1 0 6720 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_138
timestamp 1698175906
transform 1 0 8400 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_142
timestamp 1698175906
transform 1 0 8624 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_172
timestamp 1698175906
transform 1 0 10304 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_176
timestamp 1698175906
transform 1 0 10528 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_232
timestamp 1698175906
transform 1 0 13664 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_236
timestamp 1698175906
transform 1 0 13888 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_240
timestamp 1698175906
transform 1 0 14112 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_274
timestamp 1698175906
transform 1 0 16016 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_308
timestamp 1698175906
transform 1 0 17920 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_342
timestamp 1698175906
transform 1 0 19824 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_346
timestamp 1698175906
transform 1 0 20048 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_348
timestamp 1698175906
transform 1 0 20160 0 1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 2240 0 1 11760
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output2
timestamp 1698175906
transform 1 0 12208 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output3
timestamp 1698175906
transform 1 0 10640 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output4
timestamp 1698175906
transform 1 0 18760 0 1 7840
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output5
timestamp 1698175906
transform -1 0 2240 0 -1 11760
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output6
timestamp 1698175906
transform 1 0 18760 0 -1 11760
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output7
timestamp 1698175906
transform 1 0 8792 0 -1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output8
timestamp 1698175906
transform -1 0 2240 0 1 10976
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output9
timestamp 1698175906
transform 1 0 18760 0 1 10976
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output10
timestamp 1698175906
transform -1 0 8288 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output11
timestamp 1698175906
transform 1 0 10640 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output12
timestamp 1698175906
transform 1 0 8456 0 1 18032
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output13
timestamp 1698175906
transform 1 0 18760 0 -1 13328
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output14
timestamp 1698175906
transform 1 0 18760 0 1 13328
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output15
timestamp 1698175906
transform 1 0 8792 0 -1 2352
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output16
timestamp 1698175906
transform -1 0 2240 0 1 8624
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output17
timestamp 1698175906
transform -1 0 14000 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output18
timestamp 1698175906
transform 1 0 18760 0 1 10192
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output19
timestamp 1698175906
transform 1 0 8736 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output20
timestamp 1698175906
transform 1 0 8736 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output21
timestamp 1698175906
transform 1 0 10808 0 -1 2352
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output22
timestamp 1698175906
transform 1 0 10472 0 -1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output23
timestamp 1698175906
transform 1 0 18760 0 1 11760
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output24
timestamp 1698175906
transform 1 0 18760 0 1 8624
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output25
timestamp 1698175906
transform -1 0 2240 0 1 10192
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output26
timestamp 1698175906
transform 1 0 18760 0 -1 10192
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_45 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 672 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698175906
transform -1 0 20328 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_46
timestamp 1698175906
transform 1 0 672 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698175906
transform -1 0 20328 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_47
timestamp 1698175906
transform 1 0 672 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698175906
transform -1 0 20328 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_48
timestamp 1698175906
transform 1 0 672 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698175906
transform -1 0 20328 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_49
timestamp 1698175906
transform 1 0 672 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698175906
transform -1 0 20328 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_50
timestamp 1698175906
transform 1 0 672 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698175906
transform -1 0 20328 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_51
timestamp 1698175906
transform 1 0 672 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698175906
transform -1 0 20328 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_52
timestamp 1698175906
transform 1 0 672 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698175906
transform -1 0 20328 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_53
timestamp 1698175906
transform 1 0 672 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698175906
transform -1 0 20328 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_54
timestamp 1698175906
transform 1 0 672 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698175906
transform -1 0 20328 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_55
timestamp 1698175906
transform 1 0 672 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698175906
transform -1 0 20328 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_56
timestamp 1698175906
transform 1 0 672 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698175906
transform -1 0 20328 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_57
timestamp 1698175906
transform 1 0 672 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698175906
transform -1 0 20328 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_58
timestamp 1698175906
transform 1 0 672 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698175906
transform -1 0 20328 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_59
timestamp 1698175906
transform 1 0 672 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698175906
transform -1 0 20328 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_60
timestamp 1698175906
transform 1 0 672 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698175906
transform -1 0 20328 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_61
timestamp 1698175906
transform 1 0 672 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698175906
transform -1 0 20328 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_62
timestamp 1698175906
transform 1 0 672 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698175906
transform -1 0 20328 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_63
timestamp 1698175906
transform 1 0 672 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698175906
transform -1 0 20328 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_64
timestamp 1698175906
transform 1 0 672 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698175906
transform -1 0 20328 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_65
timestamp 1698175906
transform 1 0 672 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698175906
transform -1 0 20328 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_66
timestamp 1698175906
transform 1 0 672 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698175906
transform -1 0 20328 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_67
timestamp 1698175906
transform 1 0 672 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698175906
transform -1 0 20328 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_68
timestamp 1698175906
transform 1 0 672 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698175906
transform -1 0 20328 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_69
timestamp 1698175906
transform 1 0 672 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698175906
transform -1 0 20328 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_70
timestamp 1698175906
transform 1 0 672 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698175906
transform -1 0 20328 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_71
timestamp 1698175906
transform 1 0 672 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698175906
transform -1 0 20328 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_72
timestamp 1698175906
transform 1 0 672 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698175906
transform -1 0 20328 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_73
timestamp 1698175906
transform 1 0 672 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698175906
transform -1 0 20328 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_74
timestamp 1698175906
transform 1 0 672 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698175906
transform -1 0 20328 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_75
timestamp 1698175906
transform 1 0 672 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698175906
transform -1 0 20328 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_76
timestamp 1698175906
transform 1 0 672 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698175906
transform -1 0 20328 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_77
timestamp 1698175906
transform 1 0 672 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698175906
transform -1 0 20328 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_78
timestamp 1698175906
transform 1 0 672 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698175906
transform -1 0 20328 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_79
timestamp 1698175906
transform 1 0 672 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698175906
transform -1 0 20328 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_80
timestamp 1698175906
transform 1 0 672 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698175906
transform -1 0 20328 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_81
timestamp 1698175906
transform 1 0 672 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698175906
transform -1 0 20328 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_82
timestamp 1698175906
transform 1 0 672 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698175906
transform -1 0 20328 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_83
timestamp 1698175906
transform 1 0 672 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698175906
transform -1 0 20328 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_84
timestamp 1698175906
transform 1 0 672 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698175906
transform -1 0 20328 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_85
timestamp 1698175906
transform 1 0 672 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698175906
transform -1 0 20328 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_86
timestamp 1698175906
transform 1 0 672 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698175906
transform -1 0 20328 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_87
timestamp 1698175906
transform 1 0 672 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698175906
transform -1 0 20328 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_88
timestamp 1698175906
transform 1 0 672 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698175906
transform -1 0 20328 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_89
timestamp 1698175906
transform 1 0 672 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698175906
transform -1 0 20328 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_90 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 2576 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_91
timestamp 1698175906
transform 1 0 4480 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_92
timestamp 1698175906
transform 1 0 6384 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_93
timestamp 1698175906
transform 1 0 8288 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_94
timestamp 1698175906
transform 1 0 10192 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_95
timestamp 1698175906
transform 1 0 12096 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_96
timestamp 1698175906
transform 1 0 14000 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_97
timestamp 1698175906
transform 1 0 15904 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_98
timestamp 1698175906
transform 1 0 17808 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_99
timestamp 1698175906
transform 1 0 19712 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_100
timestamp 1698175906
transform 1 0 4592 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_101
timestamp 1698175906
transform 1 0 8512 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_102
timestamp 1698175906
transform 1 0 12432 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_103
timestamp 1698175906
transform 1 0 16352 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_104
timestamp 1698175906
transform 1 0 2632 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_105
timestamp 1698175906
transform 1 0 6552 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_106
timestamp 1698175906
transform 1 0 10472 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_107
timestamp 1698175906
transform 1 0 14392 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_108
timestamp 1698175906
transform 1 0 18312 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_109
timestamp 1698175906
transform 1 0 4592 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_110
timestamp 1698175906
transform 1 0 8512 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_111
timestamp 1698175906
transform 1 0 12432 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_112
timestamp 1698175906
transform 1 0 16352 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_113
timestamp 1698175906
transform 1 0 2632 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_114
timestamp 1698175906
transform 1 0 6552 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_115
timestamp 1698175906
transform 1 0 10472 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_116
timestamp 1698175906
transform 1 0 14392 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_117
timestamp 1698175906
transform 1 0 18312 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_118
timestamp 1698175906
transform 1 0 4592 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_119
timestamp 1698175906
transform 1 0 8512 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_120
timestamp 1698175906
transform 1 0 12432 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_121
timestamp 1698175906
transform 1 0 16352 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_122
timestamp 1698175906
transform 1 0 2632 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_123
timestamp 1698175906
transform 1 0 6552 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_124
timestamp 1698175906
transform 1 0 10472 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_125
timestamp 1698175906
transform 1 0 14392 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_126
timestamp 1698175906
transform 1 0 18312 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_127
timestamp 1698175906
transform 1 0 4592 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_128
timestamp 1698175906
transform 1 0 8512 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_129
timestamp 1698175906
transform 1 0 12432 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_130
timestamp 1698175906
transform 1 0 16352 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_131
timestamp 1698175906
transform 1 0 2632 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_132
timestamp 1698175906
transform 1 0 6552 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_133
timestamp 1698175906
transform 1 0 10472 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_134
timestamp 1698175906
transform 1 0 14392 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_135
timestamp 1698175906
transform 1 0 18312 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_136
timestamp 1698175906
transform 1 0 4592 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_137
timestamp 1698175906
transform 1 0 8512 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_138
timestamp 1698175906
transform 1 0 12432 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_139
timestamp 1698175906
transform 1 0 16352 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_140
timestamp 1698175906
transform 1 0 2632 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_141
timestamp 1698175906
transform 1 0 6552 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_142
timestamp 1698175906
transform 1 0 10472 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_143
timestamp 1698175906
transform 1 0 14392 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_144
timestamp 1698175906
transform 1 0 18312 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_145
timestamp 1698175906
transform 1 0 4592 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_146
timestamp 1698175906
transform 1 0 8512 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_147
timestamp 1698175906
transform 1 0 12432 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_148
timestamp 1698175906
transform 1 0 16352 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_149
timestamp 1698175906
transform 1 0 2632 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_150
timestamp 1698175906
transform 1 0 6552 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_151
timestamp 1698175906
transform 1 0 10472 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_152
timestamp 1698175906
transform 1 0 14392 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_153
timestamp 1698175906
transform 1 0 18312 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_154
timestamp 1698175906
transform 1 0 4592 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_155
timestamp 1698175906
transform 1 0 8512 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_156
timestamp 1698175906
transform 1 0 12432 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_157
timestamp 1698175906
transform 1 0 16352 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_158
timestamp 1698175906
transform 1 0 2632 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_159
timestamp 1698175906
transform 1 0 6552 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_160
timestamp 1698175906
transform 1 0 10472 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_161
timestamp 1698175906
transform 1 0 14392 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_162
timestamp 1698175906
transform 1 0 18312 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_163
timestamp 1698175906
transform 1 0 4592 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_164
timestamp 1698175906
transform 1 0 8512 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_165
timestamp 1698175906
transform 1 0 12432 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_166
timestamp 1698175906
transform 1 0 16352 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_167
timestamp 1698175906
transform 1 0 2632 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_168
timestamp 1698175906
transform 1 0 6552 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_169
timestamp 1698175906
transform 1 0 10472 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_170
timestamp 1698175906
transform 1 0 14392 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_171
timestamp 1698175906
transform 1 0 18312 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_172
timestamp 1698175906
transform 1 0 4592 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_173
timestamp 1698175906
transform 1 0 8512 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_174
timestamp 1698175906
transform 1 0 12432 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_175
timestamp 1698175906
transform 1 0 16352 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_176
timestamp 1698175906
transform 1 0 2632 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_177
timestamp 1698175906
transform 1 0 6552 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_178
timestamp 1698175906
transform 1 0 10472 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_179
timestamp 1698175906
transform 1 0 14392 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_180
timestamp 1698175906
transform 1 0 18312 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_181
timestamp 1698175906
transform 1 0 4592 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_182
timestamp 1698175906
transform 1 0 8512 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_183
timestamp 1698175906
transform 1 0 12432 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_184
timestamp 1698175906
transform 1 0 16352 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_185
timestamp 1698175906
transform 1 0 2632 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_186
timestamp 1698175906
transform 1 0 6552 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_187
timestamp 1698175906
transform 1 0 10472 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_188
timestamp 1698175906
transform 1 0 14392 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_189
timestamp 1698175906
transform 1 0 18312 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_190
timestamp 1698175906
transform 1 0 4592 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_191
timestamp 1698175906
transform 1 0 8512 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_192
timestamp 1698175906
transform 1 0 12432 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_193
timestamp 1698175906
transform 1 0 16352 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_194
timestamp 1698175906
transform 1 0 2632 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_195
timestamp 1698175906
transform 1 0 6552 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_196
timestamp 1698175906
transform 1 0 10472 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_197
timestamp 1698175906
transform 1 0 14392 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_198
timestamp 1698175906
transform 1 0 18312 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_199
timestamp 1698175906
transform 1 0 4592 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_200
timestamp 1698175906
transform 1 0 8512 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_201
timestamp 1698175906
transform 1 0 12432 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_202
timestamp 1698175906
transform 1 0 16352 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_203
timestamp 1698175906
transform 1 0 2632 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_204
timestamp 1698175906
transform 1 0 6552 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_205
timestamp 1698175906
transform 1 0 10472 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_206
timestamp 1698175906
transform 1 0 14392 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_207
timestamp 1698175906
transform 1 0 18312 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_208
timestamp 1698175906
transform 1 0 4592 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_209
timestamp 1698175906
transform 1 0 8512 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_210
timestamp 1698175906
transform 1 0 12432 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_211
timestamp 1698175906
transform 1 0 16352 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_212
timestamp 1698175906
transform 1 0 2632 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_213
timestamp 1698175906
transform 1 0 6552 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_214
timestamp 1698175906
transform 1 0 10472 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_215
timestamp 1698175906
transform 1 0 14392 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_216
timestamp 1698175906
transform 1 0 18312 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_217
timestamp 1698175906
transform 1 0 4592 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_218
timestamp 1698175906
transform 1 0 8512 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_219
timestamp 1698175906
transform 1 0 12432 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_220
timestamp 1698175906
transform 1 0 16352 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_221
timestamp 1698175906
transform 1 0 2632 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_222
timestamp 1698175906
transform 1 0 6552 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_223
timestamp 1698175906
transform 1 0 10472 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_224
timestamp 1698175906
transform 1 0 14392 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_225
timestamp 1698175906
transform 1 0 18312 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_226
timestamp 1698175906
transform 1 0 4592 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_227
timestamp 1698175906
transform 1 0 8512 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_228
timestamp 1698175906
transform 1 0 12432 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_229
timestamp 1698175906
transform 1 0 16352 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_230
timestamp 1698175906
transform 1 0 2632 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_231
timestamp 1698175906
transform 1 0 6552 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_232
timestamp 1698175906
transform 1 0 10472 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_233
timestamp 1698175906
transform 1 0 14392 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_234
timestamp 1698175906
transform 1 0 18312 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_235
timestamp 1698175906
transform 1 0 4592 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_236
timestamp 1698175906
transform 1 0 8512 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_237
timestamp 1698175906
transform 1 0 12432 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_238
timestamp 1698175906
transform 1 0 16352 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_239
timestamp 1698175906
transform 1 0 2632 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_240
timestamp 1698175906
transform 1 0 6552 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_241
timestamp 1698175906
transform 1 0 10472 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_242
timestamp 1698175906
transform 1 0 14392 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_243
timestamp 1698175906
transform 1 0 18312 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_244
timestamp 1698175906
transform 1 0 4592 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_245
timestamp 1698175906
transform 1 0 8512 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_246
timestamp 1698175906
transform 1 0 12432 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_247
timestamp 1698175906
transform 1 0 16352 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_248
timestamp 1698175906
transform 1 0 2632 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_249
timestamp 1698175906
transform 1 0 6552 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_250
timestamp 1698175906
transform 1 0 10472 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_251
timestamp 1698175906
transform 1 0 14392 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_252
timestamp 1698175906
transform 1 0 18312 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_253
timestamp 1698175906
transform 1 0 4592 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_254
timestamp 1698175906
transform 1 0 8512 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_255
timestamp 1698175906
transform 1 0 12432 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_256
timestamp 1698175906
transform 1 0 16352 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_257
timestamp 1698175906
transform 1 0 2632 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_258
timestamp 1698175906
transform 1 0 6552 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_259
timestamp 1698175906
transform 1 0 10472 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_260
timestamp 1698175906
transform 1 0 14392 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_261
timestamp 1698175906
transform 1 0 18312 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_262
timestamp 1698175906
transform 1 0 4592 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_263
timestamp 1698175906
transform 1 0 8512 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_264
timestamp 1698175906
transform 1 0 12432 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_265
timestamp 1698175906
transform 1 0 16352 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_266
timestamp 1698175906
transform 1 0 2632 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_267
timestamp 1698175906
transform 1 0 6552 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_268
timestamp 1698175906
transform 1 0 10472 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_269
timestamp 1698175906
transform 1 0 14392 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_270
timestamp 1698175906
transform 1 0 18312 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_271
timestamp 1698175906
transform 1 0 4592 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_272
timestamp 1698175906
transform 1 0 8512 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_273
timestamp 1698175906
transform 1 0 12432 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_274
timestamp 1698175906
transform 1 0 16352 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_275
timestamp 1698175906
transform 1 0 2632 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_276
timestamp 1698175906
transform 1 0 6552 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_277
timestamp 1698175906
transform 1 0 10472 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_278
timestamp 1698175906
transform 1 0 14392 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_279
timestamp 1698175906
transform 1 0 18312 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_280
timestamp 1698175906
transform 1 0 4592 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_281
timestamp 1698175906
transform 1 0 8512 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_282
timestamp 1698175906
transform 1 0 12432 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_283
timestamp 1698175906
transform 1 0 16352 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_284
timestamp 1698175906
transform 1 0 2632 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_285
timestamp 1698175906
transform 1 0 6552 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_286
timestamp 1698175906
transform 1 0 10472 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_287
timestamp 1698175906
transform 1 0 14392 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_288
timestamp 1698175906
transform 1 0 18312 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_289
timestamp 1698175906
transform 1 0 4592 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_290
timestamp 1698175906
transform 1 0 8512 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_291
timestamp 1698175906
transform 1 0 12432 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_292
timestamp 1698175906
transform 1 0 16352 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_293
timestamp 1698175906
transform 1 0 2576 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_294
timestamp 1698175906
transform 1 0 4480 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_295
timestamp 1698175906
transform 1 0 6384 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_296
timestamp 1698175906
transform 1 0 8288 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_297
timestamp 1698175906
transform 1 0 10192 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_298
timestamp 1698175906
transform 1 0 12096 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_299
timestamp 1698175906
transform 1 0 14000 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_300
timestamp 1698175906
transform 1 0 15904 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_301
timestamp 1698175906
transform 1 0 17808 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_302
timestamp 1698175906
transform 1 0 19712 0 1 18816
box -43 -43 155 435
<< labels >>
flabel metal3 s 0 13440 400 13496 0 FreeSans 224 0 0 0 clk
port 0 nsew signal input
flabel metal3 s 0 11760 400 11816 0 FreeSans 224 0 0 0 segm[0]
port 1 nsew signal tristate
flabel metal2 s 12096 20600 12152 21000 0 FreeSans 224 90 0 0 segm[10]
port 2 nsew signal tristate
flabel metal2 s 11088 20600 11144 21000 0 FreeSans 224 90 0 0 segm[11]
port 3 nsew signal tristate
flabel metal3 s 20600 7728 21000 7784 0 FreeSans 224 0 0 0 segm[12]
port 4 nsew signal tristate
flabel metal3 s 0 11424 400 11480 0 FreeSans 224 0 0 0 segm[13]
port 5 nsew signal tristate
flabel metal3 s 20600 11424 21000 11480 0 FreeSans 224 0 0 0 segm[1]
port 6 nsew signal tristate
flabel metal2 s 8736 20600 8792 21000 0 FreeSans 224 90 0 0 segm[2]
port 7 nsew signal tristate
flabel metal3 s 0 11088 400 11144 0 FreeSans 224 0 0 0 segm[3]
port 8 nsew signal tristate
flabel metal3 s 20600 11088 21000 11144 0 FreeSans 224 0 0 0 segm[4]
port 9 nsew signal tristate
flabel metal2 s 8064 20600 8120 21000 0 FreeSans 224 90 0 0 segm[5]
port 10 nsew signal tristate
flabel metal2 s 11088 0 11144 400 0 FreeSans 224 90 0 0 segm[6]
port 11 nsew signal tristate
flabel metal2 s 8400 20600 8456 21000 0 FreeSans 224 90 0 0 segm[7]
port 12 nsew signal tristate
flabel metal3 s 20600 13440 21000 13496 0 FreeSans 224 0 0 0 segm[8]
port 13 nsew signal tristate
flabel metal3 s 20600 13104 21000 13160 0 FreeSans 224 0 0 0 segm[9]
port 14 nsew signal tristate
flabel metal2 s 8736 0 8792 400 0 FreeSans 224 90 0 0 sel[0]
port 15 nsew signal tristate
flabel metal3 s 0 8736 400 8792 0 FreeSans 224 0 0 0 sel[10]
port 16 nsew signal tristate
flabel metal2 s 12768 0 12824 400 0 FreeSans 224 90 0 0 sel[11]
port 17 nsew signal tristate
flabel metal3 s 20600 10080 21000 10136 0 FreeSans 224 0 0 0 sel[1]
port 18 nsew signal tristate
flabel metal2 s 9072 20600 9128 21000 0 FreeSans 224 90 0 0 sel[2]
port 19 nsew signal tristate
flabel metal2 s 9072 0 9128 400 0 FreeSans 224 90 0 0 sel[3]
port 20 nsew signal tristate
flabel metal2 s 10752 0 10808 400 0 FreeSans 224 90 0 0 sel[4]
port 21 nsew signal tristate
flabel metal2 s 10416 20600 10472 21000 0 FreeSans 224 90 0 0 sel[5]
port 22 nsew signal tristate
flabel metal3 s 20600 11760 21000 11816 0 FreeSans 224 0 0 0 sel[6]
port 23 nsew signal tristate
flabel metal3 s 20600 8400 21000 8456 0 FreeSans 224 0 0 0 sel[7]
port 24 nsew signal tristate
flabel metal3 s 0 10080 400 10136 0 FreeSans 224 0 0 0 sel[8]
port 25 nsew signal tristate
flabel metal3 s 20600 9744 21000 9800 0 FreeSans 224 0 0 0 sel[9]
port 26 nsew signal tristate
flabel metal4 s 2224 1538 2384 19238 0 FreeSans 640 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 17584 1538 17744 19238 0 FreeSans 640 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 9904 1538 10064 19238 0 FreeSans 640 90 0 0 vss
port 28 nsew ground bidirectional
rlabel metal1 10500 19208 10500 19208 0 vdd
rlabel metal1 10500 18816 10500 18816 0 vss
rlabel metal2 14112 8148 14112 8148 0 _000_
rlabel metal2 9548 13664 9548 13664 0 _001_
rlabel metal2 8764 13272 8764 13272 0 _002_
rlabel metal2 10220 9268 10220 9268 0 _003_
rlabel metal2 7140 9772 7140 9772 0 _004_
rlabel metal3 10752 8876 10752 8876 0 _005_
rlabel metal2 13356 8876 13356 8876 0 _006_
rlabel metal3 8512 7588 8512 7588 0 _007_
rlabel metal3 6384 10332 6384 10332 0 _008_
rlabel metal3 14560 10332 14560 10332 0 _009_
rlabel metal2 7868 6748 7868 6748 0 _010_
rlabel metal3 12544 13468 12544 13468 0 _011_
rlabel metal2 12852 12936 12852 12936 0 _012_
rlabel metal2 11228 13132 11228 13132 0 _013_
rlabel metal2 10164 12544 10164 12544 0 _014_
rlabel metal2 7476 11060 7476 11060 0 _015_
rlabel metal2 7868 12964 7868 12964 0 _016_
rlabel metal2 13972 11396 13972 11396 0 _017_
rlabel metal2 10108 6636 10108 6636 0 _018_
rlabel metal2 6692 8820 6692 8820 0 _019_
rlabel metal2 12740 7084 12740 7084 0 _020_
rlabel metal2 10220 7756 10220 7756 0 _021_
rlabel metal2 13020 7728 13020 7728 0 _022_
rlabel metal2 6692 10948 6692 10948 0 _023_
rlabel metal2 13020 11732 13020 11732 0 _024_
rlabel metal2 14420 10402 14420 10402 0 _025_
rlabel metal2 10556 10920 10556 10920 0 _026_
rlabel metal2 9352 8484 9352 8484 0 _027_
rlabel metal2 9492 7980 9492 7980 0 _028_
rlabel metal2 8876 7784 8876 7784 0 _029_
rlabel metal2 6832 10164 6832 10164 0 _030_
rlabel metal2 8540 10472 8540 10472 0 _031_
rlabel metal2 7336 10500 7336 10500 0 _032_
rlabel metal3 13776 11116 13776 11116 0 _033_
rlabel metal2 14812 9632 14812 9632 0 _034_
rlabel metal2 9380 7952 9380 7952 0 _035_
rlabel metal3 8848 7644 8848 7644 0 _036_
rlabel metal2 13692 13020 13692 13020 0 _037_
rlabel metal2 12628 11116 12628 11116 0 _038_
rlabel metal3 13832 9492 13832 9492 0 _039_
rlabel metal2 12348 11228 12348 11228 0 _040_
rlabel metal2 12404 11928 12404 11928 0 _041_
rlabel metal2 10948 12628 10948 12628 0 _042_
rlabel metal3 13132 12740 13132 12740 0 _043_
rlabel metal2 12348 12936 12348 12936 0 _044_
rlabel metal2 11676 12936 11676 12936 0 _045_
rlabel metal2 10836 12376 10836 12376 0 _046_
rlabel metal2 8036 11424 8036 11424 0 _047_
rlabel metal2 7532 11088 7532 11088 0 _048_
rlabel metal3 8260 12684 8260 12684 0 _049_
rlabel metal2 13916 11144 13916 11144 0 _050_
rlabel metal2 13412 11004 13412 11004 0 _051_
rlabel metal2 13720 11116 13720 11116 0 _052_
rlabel metal2 10556 7252 10556 7252 0 _053_
rlabel metal2 6860 9072 6860 9072 0 _054_
rlabel metal2 11060 8008 11060 8008 0 _055_
rlabel metal2 13020 6776 13020 6776 0 _056_
rlabel metal2 11004 7896 11004 7896 0 _057_
rlabel metal3 13216 7924 13216 7924 0 _058_
rlabel metal2 12656 8036 12656 8036 0 _059_
rlabel metal3 7532 10892 7532 10892 0 _060_
rlabel metal3 8820 11144 8820 11144 0 _061_
rlabel metal2 6972 11228 6972 11228 0 _062_
rlabel metal2 12908 11900 12908 11900 0 _063_
rlabel metal3 15008 9548 15008 9548 0 _064_
rlabel metal3 12208 9548 12208 9548 0 _065_
rlabel metal2 12292 10374 12292 10374 0 _066_
rlabel metal3 11956 9324 11956 9324 0 _067_
rlabel metal2 14700 9044 14700 9044 0 _068_
rlabel metal2 14084 8008 14084 8008 0 _069_
rlabel metal2 13580 10430 13580 10430 0 _070_
rlabel metal3 10948 10780 10948 10780 0 _071_
rlabel metal2 11732 10598 11732 10598 0 _072_
rlabel metal2 10612 9576 10612 9576 0 _073_
rlabel metal2 11172 8652 11172 8652 0 _074_
rlabel metal2 14028 7966 14028 7966 0 _075_
rlabel metal3 9016 10332 9016 10332 0 _076_
rlabel metal2 9212 12292 9212 12292 0 _077_
rlabel metal2 9268 10808 9268 10808 0 _078_
rlabel metal2 10164 12740 10164 12740 0 _079_
rlabel metal2 10668 8708 10668 8708 0 _080_
rlabel metal2 9604 11032 9604 11032 0 _081_
rlabel metal2 7896 11564 7896 11564 0 _082_
rlabel metal2 10668 12880 10668 12880 0 _083_
rlabel metal2 11228 10920 11228 10920 0 _084_
rlabel metal2 10836 11816 10836 11816 0 _085_
rlabel metal2 10276 12936 10276 12936 0 _086_
rlabel metal2 10052 12908 10052 12908 0 _087_
rlabel metal2 9716 13356 9716 13356 0 _088_
rlabel metal2 8540 12208 8540 12208 0 _089_
rlabel metal2 9156 9464 9156 9464 0 _090_
rlabel metal2 8708 9464 8708 9464 0 _091_
rlabel metal2 11536 10892 11536 10892 0 _092_
rlabel metal2 10780 12936 10780 12936 0 _093_
rlabel metal2 9044 12936 9044 12936 0 _094_
rlabel metal2 8316 11368 8316 11368 0 _095_
rlabel metal2 10136 8036 10136 8036 0 _096_
rlabel metal2 11592 11116 11592 11116 0 _097_
rlabel metal2 10108 9408 10108 9408 0 _098_
rlabel metal3 7336 9996 7336 9996 0 _099_
rlabel metal2 10332 9016 10332 9016 0 _100_
rlabel metal2 11956 8176 11956 8176 0 _101_
rlabel metal2 12292 9660 12292 9660 0 _102_
rlabel metal3 10780 8540 10780 8540 0 _103_
rlabel metal2 11060 10668 11060 10668 0 _104_
rlabel metal2 13188 8960 13188 8960 0 _105_
rlabel metal3 1239 13468 1239 13468 0 clk
rlabel metal2 12572 10206 12572 10206 0 clknet_0_clk
rlabel metal2 7084 10612 7084 10612 0 clknet_1_0__leaf_clk
rlabel metal3 11620 13524 11620 13524 0 clknet_1_1__leaf_clk
rlabel metal2 9548 9044 9548 9044 0 dut53.count\[0\]
rlabel metal2 8232 9660 8232 9660 0 dut53.count\[1\]
rlabel metal3 10528 9548 10528 9548 0 dut53.count\[2\]
rlabel metal2 12348 10402 12348 10402 0 dut53.count\[3\]
rlabel metal2 7476 11928 7476 11928 0 net1
rlabel metal3 8344 14028 8344 14028 0 net10
rlabel metal2 10892 7602 10892 7602 0 net11
rlabel metal2 8428 13216 8428 13216 0 net12
rlabel metal2 13860 13468 13860 13468 0 net13
rlabel metal2 13524 12936 13524 12936 0 net14
rlabel metal3 8596 7700 8596 7700 0 net15
rlabel metal2 5628 8596 5628 8596 0 net16
rlabel metal2 13692 4312 13692 4312 0 net17
rlabel metal2 14924 9968 14924 9968 0 net18
rlabel metal2 8988 16240 8988 16240 0 net19
rlabel metal2 11732 13300 11732 13300 0 net2
rlabel metal2 8988 4536 8988 4536 0 net20
rlabel metal2 11144 6020 11144 6020 0 net21
rlabel metal2 10388 13552 10388 13552 0 net22
rlabel metal2 14084 11732 14084 11732 0 net23
rlabel metal2 15204 8596 15204 8596 0 net24
rlabel metal3 3178 10388 3178 10388 0 net25
rlabel metal2 15484 10108 15484 10108 0 net26
rlabel metal2 11088 12292 11088 12292 0 net3
rlabel metal2 14084 7616 14084 7616 0 net4
rlabel metal2 5628 11144 5628 11144 0 net5
rlabel metal2 18956 11312 18956 11312 0 net6
rlabel metal2 8876 16324 8876 16324 0 net7
rlabel metal2 6020 11340 6020 11340 0 net8
rlabel metal3 14140 11060 14140 11060 0 net9
rlabel metal3 679 11788 679 11788 0 segm[0]
rlabel metal2 12124 19873 12124 19873 0 segm[10]
rlabel metal2 11116 19873 11116 19873 0 segm[11]
rlabel metal2 20020 7924 20020 7924 0 segm[12]
rlabel metal3 679 11452 679 11452 0 segm[13]
rlabel metal3 20321 11452 20321 11452 0 segm[1]
rlabel metal2 8764 19677 8764 19677 0 segm[2]
rlabel metal3 679 11116 679 11116 0 segm[3]
rlabel metal2 20020 11172 20020 11172 0 segm[4]
rlabel metal2 8092 19873 8092 19873 0 segm[5]
rlabel metal2 11116 1015 11116 1015 0 segm[6]
rlabel metal2 8428 19481 8428 19481 0 segm[7]
rlabel metal2 19964 13244 19964 13244 0 segm[8]
rlabel metal2 20020 13356 20020 13356 0 segm[9]
rlabel metal3 9072 2044 9072 2044 0 sel[0]
rlabel metal3 679 8764 679 8764 0 sel[10]
rlabel metal2 12796 1099 12796 1099 0 sel[11]
rlabel metal2 20020 10276 20020 10276 0 sel[1]
rlabel metal2 9100 19873 9100 19873 0 sel[2]
rlabel metal2 9100 1029 9100 1029 0 sel[3]
rlabel metal3 11088 2044 11088 2044 0 sel[4]
rlabel metal2 10444 19677 10444 19677 0 sel[5]
rlabel metal2 20020 11900 20020 11900 0 sel[6]
rlabel metal2 20020 8652 20020 8652 0 sel[7]
rlabel metal3 679 10108 679 10108 0 sel[8]
rlabel metal2 20020 9828 20020 9828 0 sel[9]
<< properties >>
string FIXED_BBOX 0 0 21000 21000
<< end >>
